��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�}�\�$}�����,`Y�U�m$�f̾rc[eR\���?CɆt]a�B���R���������ʥ�+�[���R��0'>�ϋA�����/���;㭤3�r���$!�v	�IL2�����w�џ�p[9�v���t�MQ�Tz���6��M��R&U�֘�ntG;����X�V9���|���:�p��S
����Ǥ�.�|/�~�Gy�J}���c�W�|�Sp�ʎܷwJD�k�7����h��;�#*(Z?��Q��F�\>t�6l�X'��N�sU�ʗ�y ���bӖ�m�rC����M�P���@���Pt)�{I��Xމo@jd�t�O
F/�:z{�o����fq�L�J:�a���ǃ#��yQ)	���f/?�j������_O'�8��j=؇�(��&�9��4t;1d�����?>�W��G�4���Y�}OG�r�/:
$��p�a��ŭ�i�[�%�x�y���������as�<(�v�ɐ2�� �oR@l`��Ģ�U��b��>e�*8-+�G������)ۺ�NQ��u�̸����#T����!��r�U���HQk��o_V�Ewp�Y�9�?x�Q9H���a�>���,��>�W_/@��J
5��}�\r��=����#f���8�S'��N�4��^r-=2􂴁m�']��$-J��v(L)  W:����H<��a��#�s�X���
L��S��,Qʂ4�̩tr��0
�5W��F��\a��b�������3��
ۀ=����.XG�c,J�"r�`�� �i����48�f�y�4t�Nk9��-��C�&��+��Df;[qs>��������y��j�hm�=����^o�e�F�V4r��}e]�.7�i��-���4p�q9Qo�$/C�� �/[?��0D��5G���1�#�
#g��@���D�CZ�-�#d���u&v�� (gYYW���"�n[���� �#3wX����!ᾓC��(|\0ng�z����	g����	�HC�c �X������xgPM	`V�GI�H�pc�+cJ�|�I������9.܉�Ăq��a'�8*Z@��N# ��y���ɕ�;%L�����ǀ��~�T`-L�؈�Ω��	�T�&L���j�"��Gy�*�@a0�-���`9W�]��d�����$����� S>�����X*�孡��kgN�{��T�o�pmk�aQUVۣ��t2����alB�n��h�퐉\t����x2s��;�3f�gc/���K;����lȕ4<Y��;c�q/���e��1+�mݾ�Ʀc�ss�^��,��H2��Tf���nV�s�>�,��ԯg9�V[��^U+�)aGB�(�14�V\k<c\�!5�����K��� ��y��^^ka��e|��T0X�Ɇ>��Rr�3����L���Q�������/�9�1���v��ZE���o'\�.��s���z�~�f{���	ҵ���:��v}�P��/uȝy�SmO�'ݩY�T���&���1�:Ghqh������_�����"[(�~��yu��[�M��6L(f�!~��*+#�-mڦ��*�Xs�8�n3���. ���:f~>��q�n��r�������|�GܭLֈ�q��~RMy�V#X�Ɨ���2
�T�*Fmq�,	؋i��sO�A +�����"�� �fk�N1M5J4GƫԺ��,��H[����݈�1���*��4�4�3f~7�ؑQ���:z֝���Z�s(*�,l?�X����=f���{�h���b�3�D7Yk*�t��$K�-�ˑ��e��V���>0(q�áϟM"u(R>����J�([�ԇ�l�ڴ��qy캋��7������#/N�r~��+q_qF:4ڰ�W���8��2�wO�|q�;2�Ї����H��}Ŧ
s�hx�L
A%a����f-gb"M�v%����Cnd^x�<�j��q��h�_�'��	󻬀� F)�	��ؘ\r-�7ن�ԛq�k�ª/#m��Ё�����
���j� BCB�����/��P��	M��=���P�������F��u͘��|�sYyɷ����M����ks�ء���(,��ƕ��\�6�'���BW���_X *�E�'�a不��h�H��gN�^Z-R׍2y���(���v�U�7Wy���kE�1/%yaJ�X>���XJ�L�� �1������\�C��	���g���'lئ*I�y����yD@��c�ƍ���j;��%ՠ,gy-]�����pLȄa��O�A��֌xu�皡�O�`�6>'�D�"�rZ�w�sJ��[���k�@Zh���N������k���ěT�mc� ���E���KQ����ì��G�И��p;,������A��
��Ft
�����eŸ�(� �b$r
*X���#����	��a �`��y�x[;y�#/j�@��%����(z>�4s��p��@n�X�-x����U�U#uU�Yz�.T�B��D�h��˹������0:'g07�U�;�-ڰ�LF|wH��9zJ �\z1?��,N7�r^�y���#8��zA�<Q�l�:GPD\Ͷ���O4���h�K�|�Ӄ�g��h?.BdF=T��֬�����9Qf��d�	���lu;K���a����~�Oh5[�Q��i���f��u/��.���JO���1ꨉއó���T�c*�#���m��n5n k6m�NY���Z�z��XI���N�FXu�\�!˓}�W-	FKy%`�u>�ڮv]7�
J�=F��˲$TG�\N�����V�/x��k{�_����A�.��T|
�~-d�o0�nl���fo.�檲�Ű����X�k�/V���{���Y����6n������C�(;��P>Fh�
�>�#5eˀ7f�ZC�u$�uo����YU���P�&�}\Ϻ@�<�a��1���(�m.cM_�J:y�X�8(��xy���.~ːc�=�����kb���i������D��p\�Cp`˝jֈ��Ӓj�x��6m�
J,���	h���u�-K�K�>`���g+ Sw�=�n�w�k�~Cu�|`�#\����;�k��AIŜ]���$tjaB�K$KBy�ٚ�~ɘ�F��e�x�d�ncJ����s��}��N�� �[�2�l�$J�r��{�͓_�7���bu�1�]|��l��eRg�U:���}��h[;0�,ǣ<�"9��"������m	A�~����(���N��`�ۍ� �͹���80�gg�^�#��t��znΈ3f�Wo'��lm^��[Z����i��֙�u>5.L�f���R�㔸��I�iu|��I=�j�"f�X@�5d��FZ�E[���9:~Mɝ���	H�t���	�3:c����D��Ш�O�g��Ԧ>�*5m/x�vd|"y�=H���[x=�|n}ϋByM�j�xV7b���]몺�&9��8{��A��Ѯz!Nt�;+ ;��4[7�55�#�� ���t`�[�O��j�7?�;i�h[Υ�R�>�ʍ��T�g�H���yU�s�qg9Zbe&�^m��8ה,ZM�����Qޯ�� ��ѻ̗�6g�x�'�!*��u��T��fj�� R'#�f�I���.�=���L�g!B�P��,c�\](߮5�6{q.V��EP�����
�d����=����Kos�m�:`�(���܏�S�Y�v�^�7^���ѽm+�fz"4������{���&���ot�o��Y���%���m&��T�	��]=�"8q����pĲ\�*�!6ED�7:�s�j��㻔�Y�����"�%]H�FuS���p�g{FӶ���QT�o��$yl���kO�Wٷ�����J^ E�h�Ja�4��kE�f�?1�~6��g������ݡY�FB��O,�Ø��%�?��$<�@q-%��+�/hT�s��b�O�YI.b 1j�E��!���"�+V����J���%��3"y� V�_����[�3&S^��7%�Χ�7C `m��ɰ8u�k��!D;�1=J��P���'ˏ�����n��ĳ7R"��Ѝ�ӂ6�q��~��	�[c�[��b��x6��e��e����/�"����c� ��FI�-f�[0߄8�*[t�QiO%�2�r}���>k����FR��6;Y���Z7�W&h��?�>���$9/�Tۤ@������O�����L�R���_���a��@��q�>��������=���a(L1�iο�$+���xU6����`�t���n{�7��f�9r%/��rZA���esZgw�u\�4�,�$�g3.x8�&�D�V.���lp Մ�P��ڭ��p(��kҳ+C�@�Z<M�wܠB�Kg���x�tC�gI<�vA},��8U^�)����g�f�L�3����t��ES�	�J������uHv��lt����И� Ō�õ�Ȑԣ5ؒ�g��tNǰlP�;G�����R^��TK�+֍#�7 �U���'��3���	V��W�wL~.`U(��<7;��l��?ʯh�x�-��g)���yܔ��
[��6�Һ!��H� zZ���� QR�9�CQ�hQ�SFFs��Ŧa� ����m�!s����>��U�RLp�XnE��,��#�w�³������3 R�NE�[��J��>VW+�<'dA>�ZVX1����	We~wLIXz=�6�6���pJ���@����,�z�)�b���p�����S�TW<�]�A������ɩ 73_ׅ#�G�!�bٳf?�����B�����%1�uۊjH�M�*v���\���-�6����ȍ������n�u�����p%;3�6鳖W����k�h(��8}0��#_R@Ȃ���}�q�{��8�q�5}�=������s=(�
�Z|TH�H%V�Q�g�ue� �� l��c}���׊い �a�f��	"j麱swx-R�OŞ��^�L |R��Q�Ç�$�).` ����p�T��7�V�r���I��/��I��)b��r>*v�+j��n߹-o<�-�� ����q�cU?�\�� ����m���B��	/\8����
����4'�e�z�ʋX��j�#�~ ��G|s9#�B�Jk��/�hT�a���t����k��ϲ�����u=�����k��D�}�^iv!fnR�����b�K��w�EY4��Oə���X1G��?Z������Nl�9V�Ru�fo��]�q���3�#�)�J��"��J�qO��yt�� ���\�[)�O�yǶ�D_���̯o�lѽ����w�X&��V���$ֵ]W���<��`�f:k��	��h���m�Y�=��)U.�v9.-�����
	��ث��Кԑ� -��&0��!<Zbs�ǔ9�\g.��No�TЋ�ڧyG�}
b�ACd���}D���[ц�;��ԭ�L�KCqܴz�/�NU;ݥ�*-�̍��=Z�:�.:�@8�=>-�#�.�|~y���fʽd�"yRh#L$�W���Qb��Ud��Բ��c}k�Ꟙ����=�P>��hw�^qAv���
6Z��#hG��76�ܘcusD��s�E�Z{��nýt�B����ϓ�Ryb���L�S�`�"���d���y�<kndb��p*2���9z�}�_�[+6���	�N�o/�J)Y����y�0���)t`7����!�(R�PM8_�����r����c�M�ܙ�p�A��0��D��C�k�<���J@�P�xW��bw��?"�����@��-�xm]`T4��}ĩ�̣r�-H����>(��<�_����nSkBRoHJn8�`�nv� '�0~�I�Ag���n�Om�L�'ρջJ�#ܹ��dr�`����K��b��Z�`�/�Aq^?���m]�����O��1������d��,洅4M2q�1U��!���0-��u��_%�M]P_�Y]�_���V��~G0 �"�S�0%��H���t��O����X�����H�q�W>��$y�p�TXd�o��0	�X��y�o��hO]�c��c�8s0�^F0�E8v?��,/n�����_L��rB�:`����M�I�μ��1���a�, �1䀽�=�*݋���e�4+Y#r[�i;�W�´��}����϶B�lȀ�e椼dL��܋�P����;Ħυ��ןJ�G?0����H0&V��^Ǿy�UP򨧑�(��*�#�2n^ɾ�����{���c̶m��Ep�4��Q��m�b/<]*��S��vI�n#׎㿾�$ŭ��)�5!=�u�oTtiK��g�t��skZVYN'�&���|��M"ⱆJj��b��Ʌ��]��^��
b*�U�^G5pc�J��7�6�L��	FB�a���iR�L�b������0A�_�q5�-��<�9F�ZM�5X`r�ǰ��o��AbT�C0�+;,򭳝8Nl��@j|�Й\uz�7W��L���߹ї���m�Eor�ܤN����~����ln�YP�j��GҬ�r�V꫼�6�]��d%���N�E�P-�ܶ�5g��in��ʽ�EmD��b�B���{����T$����,��?�H����%��� I�褫�*��2�ȫB�'O�es�8�H��%}i(�jt2F��bT�	��7�k�"'x�v�c��);-}R;�ή��/Y�U�*���#(�nd�ނ���Ol�n1Aj�]�G^�r=��"a�z%��Ɂ�pO��t�jRt��&�-�C��9��Q.ةٷS;�[S�ci/������F����Ӹq��8�է�L�Bb�)IIIJ��t�P�kP�i��k>G4�.,&��@�����d������k�}����[��)�ᶽ��;z29L'�-8
(����������eE�/��Sn/����E*#8�ۏb�]�Z2z(NS����l�z�ϢZۢ��:��B�͉�F�`�R2���`cc��`����=Pu[k�% 1��y�#|
��㧑N@��vB�5R.��k���C���e�?p4wkҗ�-o��%�[�z_�r3���(N&��ӦT�x��I�"����X��H�0(㾣u�.F/N�|/OgVUG��U���b��L/��
�����7:H������<��(T�R�V3;f;�6���ٰ�&�$��G�<�$����Tڇ4vzӐ��y�}�	��9�H�*�Ծ6$��N��'�<�I?�܊�=�~��V����A�hx��I�:Ln���;������2\�0�����'�
�.�o�h3��CFG���H��Q.H����|��{4��� �K���Ĺ��V�4"�?	4&6�v!uVυr��*��h��8�t�4����`Ǆ5�A�C$������cW��ի�q��6�.��B�8��hکc΀o������b��?����*n��_V)�Pyכ	w�֛��5s>	�@�-� d\���\�UG⑎z�h\��t\X	P8����c-b����>�@�5��%�5��L0��x0A���T�k�=��U4��)��[��`�pl��e�Aw �~L'1l�l`s+�D8\��o��ر�F������⾵�d��4s%4Ͻ_9�@W��~��]Yb[���so�p|Rk��z�v��'O#��q>�x��&�3r4���1aalD��I܌{�8�Q��;��������I����E0զz��^�7��k��uw�V#��QM}J�]��n��MN�c.:��#��'�Δ.���\ޝLm��>�h�8���}߂�cL��v��rkȗ�.�^6[,��L��Ҭ姨`珱�=&�4��iEIW�L����>����V���Q�������@�/�a���]q�$�LTiw#�K���u��[bmb6kjאnHMs�wRi��� ��'�oP'm��.�ѫ3�j]�b�p���$� �y5UȟubD1����79�oϞ�[����uɰrf�naԞ�2�����[�J�i��G�$���3�o7� !S!���{��Y�j�<T1jO��r:�D!.���gYuF�6�?ύ;�v�&�_q&XCgJ�%.Q�P��~ꠜ@�.f��~T:�wX�D<V��8{�D���m��)�+��T�.�0}�\1�~|j4>x=h3�����tɁ���%\۳/�Dd�Il.߭Qi����{�o0?5����rK�c׸�!=S���i?�[0���^�U�(nd|��l��k1�cذȻ�`is�����6��i��t.�Ӕ�0�xE��!�G�d�,=v�.KV��Q��
^���V"�����Q/��	3��]��G��V�]=���!	��l+ߚ�x�M�k?�`X�g�͝��A�\q�zB���݃G]���Y��/� ���1�E���l?t%Џ�6x�F�y�$�ǓC/��T�~�S��2�Ι�o����j�/�	�C��F&Q��a��/S��(���e$�WW(sh}�}.M�������CȈ�]�lo�uU���� �Eh.`.A����4!.��@���l��\�14����Fc4DGR��+<Ҏ_�/j]��.x�מrQ&���R�R����*2�֔9���8�`V�'�a��;Tt��Jzx�v^���k���ߡQ+�J���+����.��j�6}HW��R�������핚[�{B �d`�o��d�3$�ܜ ;|��	"O�Lճ��<4�e������}qcS>c%r�;��l(�b(��C�!���(����`6��[�:��{���c��aqP_�W!5E`*�c=�般�c����:�]�ژ�	�����:T�yGY;0�p��g��;���-���h���l��9���ю���d7L�ڝF��E�}����M&n��o86an�@0X����^!ZwZM�Ge�w��"gj\Y\!����ȳ�5�=��e��Q�n J�""6@���Ұ�|����L,/c<I�)P-��l:=��ni����z�A�&���7Ri`8��8�M�)|�`�U"cV�J�E�&����O��h�nG,�< �i���gRQ=X����ŪD]-�e�\�t���/�;"�����K����Z�%yh�5��gHa��Ǩb�V�oR�`I2a/���l�Q���ۚɹ���x*�z9��d7]������6}q[�ujB�}c�3�Q[���Եqo3��y�x������: 6J����%�BH�g�0�o�M�[(|M�	v���2k�j�ͭ���pQ0>���ˏ��ܩe��[i���X�f<f�Xgw�\O"�����ﵐϖyN��SEv�͚�#>y��qG�h�Pb�qx�̴���������/5(�1f��#�"���׼9��a>�D�)�E��.���ҿH����cj�����;y��|�+���*�����t��dHN�}���X{(�j��G��:?"�`F�w�az�d��4`�?���=6�ѱ�Dx��f��.�s���j{�ST���fs�����csC�#6&^6�-'��7ͳ�Ŋ-�1[��ߙ�|���a�3�B�}h�ݨ��m��I�SYt���«%�Э=-�cY�L�T�5��t�^�٪8�T.�6�<���=K�BENf>$�O������oJ쑯�bc9��+Z|>a�X���ື_�[�e���	�#�D��������8�����jt�k_�g،#����}!ò���:A����\XCY+�����x��6�1��ȫ{+=�G�=��X�&?��RrZ��W%��Fj��g���
n�����P�7��������9�P�E��e��#�نb�n���6�?���
�I�ަN�jN��}���zr w��(��NLbm�R������c����W)��vC�Y�|�%�+<}���,γ��7��O�5|E���������f����Z��d�M�:�F{�*���҈�6nwS�٬=Η|.L�Gh׃�M���OM������Z]}���������'Jtd�`�~N�a�!��jIhՒ��f�>�h��S�0�[�K6f���%��)fF:��Q����)*Lt�̻kA\D5�^���$7�Й��t����Km�����K��}�Feq#��N&�=�2nm�jԠ��ȵj�;���Ag�5�|���4&:�H�;�֌��q�^ XnO��@��_4�eB���"�WJ�<l�v.��j���C�|����D	�����"H�/�a7y���/�'���x�9�>�L�!�þF�,"F�Llb�O}wO�M`Fz��R/IW�?��㍙Pk;�bmƋj��-�\&.������{8+�
~T�>�0���/�9���:�"^�l�.�|����%u����j���&(q��S����o'Ȇ ���j�M�x�g�����;����k�m��O>�.��Y�i?ԮwE@Hn�8�k��߮�v̷Db:<T�O�����Kֻӈ�e��<���������\�m��6�|$�m��2>��+�M���4g2��4��66������ټ`�}x����m��NFH;S�t먫b�Ѵ&��~yq�<Fw���;E�f��:�����|ȵ^�%=������������*�.�SpO0S%��ѿ�@��I2]ӿ���G3u'��'�̵rf�^�xV'p����\�L�it�'?˭V�۱qaam���h�&���c������7~2A+�R���[z/�R���]ϟ�Vu�C�_�m���$�G�����c�]�,fb�#���T\���nl'����(��2�B��e���6�@�<��8�{�.�r�څC�mvH;��u
q�~{�z�P��;tbx����n������6�Mۧ7v�������~$�@s�x4��H�����&�,�xp�`B�M�ܹ��V�j�^���4�[�InM�n��&-�5�\E��#�kD�hmV�㐶�&�j�`%65�\QF��)�C��e�@\� ��f���4�w3~(b��3�$ bͫu���w��8/�]�=�<����`�z����?!x��ymf��ō�?Se�����;j 7�YS��9�s��n�G⫄�A}��sBc�}<�?Cv��-�Ţq��&�YC�z�h<r�'c\��Kn��q��qC��/s`��I�P������pـ^��Y�R\�S�������a+�OZ
�DUޜH]�;�W$��0�<(5�������h4�+��ɒ�5�<’.�O<ii۸t!p�XM�"c���_���jy%�1,��}�蔤���0�V�v���uy9�� ��0 ��m+x�RQ�����q�$sf�� ��j	�:U�QNש���q�m~="�{ŭ��;���.Gf�����[��M�Z�wgeK
�@���Ş8V�5J��M�o�!����"�RH�:����ͅ;l�;����ό(��j_��&�0i�,^g~�a�����ȹ *�#��[c�ءM���;|������z�k��JW�q���3�T�+�������U�$G��T�YR�ƓZ|����A����.�V�u�@E�d O�"���&]�|A'������a��qK�BO�\���ހ��Ij04�/�O�_p��L���ֲ�	���:Mχ4�� :Ox�P�� ��v�c��*���o��#Z�����|�}p�E$MS�:���]�^� uu�7#���� �7� �Q�x4"ǟ�R�@���S*g�tTQ�^W��$! 0.�nI)�� z���I����*ϩ�dl=V��z�����J�&2h� ��͑fR�	����n �Y�0C��Vk�>�C�Ӂ�:�O���W?��n.�}���_��}������R}?�a�kVrD?_c\`�s�nR��Z���-Ot������	�C���#���h*d7����*����h��r5A�� P��=Z��������?��t6X���&�w]^)���|l<��xy���%��d�Z�Qs�\�N��*m�jA�~UVf�5�QN�vD��b��}p����/���t���ǵ(A��Mӆ�J&�5���?�XkL�M�]��PҺ�?v,���?&1)+2�W��4�e�꘎��X�6d�SmtT���l����/�/�{Lإ�k��Z���U>�\X@�`�ӣ֞���ώN�y�_���MA�����;0�9X��H/?@�~յ=o���z���*s���Ȟ�w�#^�sjà~'>/��G���N%�����̹i`��E�YWjr֨
dPZ���7�ǔ���d�**�����~���a���ێ�g����߼�c6�a���J����ʈ��,��U���'��xf��xU�,[��4{q�}Y�MUr��� �Z�L���uk�m����i'���J�	�`�a��7J���n�G��������!�h]�Oy�W���1$���!U�,�)�	�Q6O5v�m ��V���u�,FT�O�U���h�P������	���e����d�^�4���۪���)q���N���t:�]�ٷJZ�O��`�N��!1yr��]�)�jV�����ro��{�'�V³@�U/�j�������
��lK��~c�?������pN���_X��D��t��<�)�Mp�cIлH�	����`v��:q��Kx`3�qo�`���V��8)I�A���PǊY�{�SX�g���^��0�q���,��չ�uS�Q��\ޗ�)/?�2�U��9i1m)��}"�=�r��oW�g-�o�Pbe;��$!<���5,g�$��%�;������P|�`�0�xS�?
������X��=��3RY�❦6���m�u��m~L`s���P�:n�{"��g5����$�X�)^��?�i�ߏ��&eE/��!d��]��Q����k��1g����|�t#�~+��Jm� ���������%8��?�7�Pd���w_Zd�m�Z�u�K�F�/(�Oᒓc#Qpr�ZPQVi����5vA��yP��+�:�c�	��F8�OM�Ӽ��bp���\#.� څG���#H��&�V��;�,�,lu�@"���6�:�v(PiBj_D!Yvf{k��-�K?�ev�9�()�Ɵ�=s������mu�P3�|)�#HV����uΝl'�w+:�!>|�8i;�J �g#��|8�G�yc�(?c8�)��q���F�M�L�
�S1����N���rL$���C���tȖ��x�AŸ��Ҹ�?�5*�	�j�_���:��g8��N�w��i?O�NXQ��]��d�"t��@ �yA:|���u�O�/���vZ�b �Օ���O��Kᱚ��H�-뉴3x�={�C�Pӥ)�p���<0��^3JbtT�k���q����4���Y����[����is#7���e�pQ}��]<�_�)/3.����ʉI�$A���q��qr�W�BU��:iSz%͵׷�Ty_�!���Gr]m�3:�C|��O$̚�kZ�u� ݂0�(ֽ�k��0��?�!�m�eKT�`��E����A��uN��̾��q�P+�Ƥ�Z�h���V2Pfb_��1oC�\�	�����=�u��1�U�oyv?�3�'�p�}@�O�;��P'ցȗ��ݩ�9��b��3�f9Fb҉�ix�Aʮ�S�,|[;���{l�����	{�"�W���Z��ɣ �f��Q��꭬kK�6md�m3�z�`�=|�F�d����Fc�C�"s����4HM[���&���s��]Xm"��F�O�77��a張~7ȨǓj��vqZR�� 3����0i}E��f5�T�B�2��!?�\T�uX�ws���๠���jؚ~�L��t�������{�.l�N�����n�j�+.��x�.��Ⱦٲ�;~ؼ`�<�ixeخi��@(�pѝ�EF�י/mr�� %I�'�6YѦ�k��6�^��Ep��T�Um�1�xM���6�O��{�>����)d��&���!n$J8mT,�I��}v�����)C�ҡ�@ܧ��c��>^/�T�N�5L=������T����j�O�dBba���p�4��0������"^�e��g���k&,W:3��H�Ky<��x�vdv��&�eNz^�:i@d��&{�)ج��Al�;�T��[1*�6�[/���D_,�
�N�'_q�@C�͖�ŭVg�Ғ��J]���B=��XJ�x�<�Z���k�4J���q�qY�}@l�H�5��:X��r��jX� ��x��>��!'DK4�nV�(���+!����f`�I؜i���337V-��.��8Ch������v�n�DeA��0S֌������B���dF��~�s���;!&h
ߚ�G��f'F� ���.�z O�w�1�t��_�V���H����v�� �N*oǋc��H	��놿�������Pw�ݺ�$���r�Bl|�z����A��@YR��s��E역�%���=�����O[k�2O��"��4�7Ì��nDf�K�hv����ț����Lń�80zi-b�T@�Rඥ�?,��o����bj`J�c"�Ţ�`�r�N�F��ƺ����HR0�,��-�;E�w�vd̎[s�6À��X��ְ�Q,�^���b��7R���Q�{��������qw+UQ%Ҩ�G����b@W�=$�$yeɗ��ڐ���Ȩ�0�[�3��	�]=�E��m�����~+�"�V����9��i��q���FC�$�&��8Т�+=cbK��:���,��=���N!qw��%zR��J0P��&��0��!�����7���To?�? wH<�~ҥK_91.�e��=x��'~怔���_Օ�,]�\m�yEʉ�)
�
��J���Z��X��K4��d�/�ȋΘ�7�f�j�i�]�j{B���4�J�j)ZSr��6r����EY�8s�:�
5������u:wD'�� x��m�Qy�Ӳ]�.$��<Ӑ��>Ώ�tM�$.�3Y9J2/V6L̂P\v�W5�R�ĺ�e�P�J����q'�^"�CL/��ߢ�uB������"v��/��L���,'�,WTk����<�	|��P���@�F���8�=ý�Lw5m1�_vtY�
@ږx��Ӈ-9���`$�˜�}c���bnd��p�|��9�A��N��8�#�e[RfA�=���.^'����
)�4�����,s:��&(Ma��k5b���¨op4)����ˇ�����9����t��(����s}��%G���OS-P���~T`�3@��
Tm�-I[��h�϶|��"�!��	���ݞ��#5ګ�����J�逭=���۝�/s*�+	6(���=$�
ܜ�g�Kc��;;����~���\S�2a�1mH�5��X���v����\�U������i9,<+��} ��{y�4Wm3��%���� �V�7T��}j�g«5������f��>�;���O���V
+QEW<Z��X�1g�\�.�ڟ�;a3�b��/'�.}��,��qaq��1I��O�Rv����5��Un��������,�@��� �	ta�[4$�6��,��8S0'���$$�ůh�8����^�>�������9�yK�g��{3 �SV�^X��Y{����W�V�1
�M^�_)]���Si��B��[�
��XT]ҳl�R!�à>�l�PX�y�C��<�TxY��SVgv�/���A�XN�$�=�q�X7���=NSX�dD�	��5��kG'�y[�y~�a�鎙�u�
U<c2��5#�T������s�2�q�uX@�Čc��T"Cn
���N�]��[]K&���t��y��R+�rm&x��M�H��S`�NhK��Lq'c5���l8�jV��ˍ��Ǌ:��u3rL��Nx$J�`v�ʈ��.Hd�g�9S��jwWE�����Dy��k�s2�4|z6�H�.�-]��n֭����)�m۔�¬|H�$!H[8��A҆~���^M��P]b�*�-��vڂ����x�̦�"�Rp@'X��3}�r��]&w��J�"��1�\ԉ���A%��Qx��j8��`MSJ�|���OM�/��SO�~�ƿ�֚?��`�Ɩ6��'��%����6���$"K�m����m�Iʀ�(p����c����B�{�-�CPJx���8��
�Y��BRR���ojˑ�a��d���B�����#;��4^�ٮ�6�N=|�~|��2��;iYMl�����Fٱ3<�"<`�8$|/u1+5gK-����8�����У�C8����]$���lYr0i8_� X6"��H���"�P3�)v�bx)K��6�D���-�@4��^��|4F���S�,k]��%@�{�&/)�Q�rB2�}~���U��O��s��b3,�I�&EE�K�,l��ת�D�����(^������~n�I� �?mc��	i����aA��0i�O��j
T��($�m=��8}�/��V��.��5�}ٳ��y�I�� 8�-;EO	q}��%L�x0U]�
���;�[n����}�K_ԉl�'�V����8Ҁ��)������mc��Iࢮp\AⓂ�#�q?��2��tYZZ ���uSHh��n�Xm�W��Ĥ���O����0���~��lk<��Ӎ���4�ۣK������yO��-��S�C�Q����NLf�{3�`�^�h8�ҳ��P̀��({F:��ѮÛ7��p7�4��:�P����9�DկI+�1��F�Z�m��̢E�]�a|�fl��V04w���!�ۢऍ	�p�49�>��m��tR�%��?	�{�,��b,��N-i�
T?�/i0I�O�3K�&��7J~�B�yP@�����awb
[8��C�T�]�`x�z��6/�=S�h.��T'^��;�F
Q[���`>viXAZz��Q��[\�}�|u�KR/�����qW�E���ҧ��령ϰ��hd�b��Jw�] ��qkg����C4�ϘOr[%CLԱ�ޠ�w��$�/�.p��e{��� �[����c�����^��bm���,Ú]/I^l�9Ɵ�b�O�a�K�M?y��/�#$U�n��;�jK�\|6���8
�R>�} r"�r���bֈ�OYR�ن@�_S��+�W�y��5�̞�K%��$�jR
����&WZ�qD�H��S���i�HNۜ�˳�k�.�D\t��,��FgU�H��"�U�����`�^n�Z���`2���\"궞���q ��QŨ�.�/,Éy�ꦈ�(�y��k�����o�I؁�������V�Y$��t֋����u
q@�1ѭ����0s��U�hV���fu'K	�.��Qq�a�3$x����sv�k|��Vk3�y�ȕ��]c�(��� ���;�����DE%c������\���˷w;�5�m�d�,�{35g�%��zH�Q�t�3��j�,�e�;i)L�~�o@ {9TO:*E��N���p8�@x��9�P�&&�0�UF$.8�^]�~C��<�X�?t�mӤL�F�Le��RF�zx��%]�z.P�;���ju�_��3U��������UO��z�r�<y؏��_Ԏ�ɮ�	5���C��'�0<��~R��;
��EH4���ScD���emOJ��c��О&�u9�E�2sLSc��.�ok�N�WQ�
Ρ�U� Ë}ip�rʃ��=p����0��*BK0�r���Tl�t3��ptŏ���A��%��0R�� nHl��
��~�h�&XMm�ۏ&"Z`5�dM~��"=	�e\n�t����=�w���N��6��(懂�=�n[��)��Q��Ռ��� g"_�Y_h�$l�B��Y҅��;�S�p����۶���7o�
��������C�'�[��Ň��@��i-_IZ�y1���s����i�ғ/1�d�����{��/ml�o����R�y ;z�&{��#�$�:W):�cɅ<�c��3�Jvo���Dr��jF��RC����N|i�w� �����|�W!JQ[��;aN4m��� �/���~���7������FX
T�3�,eS��~v�ͮ�=�� �P��cE��W�|C��<�h,a���%��D�%�?�w��I?�Nt�=�-�0O���0?�����2��o�UΊ�"���&*#�Og�H&}��O�<���^�������1���o�e�}��X,���3	��[� �.��&�+���~�J��!|#V/�m���d�^bŰ� \b�i��)�w�~}Qb�����w�U&^y
�C8#��f�G�W*�-�B]^~7�YANdZ��Q��z�>y� ��܃M���t������o��(S�����s����LW�'�*Sy�a7UAy���P���w��I%5x�%l2�x����5"������j�3%#�lٲ�k��,+�rf˫�s=��ei$wV���`4������u=H�a��̦�I�P�2F����bqΥ�X�U1�����=[.@U���Us���*塋�(�:���u�nm�
�8�%���(����$����o�\�+O�~�7�w�}6��7b����K��eaE���87x8T�)�\�#�4ǧ<���}'���E��=�7[a��n�M���ZY���M�x��V�A�+ݵ��Q
?3<��nn$�Y�R8D���E<L�MK�����a}��`U<s�Xs���/vB	�'h�.oo�_�Dc�� �]S����V�5�0�7���qZR�C��.�H�U�Vu8��s�����E����]7���}��1�I���B����O�~~/�:�=�MB�$`��bBj�]��͌e5�����W�e�Qv����#щ �"�0ݦ�RD�c4�T�1���K�wo,�cůa/�t��q�IG��р�(�hf ��o��� J*�Kq?yxێ3�T�� ��;��|�^��`���������jk�=}��Z��PJ�N���xL�L����4�io=�l�!���}�(�I($�c����k���랻E����U�ʰՑ�p��\˲OT���w����H�7�W΃�K�$d0����=���g���5� �K�|V��1�x{���\�r�c#�3���"<:��l�Y&q{�R|��Z���fHD�>qן0���dF���ik�AN��Y��X���pG�N�j��gF��J�-�c���V)��86h����Z8]������9��;U���1M�x��y�髼8o��T6�@����'�]�y��� ���"�a������cĢ��O������ �hj�Φ�kE���{�qm�ƈ�hC�� �$�#�N�����5 �'��_"`dSӜi�$���6�8`��� j|Rx��s���MPK%E?
p+5�������o���K[F��u&~�V����=�(��d51��>M �u� OJ�Ty⯏�-lŊ-ϒkf��/����%��9����u���Ca�q+D�/w/���%o�)����s��д�/�}�Vj�+�W�y��U|X������К�.`����2�@g��eC�d�<���]!G<�&�X�21b������%���1��g���fޛ��1V0 �}���Qu�ś�G�G�N��=��D���&��Ҫ���b�s�z�N���"�� ����}(~1MLԐr�g�x<Z�;��An��xe
��K '�.H�O���g��^A�����K�=]i�o%Np
�Q)>��i،�>Fql�H��?O0BZ��Xw��Ce�pKԩ�-s)���&lJ#	:���do6����T
O����S��F� ���=��o�f�|���aJ����	���K��\}�dc*�8��e{�=�ɮʫ��{?,�Q�~Ȕ"s�������qX��_����{��|6�<�maq^����?��*D	�P��D룺x�E�#���1s�)����Q �ް�R�g�/�����H���J��Y��G�@{�ܐ��k�
+��P�s?�oE���N�����~A7H`�#{�_���F����!��u�gq%�,y�Y4A/���9aNI�|�i��s�JA	0?��%�O��a��t��ȥ���]�����q�B�۽�5\F�įu潣��!��п��5r�JK��ہ7�ѣS9�rڛʛ��d1���VkJ}�~����H88�L�o.����CO3���h����Xþ�t�z��W�FNգN����̖R<��ר:�	�������b�]��b�ļ�Q�&���W���ؑLш��O$>�3{T�Ҷ�(.�O����8���%3M��]SLg�b(Ư#��Ώ��WL�߼vx��uh=�,G���O��������:atM��4Y���[~5��P�Ll{+/����)� �%��(�&ڤ&ЦO�x������MX#���.C��<���8&�5=��Ҍ��
_V��������U+���dns�P
�]4ϳ��\�siI�IW2Wv�x��`t���/N�8�g�yM�:�Ԏ��Mf�ƥZ�_�������Ea]�h�d�	c��V�g�nH�?O��x�'���ww\.++)CE����`��s�&���q�9��_�� �6˽�����\�G�pԿ���o�U�.iF���*Z�Y���ѫ�=� $E��:Ţ��d ~$�4�t7��?� "���َ�x�" ����ukv�Qrs�r�K���	����~�}u|?/!g�.9��*2��8��֡�v��(�����1M�w���+X��ڛ�q�BR�S��r��=y�B�����d4/��-��o�uKĈ����v�,��6�ȏ@usƜͥ���ZC�|Xi�h������� ���g����w)rW�q D��|�)E��>���-���q�,3�`.(Ќw*����[��c�2V����~������Fo^��'[�� ��䢌�wU�`��u�a�M��P+�a�>�r��rjB��"��Q, ʃ�E�4��l%l(Ur�^R����=|�kZQ���KjG���L���V!Φ�KUdS�㍣-��ȪY�j���U�τ��R�?Cx������b��N�*��U�����R%��!���N~Ik�����HJ���&�C�(F�x:��.���f�PJDV崲�\���~�-��tKxP(Y�S���U��!�m�d5��3�DŤ��L���J���2��Obkl~m��	C C��K��Cb�&��Sˬ2�Qg�c`����u����zߣel�U��38�k)+��4%I�2�2��X'�"E�;?8� �jY����pz�QɧĤK/�ոlۂ�i�Z(PW�y�����QD*�
pؖ�n���b%u�3/'�&h��^Ӊ���t��:�ʹ\���ֵÄJt��F��+qN���#aJ�������F��[����dH�@md���?��l~�X��ϫ�����޹�5U!,H6f��0W.����P��\M�%��C�g%�ښl�
n�z�3�u8L��4��L\�7`��l�8�a�yP��z�Zs=��C��փya&�e�a�8;/���fR������,�G*/#��Z(J)�_���oJ��;��t��~�Z��sa �OP� ��'���r��C��_ٓK,�V6���B`Š���"�"m�=�Yr �-E�(��(�����U�?��T�)��� @�zo�/i�*&�\U
���-�tX�Vp�����-�P�:�# ��HLE# ���`9:q�,� e31�o&U���4�*t��G�!���$&�|w�H���6��UM4ad�;_Aer��pw�,�Խ�����T���v5ꏵ�����猤m���.W
��Xl�ݮ�S�'�6 ?�æ�V޸��Z��D�ʤT�� F�8Y��C�6�!t,�Ѱ���q�������HT�����d�%�f�3~�ix���MC�IY�٭؄�R䝅�H�ݙh�K4���),"0��?��Hu����ߢ5�����?���$�W7�RuU-�����z���k�v M{�ml|6���(�"ig�q������� �%:U�d��4՗�d�=��>a�Y��C�2Ě ��kġ��s$���U��}�U��dl��N��ߣA(�2� h����o��{ �_Ă��Ӎ5�5�˵|N��\J�Z O*�C�I��V�MF�fO���WBF��*��k
�[�k�9���E��!�-�1���C쒣�i���O߫�v/A^Pp�$$@��U�����S�S@�E̿��󘗽�	1���'0��d���T��`3i�m ����N�3{Q�����P��Io|�]M��s+u?�h��⑑�3
�R�-��E��� V������5M��3X��A<*��З��*^ ��l*�~�1rHuN���O���u+�c5�[&������	��B\)���9	�������}Q���O�������0�9ӧUcgr�����X9�q^gZ�؞e� ��BL�Nv
������h�i�� ��>m/gY�⭙9��=�Q}�= v�cAt���W�>������i#�"Z)���Ŕ����ߔ�]������!���E�`��r*��?q'�#��셪����rf�e7��y�}�֝���b�tl�8E� �3�}ܡ�UWA-����O�����O�p\vp�� ���{&bH��JG&��Z�Aj(��������HO�*0w$��4ϞP�_�m<�HS۱�9f���Y�p�JH�c���������es4���R���k����#~��i�<�Ws��� "���u��Ph��"��W�H�X}�X:ȸ����q~������2 ��tͳ����
�0F!>R����s8s�� ��3�$�:!^���"��8�N��?�E�(���.Idw�r�أ3�-#'(? 5���ګ�B� �v����F.l��<��4�1���r��	�@_���U������g���#ף�D�Ȱ���}���N�\s���j�0iE?�$S�r�ⓨi�iȝY��__���L���.��g<���f���f4�����P����3��؏�g\�$��;Ք�P!�d��&k��v�4.��C���Op&�t����N/�����qΉƠN#�+QC�o��&�~�hz�¹<�)�+����Q�أ|!�g�S���x_ �1���\�s�O3����7"NI��6���N)gK��m�-\�zI�*��n�?��]���<$�.�j�NE���7;��Ak���[�æ���e�܍^�f�y"uMS �DA��V�
���β�АQ��ֱ���*Nݚ�#���;�ȅ1>S�L�4�["�W+.\�z�M!�筥����,D��|��;��L �0i��Cb2��L�UDB5��2����K_��m<lR�W��	�A�9}��!O_�/�R`�,�x��^$J.���zb_ksp�~�SF�'N����
�����|zFb~LE>>�^(�Ȕ;*�s����q6��r�֔Kk:ʛ[����&���3����մ�k�Dʱ�Ieg.�T�c,��Ϲ����_�1��gO^ţ��⑱�}|J�o7�p�K����eA��Y�B��W;f)A��-_%����L����[3zȇ2btQ�G^5#D�E�awV7�W�6y���K;4=_�Z9	ݬhyd�T
.a�m`��#-�o�녬��q�U݊f��e5@�*��ˌiu�͖�H��r���8vT7CC(�=X=��(�u�,���g�G��K3:��^��8��9�gKL��~��^3�����P�* �K5�8@r�=�;��Z�u}�f�?��.��΄.+y�X=)}�f����H	���:�ѡM���+�!X6���g!(z���v�5G�?Pr.�n[�Bc��4�Az$)J4��R�F�C�C�FhsI������! S�ɕ&���a�k�z~/!���G&O�8�v�#�>������?=�d��@��o!����n	���Z�o��`IF�c\}2胤�ʲ�9��٘�P4�s7#��V�YLѵ�q��H*��n&����_�2O��6��0�����(�g|v�����c\�3�Vu�t���~�N4�~���WK �alx��s�]DEP`K �;pu8��z2�C����ֹ�Q��kol�����x�Q?��E�;�d��ZR|�ذ���p��*��*$�gD��6�Xt6�z?��:��5�*x�qf���m���	��&���H+y�Nϝ�+��e�Q�/�kY	[Մl?6?x��ba�;Y�4�+!&<�A��}�����^ b����5�$	[�o����>��� �[��'J�,��A?b���Yc}J�%����pVCLQT���1����V��
μ�A*�b�1GR)V�2���L�w��i�g�]�� :)\w���p5������g0c놖�*Ԍ����� \FF$�x�}�����l��Qh�Zc�+�X9/"o�-���silO_����2�kK@f0��7i.?nO	.�FA���
me�8�z��mg�=��T��r:�.B^�]�ytpq��q����4�t������
��P���d"�#���1h��
v���׭ެ&�v3!�޶R���鬌zҿM���H JN7j����6)7}�qvQuP�;��U�X��5�C5�W�.L�l��Z$u��/*���ol��6 �Do��f�Z��9n���dn�t ��E9q�άmac�]>'k��u�W���lށV�.�����A�d�<��n��cD7PXJCK�C��G���c�:T�f�;4�t� �W���� !�ܔ{ḼɱS�rJR��N��rX���z�K��B��y����8)�f�U��%��.1A~���ґW�7#L�[���:�¯���A%$he�����NK��~Zi�.9���J�����eU���\�M ��C��T��� &Is:�cJp�̅��.�x�f}	�zQ�~J��S٭����*�6�	pe��$��;7�7�F�)�r��ľ�t0#�e�
��@����V��'���FB��� ;}u���N�*��l�(��8պT?���}��ƭ��Y�Sȹ���9��Y���j�����m}���*��I��d��B=H��eP�y�+Z�ǭ�;��!2�������Y���G��v�'�w��H�4�0��:-%�0�����1|�Z�Y~�{�B.w����8����Hp�eVW��|�M7vѯł�B2ygVU��t��*p6-U��B�3��1:���Ĉ?�?U���6��%���ѹ��7��>��/yݐ��8��>W���z���k�R{�?5��=��  d��p���p+�;�|��1b�f�J�}��eО|�Q"��Oq�R�Q�3��
��_t�;����1Í�oLz:e�t����p+ap�\�F���m�2�>�P����j���K��7��]Y$O�3L�N8ٖǮ��d�{F�CV�-d���b��`˰�Z���������sے$�:�P�� a��O_��*DV�kWlŐ��/i���g����g�~���͂9�zk$йī�@g&��������������p�\M�b��0��@^qK���/X��0�v�,n9��<>'
��QȢ�m��<3Ȱrv	�M�p�w�R0�ͳV��|n��^B+T����/,����&�\�dⲵ�A]�ʧx�G/%�nf.H����c�&\�@[�Nb�K���rY����Ҥ�.^�d���_GWUxR���GW�n���u�����ğ =�����@Wq]�D�,ss��u|�T�����a�c���j(��3 ��<�5ؓ������b��[���q�v��>G�P9���,�z�V����gX�`��_��m]z�(�ό�ݣ��Ꞟ���73�᪽~�`�?�;�b�6=+[�} \��5�avJ
5k����w� m�L�����졵��͒v��u�8��Y>9�[ę\Ӵb���,���F���]v��{S���v�����f��F��S��,[q�×��0QU�;��/:G0��Y?&b��aZ{rdb0�>6F�|�����^|�p"w�Pm���ß
̭��,,-��n�e?Q�1�;�`�XC,w��&��aN��m����툉�M��uG��u5k��A��S�=�ԇ��8�G};f*��=��c�9�3E{�z���8x�}Wd��S����RYE���9j�\��D�����߷�鑂\��`�X��d?�ɩ�<�g�z�(���ݝ�tuPWmT�+�>G
�b�5�>��{-��_H�<΀�*���;�5��0���c�D7·Ӏ#�|dx�yh�� ����a2��_U�����D�l���G�����>�}��nKr�\�������)� B��{��wd�O2)�}�~�]�����E�#�#7ɥc��a�R�q4��5ɠ0�HւI��s�E�L��M�{>泎��[����z�E�E�GI��\�1�j�JD47�����xR H`�i�-�^&� ֨�Rq��fJr�� *O��`ɖ��od[&��4=�h����Q��Z��!;��i�v �*���J8�kqt߯_�fkN�ZWVBt�K�RK
�`��%�����mH�s����Fy����I�1��昵���W�s[9���d,
�6������x��e�a�mK��:P�$��2BKu�4���+���,u
�iͶ�*��F���&�8����)�Z�K�+��z]WH�tC�����ێ�!7OI'��_�z��P�zd-��F�%)�ǹ�����;�*�f���:�Z<���xi<���ۥn��xG�vE�bm�In����Fզ�T$L�����Gd�����l�<3xAgc�LA��ҠAs<l1B�9M�,vm�1IJ���l<�
�t��@t�h}U��ZN N�ީ!��v�	ܾ����BRHsKM��T`��NW*���Q
�hsl˭�#z�=�[�V��R�0m�Uf�֒4��d-�λ&Q�=�����)��J�]�h����K�d���3���.[��
(���o�T+��
�J���Ǧ"�e�z�M�.�_M^\�>�nئ��?/nsw>RWo^�����U8�hu	�ۘES)�[��ʻ7�_n�{{��iቛwK��8Y��Y{ߵ���o�ؤ��ѵ��@L��/L3=�L�s�(�5I��&���cǁYgB��� �d�{��Jum�R|�Q	���!Y�0�3����|O������_zkC.���yq�Td8Nz=�-���?�n>�! �������_�VB0�E�1�v\�â^9=���|缏�bYk^�����ô��^�&��oO.�� D�FSN\3��c��rx�M~��=�R�Q�U��H($N���yRxv��4y}���|���Q6|=~�4�m�O/��QF2���6/r��ݧH�	�bT�����OQ'y��n./_�jd�W�G�`���F~��F����^{��2|aQKc�H!��� jǋHG,(O�y(��෽�?o�ɒ�7�:�9��Yw��}-n��#b_�t+-c秡����8��f5�'�ֆJ<���EN5O���B����hV�wK��-2p,�{�RP��z6�]�>� �y2�Ց�N�R
u*L}�}�pCc��s��z��z&D��wT��[����崕�s�m��#�6��%o��Z�#2��%������=!��O)N�
)8��&�ɠ��S�?��*9zA@/`��YdǱ�ML=��h��������Od\0����.A[8
s�'�w7pV~`rmJ�+�+�4�  sSt@ ���xYD=���"[��o�O��j r�����ZJ�r�}C7b� ���N9�D�ٔF�s�Es��S{�������N'g+g��3�cP�YA8%�(Ǿ�W9�+8~xח#B��5�)�U�yV�H�'֚"_to�L�����DD��j2��E�l�ֈ����=dS�*�̦����>�Q(����D��<.v�]��K�l+���� [�m9��if�%�^+�#VZM��^��k1O��*փ�>�m���B���W���Đ<H��l���/|�gR�-�`uT���b��p��qkcG�n�M��m��=��,���[-ջXaך�D�v��)�.֩ꁴ�R��D��nٶq4`��!��X0iqQ��"b���t?�6ƞ�=��� �+{��{�#�Uw_�)֮$�7.M���޺`��Pu����LT�`��.��|�E�m��~Ĉ����pI�Z�y� f��?,$��9�D��+�o�:2�)��G���Fiό����ϱi� ]�}��	*JʄT�2�)}�}��	��	�Y�>nDK��|֋��~�س�Tl�65)q�P�ۑ��pq�>��wC�W �J�H�Ob�\辉�S���p�d��d�~+�4м֙�2_F^c������ڳE����u��L�>n`�u�ξ��o9�Pu����s]OD&��j�!?���<ų��Thd�+�ήo��v�*�18���C# ;$"9��[�ʖ$wS����T���9|O�C�0�F�5����'&����pGI�OUb[
C�]i�����\c)ot���ȹW��ʣ'��� +�֞���E_���7l�Q�f��ڽ�-[�Tu���.�D�M�� &D�i����3�8�4�� ������o<�b�k��N�U�a(j�C~얳�Y{hk7h9��~�6"��5HR*e�
�u���دRm����:ʏ�;a6A(hb���JِqpR�g���T�w��c�ɹ�҄�4:��E���>���N�I��%iI�y��-�0'�=�l���vE�klF�U�'o���5w>����a��x&���4���A�I��CZd�O�!�Gm�4�ɳK��RZ0���P+�q��G�	o�%孷]}@uM�4ˑ���ؽ����T-������6z�q?]���I�;_qNT����:��ο�}�wN^z�*~�-��0��el����>�*TAf��m�Wp[���!�K~����D' 8��.��br4�����\J�z�^|�*� �%;h_����s���Y�gj��GD�X����$�Ʃ�q�H��Љm��^�,�� M���|˟ٌ��N$	�%W��1�lǯ�����������tM��I� ��Ǔg^�j�$��5m��2��W~H��Dn=�Swvoj�=O�-8�gq1�������Tت�1]�ƛ��T�������aG,~��e�."�h`sZ�:�с�gk���T?����g�����i��,�pJz���@X$�A+%=}�*b�_��NX��(�wl���?4���?Izk�G�ql�	؉h�=�2u�D� i,Ɣt@���"�j~�Q��@el���1����!��^_|���;L��Q"�z&@6^���.r�-��O������v�c�qՋt� 9s��@r��e����Ƹ>+�p	�NZE�P�_Qe�QԦ�z/ש���0������N��W�q�
��P3���(�Կ�Z�ޭ�t��o�h������RFՙ�V�a��w�ÿ[��|;���tyV1�����[�{���3�~�ƭL��Y(�ޅ��.�,�Z��^����_�G*��
��s���Mz=�`/��P�3�JM���*�-:R�g=��8W��nV��@'HgS��;!0�-D;��n
+ۮ�℅���<���>J���!a%�URX��e��!�.I�
 /�K�k��8S���n�zA�.g��ޣB�U����,o��m7Լ�T*�ѦW&! lPhχ����f} ���i�g�^����ȱЫ|b���*�Hx�o˨�	�wa���j�דm8���J��9�E�{�V�F$A-�������yp3� ���Q��2IV�N(���S���0?1��yCB;J�X�^�Z{F�~�@oɃu���L@�����E,�%IE]ا���Հ�Ű�4d���*��n��`������e���C��xbU��l�5��_B(g3F%&�� uR�h� J�?��g�@����O�?�Y�PL�4����Цgیa�)e�1v�(Mx� �o�8w�Sc�K&�Eߐ� �(�T��
��r�6b��v���t����e �p�I��`u��1n��l���h`�U��|�(�	?�w�Q��w�֔$UA��#��\�+ٲ7z�]C��W`l����!����c�wp1�����"p�if�}�[^���m���|F��Ur��*2��_�g聢�/Dm�č�;�G��>4��5�@��JH@�C��s6�!g�h��f��zF!� �Z�1�p񅃫W�OΧMÀ0�D,�1�L��Dt��u�'�_G؅ܼ���F��T��E=hdFv��kk����klQ��mC6n�e2��Կ�0"�+����(�ՆZ�xP�g=#,�н!�^�R����!���Y��=�c���jÂ�sܯT/����Y��.q��+�.�~3��r��T�(�b��P��6����P�سwNK��d}:A��ؤ�x�j��)��/eD���$]�4�J���FZ�:��8���j��yʝXJh8�<�)-��aA�nO`7[�kf� ����]�ah�WS�r�U�b�cd㫘A���@���wCM��p�@NL*=�5�g�Y�G�^�S��ϓ���z@�)�<�0�%��ɵJ�!���2�ߺ?�8cZŒ�Ӵ��G'�;�M!$Pg�	;>��0�\�NɲD��`����"T�f����Y���2˙��f�݉�q�P�RШ�;tq$s�
����ݔ(Q���Н����* �ܭ-?`���6����1�a�D��:��j�(��� �nWȼ�GP�����J�Z,HS|�������!��t8�_I ����m�x-M&�?�m������Z�n?�W�x̝�'�I� ��Er���v����(����R�	��=��Ϲ0�(�so#"> ���Zר��7Ց.�����nyQ�V�ĭ�x�Sè�ol�!F��ԋŴg�D�z���݂��p]��"�gW!�x">�IM��~��h��"QEC�IG�uΚnV��	���O�m�mB�yX���c�'��֠l.�8�A;ᔻi�1�V;��� i+�648	�zR%��0�xD
<�A�����g;}.�cb���QY\T��ۨ�+�N����8���ٯ�J����.0%%��^���u=�AZ���(�����Hf� 0}�/��1K;ZF�R�D��v#�@Ϝ9���������cD�M1�:~B�D0R,��29��@w���ڔEmwz� M��>�6�M{��L�i�+`ِZ�l�΃t��ȾV�I}���2��b�\� <�44��ֳ�A�nq���lH��T�Ӎk'vo�8�u $��v�l�k>�{�w04��KЙ�����7�	w�cz�E��Z�b~A@�#����<��sڰ�ހ��,� ���8t��[��T�o�b���+,�y,t�@˂:��ZK(�!�[4��t/cq�K�ѲC�t��]P��ʠ�NM����4��Fmn�xL?�z�����s���YC<T�p5�*�+��-�r�eV��]�
/.�њ#1������1)9�����r%�Ϩ�DG�;���r�x�Æ��U����9W�$#&:�����"P�.���ҫ�*�ξ>j��AL%�#^r�YW$��
?	�?��Q∔�+�Y��,i;m���Y8?���9��6_���֬R�����<��k")f�n���FB��G���x�I���
�6�&7]+ !���z�e�F��ĉ5��-��?�_��L�M�������XuG"698��{�~��l�I�w$u�:H�*�����I�zK�Yw�;�:ۧ��Q�,����bҢ��mG����.����T=j���U�*�~�?� �ʝ�c]r'�/��<l��0W5Թx��C��,n>�ޚ���l^�8x#j�_#�5�B?���~�P��{ɁR�x����R��j[<�/���R~I�K\�ͬ�����6�.�f�{Xz"��{o�8tq��u�������i���|�(���m�^�p�DP�ky*)8�)}�z�g;)�c�����L�%Rz�%�%&�S��.�\����N�,�j����� �����z'�%�zW20a�c�6�s񩚧���)ھQ����moz��9#����w�����.$�9��M>JT���N�Z���:ozW���Қ�݊(�&���)�BE������2�-�����#�Q������j�V�J���͕����Q·��Lwno�Vѐ��<<��?;�bm�bg�bH�b6dw�N>�����b��xo&��M6���Uj<Q��� e��i��m�6���wm��jf/W�e�e�SNg�;S!�9)����^��S�Ju������E�6��'&VȊe�JOt��_#�T4�&�(E��e��-SXR�Q�g��~�����-ƭb�*�Cn\@��]n���^��S
�ᕢ�Ӹ'ho����<^	3��3���a�],��!A��劑�׵&B�\��5��:xc�i)s��T&�K�ev�͵���r0��ζ��[�^�Y��9�~]c������ە����c�Ep������t�칤.�7B�QЯ�d,P��c�c/\V�j�n�'��!m���ɺq��I�C�Ey�ح�:��;(c��h���گ�	��^��$�}���Xb������ 1��s\��[��Y�K�w?e���ē���6,�v��7T?�2f$uR�K��6`N|��g�5Ml�~��h�Z{��A/?n����x�R�������#�؆���YAl�Ӟ��e���\�ڣ6<�E��a0e(5�L�토�����U��K�
�1sK�z!�V=���i�5J�W\A�Y�qE�hA]�%P��QњC����l���.���ZA��	�]Z�8���g�3��{�R��Ⱗ���
w���sh�}_�k���qeA}s��B��T��������#�,�����rKJ*��}a6S�x_�R�y^�A4B�`�
�g�����a*{ejAfB�u���m��UX�\���E"�d�m�7f�$��<�̫�oQ�B?^�K������[���GXNuᏱ�H���D�O�0l�Y�v	�\�n����I�ѵ�b9OQ&���k�A@��`ry�xe�P�A����i�����%�@ZQ��FR�4fP$��[�d ���7���fb`��s�|B�d��F��h�3��c�[5����"�d�g�y��Ym�sgK�V����d��̳\R�U7L099���NB�la�Xf!�?�u����ᅶ��}K���~�à�/�B�-�'Ū�m�������p��n�]�U3��x�ӿk|1@<�xY�8h�sps�7	�')�6�b���=�������NY��"��*�cȊi�H�8'��"zS��0N?C��y^��U9i��y�
��HK�zCzW�Yz�<��s�
`X:9�4E0|]pD��5�Y�nt��ײ�N�Z���>�ky����_�>���������;�u���Vz<���~��A�_�.���8\M��9�*�)���F$it�g���ܐ�覰83�^|]>)�
㋴Lg�I������ܖ~�{;�ɸw�=��J9R�]8�a��츬ǧ�,0���0�;l���ݎyy�p��<���v(7&��60��8B��P@�3]�3��xTZYo�W؇&��
���Jvo���9+vV�`PH���F�hS�=lR)W�*�]_��� ZBl�|���M��[Q�*��a�͋��v�x��ޘ6��E� 'b��H�~
}A��zk[B�W�9M�������P7�
r[D�4��I����)nߦ�ܕ �j3�s�w^�������{vc�hb�����Lk���р-�m��A��' 禃�	؂`��;���|�ٱ~�E����`Hh]Dy�W8���23�bHHvf8,���j����R#�N>�ч�ޫU籝>)��[E��0�A��;���d���8������WC	�0�%��Onz���?L>����%+õ��P��!�Ҵ�7�0ʺ�&���1��x���[����o؀E��%'��.�4�s����>Ki�u~��"|U�S����|�c1{�����H����)��Oؼ�D8T� ̤'oL]݊�qL.��ݫ��E���v(�E�9���~����9:�*�5E��w��ۭE{�F���U�'Lq���H��ى.'d�G&�s�R�(�(Jԋ�sh;%��GnYRP�T�f ��'%�C�,Ŋ-a.����L@T�E�5����k>��%\�Z��L=�^3��@�u�&0Kk퐟���+��^����lj�߼�P������O��owȆ9֯v�}���@1'�$�e �٥� H��1��te�Υl_E��lW�A��N��}�[�Q��
-�Gq:�u�/���x*P�-j�q���/�G	sɐ�_�\W����[�fM�#nW���[�����I��R�Ò��Nu�+�s��vq�95��A<��Y����{�)~��d�0T�GH�*�a�5�0r7�lQ&H�\Q�wG�3e�*O���7�-W��X�+��x�x �B���yNQTD��!ˁ�j�5�c��ң�{��`�-���Y���J_� �z���3+�LPQ��n�].����Ɗr]ӜCQ�a����'�b;A�J�ѥ)ԁWj���*_��Q��#i>�_�>d�Y�^�KwEU��p5)�F9��]��*Y�x�����Z�"8�`������;(����3�WE�x]��l)la��`�$�����>,ƍ?Q�c/�}�`hQMLѱJ;j<�[~���},�!K�����um���#!0���Wz|#s^O�ḊR�$��8?��ٻ�m�t��YḜ�;D|���� bH����-�k
R/��(�~qfoF2�9��g��a(8�#���48;�{²�("�g@�E��pn�]u����,�F�9bˬP_=f��K������ �I��'��$[�d<л��wV���������K�
��ņ�d{(�8c� M<��=���
�|n5��W���G6P/��5�NT�DիVJ���hش:j ɬ�sz�MN`m$])Dc��;ӀJpFF� ��=�x��A���W���X�I=��A�(]���*���c��H��>Bc[����w��ي��\f���������_z�G��!K�����5pq4�}�_�3�]iڟ>�	��E)�M5��Vb��Ś R��:��TȪQ�濿�(����]OxԎO�K��Ҩ1erY���1��9����ns�
�z�I�;��3h4ͳo��DЧ .z^�` �g�m�K�~m�����A���ecεKyZu�E�HD9�wK)3�j��o@��(e��9�*����5���rc_Eu,�n�9�YW����1��<kP'�������T3��~���O��U���� 1]=��*�@��/��H�9Yx[j�tn���	S�!h�7�*���v,�e���r�S�A)7�ݛzzז�j��5�7cŻ��*!�s�1��B����߬�7s��ct����m��`��������|��hk�_TA�}4$��hʌq=��ף�L���Z�]¹N�����-F����zG��:\��4�����h�������d���D+��Y��%1^�#G�9������+����j���w׹¥.s݉����y`���p2�Q�H�%[�.M�8&�ߔ��(F.�z���G+hR>OM��;Q�z�ŻF1�����(s���L�W���`'�2F��8���V#����0!�vV��u����5�s
�l�<�a>�8��9�`�U[���7�����6��*|FK�,��Aoq1�TZވ����I��Ѱh&_( i�KR��j��T�����s>����|u��H� �_�%�Л:Ѝ\W��\�U��bdį,w�K�g�/s���n}��s��7��9�SO��!f��#c ��HP�ֺ	���H)����E��\�����G�͵��:�>����#F�In��`�jh����NT��Pby���}�w���MZ�QE���+�����i��ը�K��0��%��DV��D��_7�9��P�K;��팁�,�O����/���Ƒ�x�I��[f�Z�)���=�,=y�>��l}��9�D0���nM	|�"��r�G���NZ��<('��%�i����P:���?�3������c�L�w�/����o�<5����{)�����+:N\�a��*w��E��>F���.c�A�I�&�A��h�������=��*����X��@�	�BQF��D���KJ�3hBdKv\ �<_�"�o���q� �^��#^��H�Z�Gb�1[�Ќa���f�b0v�����p�>'��MV�:pLm�9	��a��A�՜|	_M{p�זdIW3�b.Y�/\�wC��� ��⠵�pd]|F���h�x�KW�y��D	�0-��%nxT�9w ��9X�\ÂF�O@�[(����k��t�]}��uu��3��B~7X�6E���T��}.�q��K��W����$C��WK��G�T��&As��I��&A���O6� mJ;�s,��J���c1��܍��T}HD��;���ဍt%���+w�(g�cG��\�݅z��ɨ���DE�G�R���7N�rZ���}�[���'���&_�г\��$�߷���1�3��}h�T],�B)�i�����Κ�>O�]�=�#P\V3�����Sh;S-�1�bK־{�͔x1�[���Ju���,�N2U�E��m�w�UН/��w=O��g��j��P�����MP��HM"8� �'V5���;��5�OX�*�`��@�#!��a���B�X������S^���;�R����(���S��E���^*��]1�>��l$�_*�JQ�dj� ��S:T�Q���O��6-� �9<ݧ3P�$N������fI�'�����n��[�}�-�#��t�;�4GAz�;	��Ț��8	���q&��m߇cl���8F,���|.U�/=o���cU���F$�e躹m̆//p����,�[{����g�`v��>g�J�@I�B��6�0�;�~I �82^�t+�x���Aa%����Y��pom�M�B����\��h�����A?��~���"+����O��6�5�F�@�H�vPVJ��%U_[��\
��h��R1s%�Q�n���0�������1�/��ݸ��z\.�E��6qΖ-�I;�gT��n���e)��JYoO��옡�7�p�����=��}F�nkqbE����Û�'$�%9<9�Z��Z\�u�*{��6�:t[�_?`
��S��.#|ʷ���%e&G.�5����&@qY�c�G��o/�D�a?��"sl��m�4�k05�2��Q)�uy*s�W���ε���F�]�s�F�r`���	q#��y�[Qe���Y��<;��p�^�aU�禰�2�~���2�\���=�p����P�T�����Ƥ�dp���y2(��L�J���;q)Wޗ���D�]���8��A��
�ۜh��p4�2g�>�d�Q�=�rC�ΡFWh��*2������|��/ �����C��VJ���Wl�~@����)"�n���ei 8��Ms�}�JEk7���eQ�b?�	1ώ1�Pv��������m�,V� .r�W���BBqNԷMH[��ݹ��s��gw���cDӻC�����j����e�X8w��b�Bv��3�1B��<}�=f"̤���>=�P�6���[��"�(Pq��h��y�C���'���o�
غU^�`�>���R�&�/�(��r����t��F2<��/,�(N)֨�*%\/)78�U	��y�D�I��BndT
\)]�@�<R�c7~��QP��T���	[3�Iam~�ğ�T�����+��r�_�x^_�ؙVS�yl:�u'�=#5zx�%�d�|ꙧ>�%i,m�&Q����{
ټ�r@�|��`NNe��	�� �f��OVzϕ�
tM	2�/�S��u'k�f�������&꫎��F�ȇ'�ٌ�2��N<���pc���Lz�,�D�J��v��U�zx���ߊ���r��B�o��g�	��@-t�����?qJ����?��ռZ�@^���Ձ�wt�U?�2*Qi=D֋?�p�v�M����1o�\�Sqo�S�q�I���i���r��8�{\G���G@�'�=� �l�	tj�ȫ5����b���5�mBO�J�\�Z�ߧx'��4�9��'x�LS͈I֏'|e�2�G�a'�s�(e5�w�6�h������x����o��_k.�B�H��n��܄��x4B�R3�׸��8��k�"����9f��Y��^����`5#B+I�gqX�;� �і��f�C��2�R�j�*��\��Q�ePjb��D�H�e۟��+��k�Y,\�d���Y��8`/�q���䗢ɠ�-|���ܤ���(�AH�Ac��$���_���t�/y�B&w��fݳgUVWqKs�jq{�-}O%�����5�	U�̩�����GΫ?�{H�qMq:��\C!��]��< ��.r�]j�b�!y)=�� ����xl�}"��Έ�x�U+恀�몦m?8A�$�O��oߘSK��R�N%bu0�����b�@_k�m��>D�?[0�{n�4���,Pc���l��f�p͵��-N����B~�j��Ň<��zrL�7��-^�Mf�6�j�K��5�(#s4��+��_ p�D���׶mE�ϥ'v�P$y+	�F����m����OS"��Do����o� ���f���u�JiaY�.k���}�AZ���WBg��\��h諉�,�½��4Kj�;�D�1�0UȊ��/��Yz��� �Q�z:��B�\в��Xf?�H�&�5v�	��LP�@kP�	a2K�}ޢ�<;Uau�s5�������A)�H��fΆ۸�ޞ��]�RJ�f������������m��#$�иQ�Gˑ�3Hͭ&��$z��6��!��P�dN�U�ܩǺw��;St�v@��Y�b��c�G��hN�vB���q�o{h@��S&
��	Dn����tO*mA��8������t�Y�W_Z����7���l��+�jr;�i0�ܩ�1J��m���G�W���yo+�]�7�G���tUx���5x.� �Y�,Q��RJ��_2�S�<*�����`}K"xN2�]T��+(0��]��X^`����k�-̙?X�1�CVF�8��R������ ��2�+�(��0*(�4�t�2�@L���y�N��P�TrǞ����̘K��k�a$v�/f�r�Ǽ@����24�ͫ�Su��u������3���ދ�u\ys�M�i؉��+ܵ�ݿ�z�eM�&	q��6��6<�x��v3ӱ"�ʨ�p\���aN��-�?�0W����{�h��� 9d�ɰN͗,�� HӍ6Y���Ț'>b���ܡ{��b��S}�ȮZZǠjOH��)o/V�2Ql9T�2�b���T�����?̻�,k��ʊ�DGY�uK�4��򓧴q���e�p���p��%����-
�F�-ntX$�;A����`Մ��}$-~��x�􇣷ѽH�����@�:h�_I�@v�N���QJ"� ކ^���ӓm��6U�N�BN���
AJ��ǧz��љ�)+�� �F@�"RO���`� ,1��û��w�.-�a��&�5��*E�lܪ��7a�ٷ���kf.���Lձ�ib��7�l� x� 6�E�J^d��Qz���~	�yP���:6P�Ů�>Pj&�����Ʉup\�p5��~�a���W"e�9ݕ�ZE��K��O;�E ��]n%<�q7�i�;l)����;�V���H�	�b-��9���,���؟�������Z�σ�"��IsW���� ,*~n���J���w7Fsg�{ƒ�kۺQ
)S�L�x";�=l22�#bBn���i�yK��B�h!��$�W������ڨs�}�����'D�%x?��Y�\oQj���\��(�=WC��G��M�x�y&D�����&c��|�����V�u+�S�x�r�8N/��@yT������E/\��`�QpS�nO�h��a�"bJ��!ޚ��J7Ż��)r&���l��v��5������;�*0't�z�&��5?�Eu��]F���7����:�$�=ylj�����lD�^Qy9]X�"o��h��䟞��K�H�4Ӫz�JW��vX��/NRm�G}��˦2��K�)�m���]��;g��-�(�8�����fgh
�Z�S�V�H�׳�T^ �}����Վm��	GN�h���7rEi�ӛ
���ΰ��*O[t��*͸����V�������n��ZM��q��'�p�$r�ϸ�-�l�1�%�nL��(�H�NYo�@�Z�ǔ�S����f�^�H���9Td]��R]b��o�PƆ?�k&�B��L���^�C�!��ݦ��&��Lm;g����P� ��D䝏j��Pq�yY�y�k;K� d����Q${��^ ��2�JFf$�2��,��y��g�M�%��bϭ���H����>��x���R8g�jԢ���4� aC���骕���e��5��x��t���V���zU
�Z�χ��t��� c�K�D�o�@lG9�F��NLM�!j4����@mK$4xw��A�ձ`�#� �uh��;��1�� r��9i�e�L�VP�L�����%p?P�)�K�i[�A{�5���vr�OW	$v��r���F��;��w�������H&�# �<�����<�����9A/�ʶ$�]�kQx}��
V-5�P���93n����O3�"����^�������mS(5Sͯ�k)݄ڤݐHhh�,ַ��[/2ea��a��uǈwW
��P#vZ���Ne�82n.��G�F��n;Ѹ5��G��++}�ܣ*�A�Ә`��Y���q��=��)��Ĉ��@��%��3QG�rY���"@}�4Ӆ��2`dh�{���J1i����4�|���E���@N�E-�+�^j
�'�ű���P~9�1Pj�t�1[%OR��Uk����BF��C}y�Q=��X����Q��ɸ�aD��ҜM�߯�Qe����������A�3���2@֌g��\n��0����^u�-xfʑ3d1*�]�kk��>�H�Ac��m��^Uw�?��Pt(mX��To_m���,��'�Dу}]y��5���*����ғV���.R13e�![ݭ�E�ʲ����d66�H���>�#�*m�,U�aL�%�C��G,)���������5��Ɏ�\w�"��V��C���!ܤa*r�T��/q�8B��0�����s��Wc���Z5|2�k�]�OW<�:�4�b�7�9�N��$���Mӭިl1�sɄ�</����`̎�����ə#��sJ�9����&q�X�q�Ϳd�S�N�#��^!0�)���M,!��"�9f��4?T�Ѽ��
�(㩼=�#7��(U��:��%X}�l��{H��6��������WP�b)�Tn���0�Z�/[E�I=�d��J��e�LM\#p�煞�~-8$h���eJ7l[fM����^�W�g�l<��W����yǈ�`?�� N��9ɵ�m��b�ނ�a��sVY���A?D]�EAԅ�yI�ۂ��&��g~����{M¢��?��0���OEbX&��Y�̫$j��>�~%�Q�Y�b~" 	c�3E����� ���3����!��xC�zq��S� =���:$7��jlJ��S� =���*��c��Kă8�,�S0�6SlIW�� 
�}Q�|}D�� jB{븱�U�Z �ƍM�9�ȳbg?�!Ź��;�%���I�#V�R��`]�K �=�x��r/#��
�������qRU�I�+Gv����X�{�&?U7��F37x�W�0]�ul����I�R�PMĥ�u�ڈ���-�˿�R*��Å���B���r{ *bsz3Z�ߤhAS��H�1HX����~T�B����]���Or�'\�i�C�A��-�=����Úw��0������ �u��� ?Z֙>O cY�!�ġ�7����_��z<8z�༜�-eq�t�<O�dzo��#�wC�+�ǲ�1��pϾЛQD ��>�Ql��<4{@�L?�F��*@ xI}�dH���3oX��f3����G	,U�/��h�Йp�l�[̸��c��BѷQ~���'���J� ��vf������=z�fY���2��P�4�u؟|�FnGt����7���ߟNG�P�����Kv�}=���O�C��C�B$��(�Ɯgo�h�4��uk���ͦ���K����m��-Z�e�\�"��t%f���E��1'�;o#��g��<}Z�)"Ҕ�MgE,�=��r(vr���W�tE:���#݋;l|�7���Ҧ۴��믆�H����r|pw�W_$�<����Q�p�Kg�j���f����~��RDmU|p�~1��e��+N",��^�iVU�s6�Y}��QI�TCC~��� ��[*s���G��t�%��3�������2�����6mڼ)������ԯ�H8��ZX���Ӕ"W�}�E�4_��z�+.CM��� ʎd�k��[��	��ަeE`88$�Z��;fAgGDl�ALN씶$�`Ge�ʈ�{X�PvRG`$QyHҾ�|{�$�(�H}X��^s��>2t�z��I�Mpϱ ���
CKF�2Mo��`�����쩚��<yZ�AuG��s�H��e��m&4�~7v��DMloy\P�C��(�:�n�Pp-.h��^=�_���]���㺛�M�8b\�[l6���<s�zu�N�ޒc�S݀3&�~����\�Wq�u�(㑝��+r(���<�wLS��1���������M�h��ouM��1���5�8?�;Kc�߳گ���N���1�]+(ߟ ��k~���c�-��y�R|{��Ob ���4�n릕M�w�FyI���h5�z�(Z.��_mK�7�?>Dn�5
�~	�=�>�z.�
�F�<Hv!L�B�O�X�ʁ;C�1:��ܮ^3(���)2]�2��E��fqݽ75H�٘�yY�&/��RJ�'��՜��������-7�Kפ�۽�����Y}%RI�دvhQ�2��d��.��l���}��{zO.��:շs�F!�^�xv�����g~Ԉb�\<k�l�[�׭�q�X�h�X/�.[�Z�a��B>��#I3��l�������U����s���F,$FH�9��6��%�n��?SH��i2��������������iP���l
E;?����W9�2��h�?p\��ZC#�{v�W36w� ñ�0�w����ܴ�����
�}��7TNw,2օ���t�Ք X�"GT_RBAEmn��`o��� Ua,�����ocS���X?+]`�<h[�҃�j�Ĵ��$)-�HV2ӳ�F����g{{fbCC̈�z�H^�Gm�D�xMQ��plӰ�[x�3T��!)��Pq�? ���c�Y�)�07�b[��x��,�d���7v��lCU����?>�J��*��ĥ�������j��;-ۤ��P����������	ؙ��<N��^�X�݃�BV�H�@Au�x[�����q)�o��:K���N�<�6��pG��+�����2���3(��dj�GR��n��NH�(�.άǀF�(�5N�3߱m0�ӻ�$d��,X7nPL�TU
�|9�G$���L���NhG~�� !"h<��EUI���
(~;�Lg��\�r�v)����)f�	N�����~"�6�B�(�~�f�Gz�ɞ��J�u�ႇ��Q4�0f?�:��iJQŰ"���(^�4��}�@Ƙ��w�p��"B(UW�2����֚,��O}�@A���n|>5q_H��ç���A�_�n�5 ��;a�Y �Y�6 �Zw(<��˧R� �&;�Pگ�8D�#�n��M���A�D=S�g^��x���a��l��ʹ�7v�W�$}׃q+���y�#�{�ff�(" O�6��T���u��	���
^]��p��XC\�x�moP���o%JLDP�\m�s��"L�S�l��Շλ�Fή䀊S�C��O���p.��ri�l�H���q��*����D�+iy\w���_�!��Aʟ��'�5DG�� �b�fU|��%�M]��1�6	x_��E�af�c�ϖ�)��O����qyl��Z/bHf
���*�w��A��=Q�[s�&�~6'�i��H1"�I-��W$%�4������'sݢ*�ڹ]�����-j{��UL:���?$th��.��Oҝ�����'I~�Wq1�n����Bږo��Ӻ �P�T���50$4�~k���^��!#��ĭ��i�74}3Awd�85�0ހrG���U+�>�,�"{�$lc���4��������ɓJ�/��T�������^UaC`�l�i��x))����5MY]�ASI���*��42P$%5fwaX��M���Al����G�����E�`E�(M4%�zc�V��^����9k/�	�{�X�pd�ɫ�����OƉ�\`vt2P����2e�3dJ[����}ܓE���>�������n��?f飓�K�
�
J��_I=����I4W�5�(�أ��3F���O]Ҩ2��F� �D<�V[��Z�a$I5���2�`B�e�~�1������S�'��p.w	Wz��z�8�G�� v�t~�2��W~YZ:���&:��5�!����x�?��0bo��Ez�Q-�C�G̷vN}C�"�E�2�|ge��Wت-/�Z��楒%�DQ]���|�n�"�~�_��{�:����b�%g���0�Ќ�$$�3�#��=��E�����ꗚL���`�����cR"�� �x�X�u�������.��l�V��e����٣k�tv4���*��8y��8I��J�Љ�#�D��O�\бѫ�8b~#��y��c��Ҳ?P���l��O�b����8pK��_��G�} ��oC�5���C�E�>1�}C�1m�	�D��Y��S��B����r��}�W��i��R>�=�����v��(�ls�z�;���و�s  ��.:���U�q�d�֕4-�� x��3��S�Ch���c�4F���N��'m�G���\G!ϥi;
8/�R�����;�T[�AQ��^�c&쓈� ��/7������j�ц����F��-c���5�e�:(9+�?D�6U�d��ҹ��%�����l9}�8]�)R���������T	R��y�)���{� �]Ҍ��[X�E�=Ę{�R�ljԍ��\�B��`��'+ď�->����S�Abs���F3>~���̈����oB"�{���5B!^s���g	�cj`��-f�X_������&5��용�R����F��
�%�Wk��(S��@%�9���Bm���BV��}G�A|�\x���P}�~H�L<�<�� ��nl0&2ڳ��Ǐ8��A��l��5��'��U�FD��$���=b)R�x
M^�/�2��fb�Y7GF��s�i�&�@9���5�d�����-����A�6�#4�Q�9�|��*�<�ۃZg�4i�ƼC��K�q�ƙ�`6�� �G:٤��#��a!�h�ʃO6Z�����:���QuH�բ�r�O�k殯G�2����N�]=��.V��WGlt73����)ܚ\o��.;����tQ������o�x��qYWj4�����aJ�0�0XZ�$�1S@��eJP�:�;F!��
1(b�@c�6��C_���g�?��+��U��Jz��H{��N	������FD�)�&��]ЧDa���c*�#�bg�����g��{�;�4��#+���cd�w��y��C�m[�36�dat~��~�h�G&!#}�@ұ3 BT3�
�g�L>������w<	i���_��Sr�2�l��O��$'ר�QRWZ�}6U�I��R��U��H��_p��gF��t�S�IJ�&������#II�v8�(��*�
�J
bs�;n�<#5d���;VjK��Q�$xJ� X���
�w���"����G�Y���ܓ�M�<z��g�"�3��	?0P���� ��Z��S]�k��Y�"$J09�������EY�]q48�S�I�#3�/#�5��2� ����s:1"�a��J�	��ɘWP
�X̗��j��U��_��ރ���z����Ky	���꫶��By�3,L��+��W�6rj�X~��/��È�vJ����_�$W6K�;ӛB]�ց2�x��2���;E���՘Q&w�}�-d;���!ȇHo��<����H�����߲�!��K�D� ���C���?�)�G�y&Ht���R������o�c��g80�G�a�Jo�jRs��s-��#��Ы_2���)3k(�-z����P*`*S�k?�D�!���ݡ^�~�h�wb}���*5�`I�����G�o�cq��<@M�V�_z07ع�M철��(շ�N�É���y�퓵o�'2˜+%Ǔ�ଘj�P#�Jt��i�X�n}������G>��+�F���Y˹1s����G��w2�
�bi]�����]�T:���9���hd��$(y�[ԇ��Y!XCW�t._����:�'2��o�s�F�u'K{;�+��Cfǵoo�[�Q�Kb�U>��e\V���8u@}r��V;�_W��b��S񊃅�]�y�����-�K�	b��j��G:L��G.��<�7�L|�A��	%%#'p�H��Y� �����"�^B_�Qo;��{3!*k�k!��;��6�̝���T�{э{�O��@���d��f��{����J1�W���D�%���;�>@�x��Wo�@9e�5��3);0a�*��	�0%��t��[N����^�����1�+D����H�K'	h !��-����	sȯD�5�6��y����H9n6]���{�Qp��Xح�r�C]��f���9���m{?#R:���"�(�SN	J�!�v�.���o�&N���硠�-A,{3g�.N9&����ng�{�a҇ix��_I]*j�T�e��D��|[��Q�Ď�N��t�7�`$3�楳P���sa ��~X1~Z�c�9��� d�n��o���1���!&�\~k�����:�(J\ZFu8�?�3��7kV�0l��'+�
Yz\ǿHʾ��x�D�(�M���B���\�T�=ېoe}o���8`ks�����q�]��T��\���ԉ��'�T�jV���	�E���b�H���=|��%��w~���X��ȹ#�x�e���D�A���A�,;n�(o ���.
�@G13s�=)#��h	D���?��6ۖa�z皼/X��LvFr!0���g��$�H9�����X<��a�^�ֹo��7�&͕������o��
[`���U򤠿��w�����ګ�H.��Z���.C/�g�M-�0>n�)�LHdZ�P1���:�@��\�th����0}��Q����u��EC@$�v�s��J����;�ʨ�F��=D��RN:�n��/���9.b<�όaz�WA��.z'y���uO��*�0d&i������w���vI �S�4��a�c��֪|��P���8�(��D���w��_�F4_w�����nܭd�-+}];�N�
����(�DC��SW��d�d2��
Hj�w�,9���Z�4�<��9<������iyK�S�+�[�*��3N�j{~R��`���w㡵�/$��o��1_����1_���j�`YՎ�Sg��6���F\���,h��u,#��z�o#jĖ���s��e\��ә�Wx���e��O�G�	 �h�O��'��Ӄ�D_Q���3���y0�OdF�c���ݸ{���}T��1o���BE��`E1�G
���F�O�r;T�U��g�񊞌\+g��R�Ӈ�)��^/P���:��P�������Ƥ����wsxi�֚���A�\iT(w�6֟Ƶ�����/Hc!I�Ab
v�Ώ�|�gE�&o���F�y��BȐ44LĂCG�w��v���"�(�[�u�ʃq�PH4�v;f��i��'+�0������8�8�sS1i��cg�.~0e=�L$w���t��p����b짇XŠ���.�G���n9�Z+����~L�XA
F �gс�XA����t�=� 0,W9�rn�����O��X�f��-4��������?r*.�8�{%��ʴ[^�W��'r���4��a�~�2p9n錱���R�����Ծ��l��G׿k1V�@���iR�L5ˬc ~�_�a�|M>j�i�\�~���d�#^�JO@�E������0R��Ld`���|F_.���J"B�X�A�F�kYB������:��(�o��@5����q�Tu'ar����>������V��G���Q��\�p��L�E�`}��Z@ ��oA(9��U"�1L)���>Ǌ�j?�3�͕�l��}�7�@���j�y6f�3F���g��۶��;+�ns�|�a%Y����	
�������A��Dڄ�s���L�j��o�SBҩ���-m�wx/���J�e���̺^o��B^�ܦ�V� z!��o�����T`w�6n��@�aL����� FE���-S��2:ݩ����o�q�Q��ʓ�!�F:�\�����^HnN���\��G\���hx�\��ӎ߁Mͩ|��D�np����N��5��"Z6�5*)�5�����H�F0���~%��"�'������VU�!�N�2����m�U�f���X��q�ˎ�A�����w̦��3��,a]�����U*LY.���GF-[& �t��Z�h�=�PX�N�X���)�ZRk��u����it��|E�`x{0�:��&Bv�W�����ѳ(WZ�"X|�
Z�^����h:��b���rq�ō�U:����P/�ˆ�@(���,�E���'u���uQZs忩e��Uz��-�	�x?Z�9	��CK���2-���{�?��0�����E���񔦨�e�Y��Єt�8v�s��D����-�Ȼ��U~���>pF��W�����<b%M�|9��ڿ��Cۜ["Nx�E�l
rH���IdA��@�A+�J���N��X�(=Fr'!&�)��c�63�Zq˶��;�׌O��&`��&�|*N�w��Nvixq^4��j����uj�z6�\���K-f�q���h��|�T���B�/��d����a���|U�<�����o�����A�?��|E#�v�C����|C/qR�!H����v3~��'>␪H_�����O`9����Nt`i��_Ӫ9թs#h����� ���9y &X "YEf�}�s�~�K�%��,���$�����I��i���0�b�����"դS3�2�܌�۞�Ꚑ��,�
>[�^L@��-���NG������ŃG,l{0\�/g/,�P`ORBI�/P���(��?{���Yށ���x����m�<�1�wMF�KayR[FW��ڊ�S�ώLV�RM�g;���y�l����׾���q�	cT� L�wo��6���f�+�Hns+jv��GO�:�b�b$��^�vH��������8dss��g����l���+�w�9��`m158�8�T��Q����o2�W���"�0�ʉڐ���]�%f�c��Jy��NN������x��� �Fa�$)o<K��
��|���k汘���T��o"P=���n�suq��#A�T͎������~�����O�5�Vl����J)d�^gӣ�7#��ؠ�#<:�uyʐq!�[��a�>����(�<�x�SOgOEc�[���n���G{�D	�z�5>7t+v�u������m�H���x�Hj�v���ԓz���so�`� {��L�ƕ���r���E	����+c�',ҵ]�&=.u;Q)u ����ki�-�JT�7�wW���*����7"O��W��2�	s֡��|E�ǅ7�-��nV�0�GW*@p\̸�*�Z��e�>�@4N؂��X��~K|�a�hFF�Z¿�������t$4ޞ=8=	�L�6 �jw�%޶U Ȑ�Q`��Y�^�;2���[�S��Ɵ�I�Dnn������_CX�<�T<08}�"k ��%���/�a^f�efZ	c�.9��w���~o F���rA,�����۝̴�>�	�p����);��[�� �p�[���`��O��z p��p�"�����;S�ۨ��tɌI@�o<���"��,]����4U����ۈ�vP}6��$�4q>Inꍋ~jS��;�K8�ISD���`Sjm���6NS�s�Ax;+����T�c�>d�]쌔Kc�=.
��2�Hg��f��.*�n����6ۀat���(�#x!�����:���(��w�r�b���� �X\��Ťvi��1��T>���D3-j�(�!�Ŋ�?��
xh�*��E�ʊ	�qU��g��tU�\�$��;�w��\��Q���>�������@��%QT�yOg��>��`$�1��u]��8�;|�����B��-�����J�B&ˣ�u�tHJ_���QTb|I����w�B!��yFxb����V- ��������0��V8��� �ȯ=��.Al�M�5R3<�6I���r=�ɂ
4�d|4ܪn�X�̵B`3PR��z��`2T��^���"[� p*�p�p9��e�8�7�3}�VS���h��g%�*=#` �l�#]�Zd��k��޼֯0��^��4D�ii:)�o�A?��͛Jbt����	��xDES�`"�^Q\�:R��W���j5�?.�(�@V�U�b��
A:\4��9���;]�ܼb��b�CF�vt�Wb�f��3�F�,Z�[��ͤ�uD��*�{�V���T��#GB�Pk����:��jE��b8"���&�DZ�󸀛1R���s^�R�-m��<l�ʍ#Y �ӈ��/	��v�a�)���T*�K�~� �!]:�,��3�ոuۍ�v�S��l�0��`Q?�� �u��U��oZ1|o�%:�ܓϭ���k�����7}�aŚ���55�[�&��mW�i�Q�8���đ�
N�����+#h����Ş`�R������Km��o��ri�G�p�{��o�t�x����%��|Mx�(�XWBr��S�)��&!��>�@[OE�vm�]�;^�Cɲ��*vY�lTp��Sq)u;m/�Q�ɍ��v��ަ~5F��\&��I����L�xut�H���k�T��u�����P]����Ǡ��\���I��>�m�_0M��5J+H�go��/G�`�R�Z?7�.��5�fk�A�]?��%s���XT�M63�@��cB�h�T�6* `�ڪX!n�����tǻO� �H�o�<F^uM*/WR�3~��1Ũ��G#�#���4nl��,M����f	G�o<	��h����Y�X��39��E�#5�w6T�D��@s�Q _Lv��x[7�J�bA+�y���4�cn>�����*��)&L���_��^-UJ��M
~��e�	�Jq�M�w�{Ήi]ݝ�#yh�?[e�^@�?�}6���k-_�a2��@,ʩ���J����A��Ve�G�A��m��mP��-��s9[�1v-^�fX�3���v�U%���FӉ�U����I�k�3�^�Oۃ��	����G��`c�di�tD��������%P�S��OK����iD����O�O��t� �#r&������K��{��9���$]��;��$3�1��"�Mq;�8���9P���.������K�!��L)��Q�s���Y��~�������O��� LKis���qݧ��.״51��#��]�։ZI9t?&�����*�b�A�Cd_n=�AӴ�Tb��tG;�C3w&���CKba&ͬi{��찮����3�/��:�X��\����f��f�Y'\��G�l�	%�6�e>�P�+A80�ӌ98ݮ�iB�y�-ZE���ԑ� ���\�%�h�>�*/,��W��K;��Yt*m%�p@�o�P�������j����j���)@����[�S����*)@?���B<^���ueD6��ޕ}m��{���`��<�	����v��ɶ��[g����)=���JKg�xK�aդ�Q�'�]�!�4�f˻?\=mGY/�_)�Z�=�D?ɪ���n��X�L��������-dV�<���0�q�۹)U��i���Ur��s��Q�;���/<�bil_B����,L*�)�R�
W6\��zVZK����4*e��%]��3�wt����;x�ws�$P?{l;{��3UF�ňj�UO�?�w^�҉$��>���Ӯ�Ō�vN�4C'm��c��w�t��܂�U�I�b7;#�����(�`����eԌ�[ƃ�~��Q���ո����z�`�������t��ڨ��}��L���y����#5����bv���nE[�c�M��Ay�B��	�3��Gu��V�O$*���H�}w���?d/����D1s	��M���#�u���������M;T1�xXN1;���jչr����w�G�F��<�+�8� ����`U8{�})A�K30��4�Ќr��@���Z���V���6���������u޵����?�Hep��%�q��y�� q$j!�L44��Т���m�<!*���\���B�phU�艽]��gғ�uݿ�S�a��?�����=J�R	d��N@]���n,��eyfI���
����Z_�^����c,{%�UE$�i�t�� 3��4v�o؈ziN.�${*uue;����o�U�RJԍ�����lY�ӿH�]Ւ��F[��������k�HY2֕-ni�iQ�����T��}�d5�8c�����;�r&�ޙ6�#J�{	u���1��ZJJc�\G�^r��Ḻ�
]H��ul�P%IE|��g��Ŝ�!�m�!�������N]Z�j~قr��$h��{�d-�֞�O|��,[LŮ0F׶�_��Yj�6�Y��o+��9�NH�h�C�����yɸ7/3|;W���}�o�w#�bA�WE�N�b��\� ��E���o��KT�
�ES#�W�Օҷ��*֮�z�|��gO�	���ԓX�%҉h��I�%�JQ��_�@��	G��_���I�iY��^��XYU��^��(]0�ְ��K�j�`������"[_�M�~���a	�f�2�c/�F:��.h>nI@�'K:R� &ʙ�Cc�1UUd�j�Hz���'FIC�.y���xB?9�Vd�%���nLj�ȳI�
�]�Jzv�`᫨{�3ˮ��^�c5�_f��(����:��g�)Y��Z���b����=�w�������7��
vZͧ���+���E�ίf�Ŀ~����9>��sT�E(���\|wx�=`p0C�1Ox��G6�y�_}2�7��e�u���[��i�9S;��^������*U6���cm�B�A	:������҂��0z��o���Y�d��7hA�_@�3�����]�	%����h���j�6�˴Y�>���`�?ߟ%�!����(�PF̇<
�^�Rq���Cٲ��\�z���?�M�w���e������_P�`A�.�����u�)q}a�AH���r��~�rӜ��[c'y�5'�>��b^D:�F���t��Tu�/>���������>��qtD���o�u�QTɥ�i��`>mM�|��3����K��X5�c⥅v��[������a8A��Y�<��>3p>�v�����5םŞ�PHp�*���Z-�1�\YA#����$Ҝok^b��_���aM#�f� Wn�Ӣ�2Lb���"r'x���zp�G�n�ó��;onB��j�f�v�"~�g�o��|<�<\+�'�cnp�
?܏
r}��i����#�*�>#t��Vej�>S2�w��
��ޠ6?Dv2:6�8�� S���1u�4G�B�;D��K�3_x43nD+���ۓ���u*��b=��N4�X؎�8��JQ!��*�.��[M(�g�~m8y�$����`�e����!���y��(�X��tCO��)�����1�\}�h�n��V�ӓt�j��;;�Pu�@����{�l\�H��U
����ny�]6��i5��^Wd��7i�Q��1q-纅)u������]�j�e#n�c
�����-wףoȼ$Q%�a^�5v��}�,�e��!��-3�Ժ����e�Qc��r�򤓞�s63�����ݦL��O�}�����6��c����5�:J
��U�g��2�F]�j;r������1*:����G?J��c�JF)�l�F����QNg"�ә)ޮM7�!b��Et}��#�lЧ WV�rUN`#��WS)c�-���f��8�c7gSE���*��	lƿ����Z�N%���;�����m��'3����f!۞�n+qy�&w>�|�<���4Y�����O&���(y�Ra~�������bu���Et͆�){�E�S�L�S�)�4����aUV�9��u��G���
]S?!
Ƴ�lݐƹ7�İ�l� Q��|�{����߈���������/DB�;�b��>V�]g@=��?��o�N�������7w��eܸ�a&(|�l۲j�Y= "�aV%�����|-�4i�F�d��+p4O	S����o�? �x�0��,�#�^�X�E	g��h���:W�{H%P	V~Hz!J�ʑ��pF�J� C��ܭF@���c.q�¦u��
�oN)G�o�c9�����.���w���rP4=4�<��g���9�����H�;-h\�p�&����m@���ͺL m���[�|+�.�z$0�����qI%�?����F
S�ޅ)�:�kw�ױP(�p��C��6nQ��|�5�D4SVF]R��{6"���p�ЀN�V�Fhݛ����ųH�VEW\�%��6+���N��-H���Z��8��6�"C0p���	*�$Xl0A��qr)�w�E��� [Ɛ��~D����4n�{Ȧ=�b��(���T���h]?風�B�4�1�ôJ��y�}���?�_+ٴD��D��9��z�#��&"�WHacC��P�[Q�l��*����'��(>�r7SF-S��	c= t/��\:%�9=�8�9r�!!6���-I�4�
��Z�-�Qz��B�V K��BC]�	�ۇ�1��¯vD�J"{d��g1~�kV���EE?T���}n��P,֯����8���T>��n7���YQ=U}~We�M�%n�����h�/i�nzAU?V/�+��[��FB��<w)GJv��:�`�����Jt�߷��)Jd׉��������)nqf��&�T����V�BH�g
�o �$H���)A�T>,G�a'���O�L9 �5��ET�K_�5u�	/�w(5;��IWy�R�{��b��[��yr���˵���9�;8<>dSrV���M�X�u�;f���;��B;�iT��3M[^u�ȵmoR���6�%t��ՃQ�C��D�8x��!�L��o���,���,& @#��T�|��P�"~�EZ�5�P�y�0��瘕"|��s'%��g�ZYp�E�/C|S�t�u�&O�����0\ƃFRǢ�����
���s�����\K��#��.~�r.�~��V��k/��m�u��H�4�|�)�!#%G����(��=��h�3~�T�@͹~)�9~�X��*E}e�[l���d�6w�iKGr_�nLs�v���c�<=�@:�������kz������L�Z�9>�1rJ2�F�h���� ε!���,W�M�o:Q'd����]@���؎�U#�n��z�a���T	K��kjI�޷�w�s3�	&��a�`	@Vˤ"k�
A��l���Ƈ�h:�ڈ�mjWRr^c�ZPn
�0.�qi�MJNo�Y���*�7��-?`��}z$��j��7{>�=1l����9�ct��V*+rNc�֗��R<�B\h�2�r4,��]��334�$����Q�
~>���i��	;�X��CؠW�-Qx]%J`��)CL��P�6?���.��S��$z��f ����f�����k�:KY_y�$<>�*�t]��6C�,1v���ѹ���ERNL����0%��>f5Mܫ_�(c�Լ�[� �M�/֖PX��+�E'�q��)hV�������k�=D8QƵ�o�������SnXS�m����q�<����(�2y�JV�j���j$�8���J	��qM���$v8	>�?q�Ȫ)��$W�Q�\�_b�A��Ϊxo��� ܹ:@}��я�l�n�GG��H2!{�'ޢ�\��;-��5�e0*)cy�N)1�mcX�����;�n�F�}_��:�����t��I->9c�������&��ѹ]5�i�vmA6-��c���h�X�a}}D�Y�u�&�d����-KL�f�|��o�r�����p	���`�Rs9Y�i!�����F�K�4��ۅ�{S@��D$�!t���!�Ȥ䱕��s��1ϛQV5
RN�[��{�7�;s�
�X���XM���(�CD����4�� Č�=��&z��@�9m�Z����y�*)�ʞh�#R`x�G����ˁj�;�6�� �(�%�W�,��粓۬s�w��V��>���⌍��L9���I���t�Y֪Ɉ���2`h����+[���s�U�,f��?��$-
���:�RÍ.�É��=	Ѭ�~�p�q���3��ӧ	,�$��1���J�^ϡx,��{4���l��)����d����|\��G�4X<���秖��cθ�D������ܺ#�=�>�@twX�Y����x�7j���x����۟>Bf̱�C�5�)�Q�Rf�5�^֐�'߷2�6��1&� us�:H=������c_�[�y��˭=���������m�E���
�#a/��-G��<�H{����}����?T{�|�3{0�b9DRzT�9�ts��� 6 ��& ~o�\��Y��\�q���c�.�>�*���̄����ʘ���.�������_o������/叡�`�b{l�����P,b����j�B�(,U�[���><�xڳ�/0�4K���m�����Pg�L2��ZJ�b�������؝���*2 �f����D��˝y_�k>F��[SOކcI~��5���N���+ec��sF��~�t����Q>^E�+C�4e���م����_X��U�k-����=�����.���&d�����b���S8+���^z(�K��ү��29���ׄA��ތX�a�KT���,Q߁��}�5=�}_7L��0?�\d��������˷J�5�Twu�㣮1W=Ĩ� �s��@����{ ��&4���u�{��<��i���2�<�+��%�d��Q�w|Ά�@>�d�p��{��I����E?s�^^>{rz�Y>)
��M\��Ǖw�Yǡ�2-ڣ�iI�:��M��e��f���bW��r,1�Ц�pd|rz���D����Li�s1��!t��Te�F�!���$Å���/�`��ۛ��f�Kr�ű�gN�R+��p��Ȩ^@��� ���u�
A��C�12��=lz��N��$J���p|Y�qZ�������wAkǜ�"���XOST�[�G���k����(�t�C��^�k�Ώ�r�8��_��~�E��ԣ��-l}��c�:���� O��Gm����{���#d���^c�o���K܋����P�#dk}W<L��Lb�Tn�4�C	2
�`�wGoq�ԏ�ee:B}��T5�9 [{����<�f�2k~B@��E��G��`����V�"��<"X��%��~3��s���\;���rb4����4Λks|T�Dq�,+?�:���9<�	q-;D&��m��ή#�uwXn�	�t�y�Q�����G_�G��2
<����2�1����$}8(�R�W�+C���9��CZ�Z��r�\���ѳ��$�$��c��i-|�F\5�������S�d���V��\>P�*����/e��b_�#����$���d �:r�kZ���W��i�Q�l,��������%�x��1��vA�?8"Yrbt���r��\�~B�kF��t��g@��L��"��Ά��lVV��nt>M��<�<I�?iqb]D<�Ia�U��Ɩ'@��J�[>*Go�1�ceTp��r/]�����OA�*wC�W��<��>��b>�� U`E��8D��~s����G�~ܞbu��|mKm�~��ZJ��Ixž���O�v�8���mЇܯ�/o����㳄��ZZ��j������j�V����wx�ӃrM�����Zo��?k��g>�#c��L��Բ`	p�?L=��`�Β$�A�
7'#�M����<�����Q��@ٮ"ԦF�%��ʖG�0��vl��95��cu!���f�\��iKS�)�~����+y3�y�ݚ����������P�[q�x�w�[�Px�Z03���x�$+ț��h�C�]�ŝVQ�_sUY>#�)/y�S0_P:�5�#��~~;�d�X��K�8?��^�hXDB'+�Z��Mpwk���X���fOR�p�Cف��ϕςJ|]g���	�����m��e��䎿�2&���՝YH�iY�� �%G�q|�|���T��/s�	�Eh����"��\�I��O��|pZ�=��e���H�r|v�s ϓD���ա�c���Ȭ��k!Se��1y7����m�c����w��H�Gś�C4+�nY�d��ʥH*�%O�Q1&���$����I�8�����!�H:J�1�1�S(�=�z��b��XB�0�aEK`ȿSU{�sc)Mb�~&�&H���3& ��d�zv����(��luJ�!S��;���#Zz��!U��t�����a��(��(Ǆc}uC�y�����oɫ�<�60��%o,�����~)��~��k�&Hd�c��HLg}Qcj��p�Ｄ��1߶5jar��Oh��pz�/��8�G�/�hsєG�?��^%�f���b����^�ꄞ�<�TUb��!��0!U��'�yX�[�fPq�1��G�c���{��q�Jw�2L��r��1���*F���Y�B�GԹ뮑wo�^NP�[ǂ��J1AR���SX���%s �G���{V�E��\��C��������B��}�监qhyyy.�ft,���R�)�ͩ�(��ջ��u������}qH*D�.����h���\�,v�A �%�x�[89V�x�b�*)�1�����s>�+>���0��Ad��0��7�~�x�H�P:����tge}�ğ�9�p�{��dWy��Y��(�:�>��2�qP[�� >?��\)�v!�m�-�J �\��g�^̐q�$AP1�%�D�����C<B�s�K�o�oc�"Ú��ѳ���W2��rXc��MN���C�����~y<����^OqM�)�Hʲ��~3��%(�T�K�4U3Xe�|��q���&�J�3��S��[	�	������X�?Gmh�oو�(sXg8�p��Sƺ��)W��|�'0�G��)^������� &ZZx S����P׈����F�6�*���zĊ���r�BWm�	�^_��o]S�]"�=M��@>�OE�2�Vi�F ��!Py�d�+�%1d{I�I��/@ì��Zsz�!���X��Ӛ��e@-Q�k�X�z*%�1v[|&4/��@m(of|(=��� �#�a��L/��H���mM҃�#yR�ID�-AL>��WW{diKwI7T@�	��,��7r �|9z�la�V������2����Xb?_��Ӡ~�VG&��&c�������P}�e��D��廃jM���'2�S��-|�~���qi3X&�Щ�㼪FG�r_窫�v�5y�n�����.ץۈy3��'fx�:��"3
QB�><g��k���Y?����^i��`�t�d,�
�}��}�6j��~5���(��h~�oh��w}��=Aҹ����wM�҈ݤ��d�ܕ��ͦ����d)mi[,�^PwP��7��t��]��k�xj>~6��)�,���R���>�/�9���H!�ʺ�*>&y�+��5>����R𬾫����ug2k*��"�Vl�Zu�!����ՉG7��L�qJ�tP�\�-������ӊ�ԁ6��)�w���'͘���c�_86��E���6��,2���j.�5q��8�/����y͉LS��"	t�l�߬j�߉X�]�<fEu�&<dM�r�B��;���:�bR�T�{kCWe�]{$_a^F��L���h�AR��V�a���%G��OsMq9� 8������fݷ�����֚D�F��`Z�A���5���|dL{�܈�_�T��|�ANr� v�G���za�y��sE�c�@�5�}�H�0|�i9���|Pwi�5t#�ߒ9 ���wi:���6��iBI����S�-OȔ�V���c0�io�c:�?qm+E�bơۧL�dO1Iv���^�����]A�8,����G�ÿ��n
);y��:sQ�%��KQ7䌑It)�c� Q6Ǎ-k�V[�����@X�Qߵܨxbkߚr��ɪ�m�-f��� /�F�y~�*a����l=��T���DN�3�E������c@�,=�
Y��<��>��j]d�)��-��"�曆�E�H�(�4��	� �/��d��*f��u��m�k:-�P<(Z�^�*M �x����XTT��5{����S\�I�@I2Le�IT$���Wo��1���s���v�L,�*���� Bn��'_��о�Kq�}eW0�INx�/���/�@���A9{��ȩ^�=}�2kD���a��f�]��Q�J�<7��)k��1+!��_\�nFm���n�@BYO1 �sEh���H(�ԣI�����DDӸ&�2H�Ư&�?JGGE���k� C�	��]c�\7��%s����<`�v'�.c�7� ZI�$���W#.)��E���cGB�M�D���aZS	�
������^=d�ѿ�<�R�V��H	U
�x�EҦ| ������VgZ�J�yߥ���-&_��0Ǜ���YX'7)c;���"TS�&��������]�n��!��I��`w9f�T��fG��:���ԗ��70��'c�!���m�*�r5� �K�������K�
d���\�H#�z4�Mg�06Y���ޏ,�ТZ�Hs�>���O�n��uIn�~G����oi�u�ܘ��dRRX��c��OR���nԀ����:ny��7�������n!R���\��R�*�;��_�9?O*�B�a��ϓcu�������(0R�^�hF+x@*�T�~�3�ѬL�y��>wëQl!U�nKIJ`�+Y���w�Πp���M ��1N�' �MS����� W��颎I��Ee�W�8�;BBl�C�� ��i�ͦ}£�.�+���+C�#Z�/���̀�F�Ӈm���Qh�Y d�9.ʱmDYLl-|�
@��L���t�ky������Qq_n���'�R�������l~��Bs�[4��7�5\j��$l���T�P�7urܤg�h^en�}�%tk+�g>~�nԲ��e��F!�0��}�]�X�i7�W�@+c��m�0��9��K��ŬVN���w�>��!i�E@�@3�B��O�Us�@�Y�� �[��d��ù���E�5��9����a����ۙ���S�I=p��H2����jN}�Y���5��Pi�����TA�5b��s��<����뚃�*����p��,p:���}�e ��D6hv�-щS��6�� �����d;����yk���(�����~9�TmJ�!gq��)$��;�^[���a@\��?f�tJ��ə��,�'T���v�W����-߭+��\J��0�ݤ�d ��J`E5�/fz~���7\���ǩO����h���fO�'"���@�x\�e�bqD�E�͂4�\n���'+�KW��U�S���4ަb��
�h�_4����α�`�N�e�Z#S�,���㯤���z-�eH֫C攀�/52����O��ƀ2��IR\��
'�zJC����SǟM�4��$�}�.���|��\=���hu��f�&z�U�����{D �{s���:�c=8(���;<5�R��zL�M�-�w�j���6��' $#X��}D����#9�X��kd�����F�O�/������Xj|�lH��D/
�_��ۂ�x�L��Ǿ���h�.&
���@ �,��%m
dE�6A!:��n,\���#]�g�]�x��b���ý0˴d%@��n<�@ O
� ߇ݕ:�&�J��N{X��ޖn�|�5ZEd$� �8�8�A��kx�(L<�X����3� �4/�!U(b�;:k�O5M���&�-g��Ň���'�+�N������+��Be�W������wݖ�WՑ�D<��bGj�XU�7�7ǅ&��~77
��8x�e8�� �z ���5�K�i�������� 9���ֈC�D�j���M�*%��Cl���n3�=�����@�1���MJx�~�7�Dr��%�j�����4Rx��÷0��;�B� C����W�6.�������ʩy��w���f��[i��Gc�P�{V7��g�)�t��Ƀ��Α�6��s���4ԁ�e#��5d��/����W�w �e�T@�����4��}D�
���	�'s�#`2J��I̷|.rz�5��m�˝���&���t� ��
f{X���[G�|\7��_��!*��纡��bȥh���qU~�.�1��|	�1�b����'~�մ�?&ٮ����}z�!��>�A��	#;kt �3�F�S�h�����dg $��T�f����?��W��܅�x�']��F�x��Kx���9ʪ�[&�һ�Rl5ON�����yX'?i0M�/::̝ӫ��C6�TvŐ�V$��pك��v��E�5�AbT` q����<��D5u�B�j[���D�)1�L8J% O��ڹ/�: \r�ƒ`o���������պ>��E����k�~.�"x�����m�@8*�rN�!�<�9@���jMڻ�B������i|k�ꃪ�l?J���G"�����h�rR���5���lziL�6>d�4枆#��~F���|FW��:^���ĳ�k=�3H�3>h��e�Mm�6�V�õ�����K��'���S��\�MFV�GX�׹��]��X�c�,8^f!��z��]����9Swv�t�?�Ǜ5��n�Bqޝ��.��^�ς`�Z��%�¥"ՄZ0~UQ.����Ϻ�<���
����e��<�Q@N`�8�tg�TX�Z)��.��ɢ�zc��2=���[�d�AU��r���IkyY�u�UY�P���`�~���/@m�p��(��Hg|�D}pG��Ɓ��j=��9N�{<:��3a��σ�Z��1��r�^Ԗb�]
Գ��ϙ��W�Lu`�EPS�v��J�ںpdGu�϶g�[!{O�W�.̿�
T�:�7����q���tE�.@)�?ئQ8�Р�TGA���F��\PM,A�h�4|�e�@���Q��w>�L��;MJ�Â��آ�i��S�1���`� E �;-B����k.)��:-$�`��JMUV�k�t�]o�{F�[��]��*�4�,��zOE���Ƞm,� (K�,�x㷇�\f�/g�p�կ�^����Ԧ�Q�18�U�l�+�v@2�H@���s64�EM2� ��|�%t�0� ȸSH�`uJS(C�?
��T�μ:�d[|�\2'.���s��ni���蓗�����VD�[H�J�mI@���Z�����S��9��b|��]&��U̽m�8~É�����=+�)��n� 2����\˖�H<��XԹ��C,��x�vІ���T�.�M���G2 ]�\�1�=77�ǁ�Zq�X}Em�G!��E<a���3����
ڻQ�kp���Aqi�'��2�˲��̫��G�5��ko�f�2��������)_ѳ�ׇ��H\��y��Σ� �%���{�*r�U�����	�H��\@�z]G�Rہ;-��x���DfHO��#X]�W�g�Dd?�k�n|a6���>�B`�Ɉ�$ea���d*M��?8 I��l�K�%,���Y���vD����JD���t~+l��CL^�!~eƏZ�����s����$Z,�TbÎĬ����C����sh������w����p1���:>%�xy����G�|��"�r����� tACo�U�r���b���J0}dY��$�shE�5���	
���m��F�w6]�v�B�IV�6l/��V�B��ң^	j�
(J�Y�v�.i����g^�$�*�Ǡ���epl�5��f�ۧ�3H����j+.��k#�: U����n����H��d�FA�8o&���}9�3���<ۜ�,]��6rߕ��m���5�i1�Dh�^X���$��R&�� ��� 	]U��t��ᕎ���]�����3Nb��e��b�K?=r�t�W(�O}C"c�L������ɐ�ˇ@tk�Q�#IK���S:��45?�G�x��`u��p���1�+����
���*�������\��0^�oM/W\E���!TՌ���,�h�-��7�PepsnDF�a4��*��6��TUCW��t��:D�O^���P��I�I�Uv8-!V�'�PvNI,����f	�sߞj���[^s�zӫ����lu�����H4���3��ft|)m[����v�i��L���Ͼ�C�Ʌ��J2H^� ���Z�y�1�]w�>_��bd>�R��@	���S�#���P���i�X�=�Z�oaLD���������J�G�n�5�uGd
�Y6˷ڊQ;ͧ���li�_�"�d��UHm&$@�L*ηy��K�*{R�����t��R�B�R�8�ZP�A
o_w���T�	�g��u�/EB�:e0�lX��c�W�L}U��?<��\O_�ʧ����m/l)�Ƀ��hX���7┾���X�u��Ö��}���T�Sa�ޜ�3a�\zk]�$��LwYxg�0owL������|��tٮ1 }Z�݀�A��;dA�+�EP�?38��S�I��6���05���{s�)�&�/�C:4��¨qF+��\�fC�;�b�8�ԻR���c�.�m6��4T� ���r��φsž1J+&*��߯��xcz���t��#��XE�Om�q��հtN�H�^�^
��6
��������mK�΃���L.�hB��$t�7�� �L��zT6h��TY,A��3/\oe�۞�	*�k�U��
bl��j�"�f�wg@u�
����fHI���#Zy�xG���{}���U�� ��Q��y�PǝXl9ֲμA&�O�ߗ?s�j3E~���䱰r{���0!���&���z���ԺZ�Rr'��p���H:o�T7z�������~o���&>?���8J���W=�"3��'�"o��ac���p�������Jq�l�J	k�Z���g��N��"�"�U����JqW3�ӹ�,[�EO7�����x�������"�� NG���W��\�q�^�����Z�dcH�Ι���E�eז�.��\������q<���s&����qZL�,�8��,r�n���I$&l�+��� =�D�7�\_�%�(<C��t�ZDA�]���̺2>���+�vuT�>�	�-�=�AQ��W_�Mn����A�.�̘�s5rLE����r�SЊ���ؽ�
�&9�������Fb(�Q^ʥ-�C���!�g�ͫ$�hW�z��Vπ��q�a����!�5�J�hgw�������l�D
�\�rB������F�Ϯ覶O����`e{d堾}�]�hv�3�/��D ̞b�����z�/�qG&�(���$�+q�{��}U�ݲ�w���N�S��"�;ב(H�I�a��"XJ�	(u�����] �#��!-?f�m��PI���צ���&H��&�-�9��J���H,��>��aj��������r&�h�%�gWuune��:	7PG�����vo���ૌ��#G�;�X��q�;���w-oF����s��V"�	>m�����bf�%���FA��(j�F����r�tA��`�D�kL^�n�cY3;��@G�#|]�o{��} ������"�Ҁؒo�X��7�v]ꨧg�R 4@��F:��8�zD\@�^1n�F��k��0�t> ��si!P`t���G3z8%"[�%�,2����W7~�`2?�|@dlq�`��Q����V�Ntj8�^c����_Z'�_��Ė6�h>��:�*2,3@ቼ��Z�B�,��O�����4@��g�I�ɑ�����[��ҿ�ѓ-�C�v�x��n��M�gj�� �ᕕ��ӷj5Cm��̪x�c�M���M�M$8aD	ۃv�|A�z�%�!(��*��/h`�d��3�-����v��̪�V�, ~��KcMT���P��?��%��<���Q<���fv��.v�;�O<���cڥ���C����ރ��x@�d�y��.�8t��-�,{��$����6���F	 ��|�ܓ}����b��ю(ց�+�M���S�H�Ĉ�R�����~]���@P�ƀ����?F$��7���A���
�V: �o����������%Q��$�����r�'�F��0w�/t��=��p�o�WI_��.��q�$�3��g��~����c�����)�EĆ�P����4^Յl(��v�������c�X	�
UNv��J��n�^�6R�y�dA ���U4�{�����56�&q�}х����i��ɸn�����X�Dn2 �*WT�נ�u�=
��|�0�c��E�D�L2e?��͓gdDz3ؔ^�񍻌_%���X����������W2���u�q����W�3�Li�F����L�Խ�fB�:�{B�	�"B�N	f��=��g7^�0�m8\�Be�v�߬tS��l-�eQ�/���A�`�����x�<��y �S2�����	��Ò�@D^�
�_��}�gI�mx��J����,x�Fm��
���Q����b>NU*{T��H������I�M�G@�u�;E&\KZt��Dţ0Ԉ$[}oSb_�)z�O4�v.��Q��*I4�#��6Q;�r���,}�]��q��qQS��%�݉���fD�C�����+�%U��yߺ�6k���y�E!_�*��P���;�9S	c�=6@_9S�	`6���w��!�wɆ�hFX8 ����}��׉�H�5R��^Q؎N=�1�r�DU��H�2���}���S_��| =����*�����R��(0�3Qh�coD��$��G�q�6�s��:A��ZH�cY6]��Ͷ�е�[��������"*W��^�x��> j\g��7���.z��v*�Ӎ���$���=SS���2%-D4Yb���7��76l�_���ڸH/Q

:���K,2i{�iTz<��s$��U����Qݲ�7��
-P�̤Ѽ�����'EFuK�����	1�
�'����գXa$�W� ���S��w�|�6��+s��Q:�J`#��~da���Pn��-w�^��F���������r�v,��R;���qJ//�:V���6��w\���j�����B��� ,WPpR8x<a�뼧�
����1���qm<Bf⋧5���l��5��Ew �z�G����il׼��*F���h�n��⣗��,%�`O��sv����?	����?H�:�Ћ)��am�5i�\"�0ZA&���J�ls��Y�[SYɏD�»�-�(���v���B4�^�L��Ɋ5~���O�ʟ���B�짳��+�V����� �4��_���j
uV���<�x�c]��z\a'Nrn
7��R	5������u�/D;ي���	�d��h�F�Zh�q;r�Oik{���X�g��>��C�f3�S���M�p�w��n05�P5�~u�k{,&�3�V�a(��nm '¢�-]�ǂْ[�:K�N�Wf9��X�[���-.s��~b��`�|(�]	'T�27�}hQ�~BlH�&Z�̆�o���SF趧� |����Ғz�s^i�T��0�4�-$�C��ʨ��O�-z�Ԩ�yIʟ!x��m�ߜ?u���um�'�H'�n (�V�"ֽ�`��. [}��vC	��k��^D!ג�D��C�$���e��6�߼<��	�?{��GFK�]T����y䗋~}��횦Q�B͖�s�!�e�*�E��l�#��m:�=���[��u��,��(:��֬���@͔9oh�+�P1�D�qv�|%�J!�G� �g|�!2�.4�Zxx\���|�~�$�ٲB��)2�[S��\s�" �!d�3鞾;x�	)l���X��YV��+�[������VI�?�$?f�����*��G�GY�N�{b�-�2M*ar��4��`���wB��w�qy̠8�I
7aw��,x��Ѯ?+��ݎ��"_v ;��>x:�w���?i>�dY.��C��,�(�1-妍����y]���H���
6�:�J�b�TA����S}i�UN��x�_�zF��h�y-��o2�7��� V��:����7lǏ
�2a���']Ե�:�o��"��3����+..�k3c��_@�t[��2�&�������Uǩ@7[���A��ղ zQZZet0T3��R��@��QQ�9�\sC�T�N��p���(#�\E�����KGp���q�j+��z�9?�[�_������6��{3�|��N�A����^�����b��\�Gf�M���Q^~�XJ��y��Nm&$�hm��\1��_����tUd�oG>O;�R�S�@����M�T�����.�Y��	%T7XR��~>�_�[˵�A"��AA�h��Y:���	�@���m�5fc��XF%v�NI�Q��f�Z�3oF2��ע5S�$n ��Jz3��1%�Ѿ���_\��]��t�Z7��?�����<	B���L�apFU���M+E��J�	?�1���,�����ɈI�v��g��NVt5B��v�,a8GԄ��5tCD�b<w�܉{�����h<���e���X�-���ur�)��ƚ�&���"'E`�����mk�rV�1b����-��fo�I�4B)E����J(�j�s-�2�_.�l"��I��w�&�[>u���7l��z�̭� ��k�O c��W9��GW	MkW!V�Y�(���������~<��$%��w߅%e�=8	S��PIRI�5#2f�1{ʂ�n�upu�U����à��ݽ.׾�BXX�9UL���D�����N���tZfj;�&�+��2J�_���fLl�� m�o=�eS�����CN5f(�҂�qo@�i>��uh�p���T��{��#漶��\2c#W�?��;i"l��>�!���A��":'�Y�Q���<}K����,=�H���w�f���g�]h��>*�Ť�q&t�CTJ��7�C�]`q{��|2��۱.��iuI�D�Nk#_�-���n>�~��S�-�0j�ג�4���<����`�(�JW��
f���ڴ�z�
a#5<� ��7 ��an�]����Y� �>w�r���?πe�ڃ8ۢj7w�_���	9�&LZ��pI�}���UR@
�C�uU��IJWG�Ɔ�V��4j����0���m-���wW��WP��a�Ҽ��vۓp�ZAw�A��}~#x��7������F��;�>�N���M��o����L�j����< �0ery�2}>aF�:R��+wG�t؁�w�O�:K:ړrI����ki2c	��_�o5균�?(�vM�tA���ge�3��7�`� YzW6�\����q�*6���̥�55�1��Q�����}�b!����z���Ы�OI�Sly@�Y��O%,q�i�#��I�I>cP�b/��1�'AFE���J�*c�M	��Zo�?�n�f�`����^�eB,�6�f_�1�n�UL���M��V�̤��U��_-�Z����3�;6XS�V9�Z"(���_�7�ޤ��͵rY�hz�
9D�땤�'��k�6�&[�I�(G�6]+yQ��Q��{���)�)19C���������^�tZ�Y�*Q��v`|d&��&u5�lj�Ց!:>z²����"B��QVl1w��YS�����j�$�W�9'��.ؒ��Jr����~	)�;�,�s*w,���hg��6�����Z�k����(��ܮ�{�jk�қ�b*���q���c4�Aվė^h��V��!��Ha����:0�1j��xA8H[��(2��;�>�����'g��[����gD��7�����VU�@]4��D	������"����@��"���ȇG�vn��V?醺��T_�����k^x؟ؒQ���V���D�F)W�����5
��}�wf8�La[8����FJ�
�_Se�
��;��}��J�Z7ɉ���`���0��6d2��wK�b��M�=ɐ@ӎo�����ꡋi�7r+è�"���R���9���V��<J��n�b,��QyR�Cf�����nk���� ����|�%K6]�{֤{IL���הX2{N�d+�Y����Y�o|��s��1��?�0��@'�#���F1��h�܆���俘B�I����;�x_����r�#U�ſ�n	S�0�#]>ڋڻ�&A��V͒-O|��l&���Ƿq{,���/ ]�,(�U�H����~։ �.v���[����n��%<̴�q���O�\���G��P4�X7_!�+.{��wI�
zo (b��aZP���d[&���)�������w�אdf���1�|�"��a۹&��q�*��<*1T���k ������"�yt�AIg;GX�6h���I�¯t�����<GT�����S����7���0��Z��;�ͫ��?���(��`��xIi`v�:����ևt�jL��JՃ��LD�9_F��D/.�gfJ7c�.l�"��?QW�������A�=D���|�?V> �I ��^7{���|b'j����ܝD��Pw1���A��V�U5�PyZO1�v�)'�R51�H�:��ch�5����Qb�� �E�\(���C�Y��d�:q�Q?w��)NX5�OY�F� Nj��P���W4@����܆���H�s�&�d��B
�aC-��F!e�{*����n��Hi=��ϱ }��d�"d�ѫ�cm��5RF�#�"�&-M��[Y�]��G/G�C��G&<x@���xx��yGtݓ���L
���X��},��r*f�=�#] ՕYv=
_;��_ɗi+p�_�v����Ou}Ɵ5`匯�H��)�"h��g��=OBj[;Fm�ՊY���Y?�G�Va�{�)І�vr�R7�F�v&f�'r}������u�'0�)"6����JR 	J�k2�sv#r��DȧY� ��p1�#~��o��.�/9A;������C=`>(��B}�JV��a�]��L����h�)��+Ŏ�,p#�����ПP�A1��i��A����-zu�#e�Uz}�i.|1�7!J�o`�n�YK������#��͵=�7��ۍ/zU��"��{cn#p�HG�N ���=p���
/#}�@n��]��g�R]Bw��>X\})���$����W���B�lh�����3���K���IĐY��S~H`'ӆ����	dg�*��o-�ȑ��1S��7�����ry�?�@�S.�����e�Ϛ��y\�y�h��-շخ�������{��<2k�e��+��g�,���.�Xi�L�i��ʛv�`?��X���y�O�t���-S$�j����E�ǝAp������!�#O� �I�A����U�44blo��Xh���w|���<9�`c��f�Hs$��Fۺ��%�BD��c�
�/u:��2��Y��E"�OGV�
�Q7��K�.7kg��+�M;tk-��	�ݮ\���.왌�������r �ǧQ{�9�:���N���t��ԃx٦�qX�<v��xQ�	�i=�u+{��4�8��n)�EO�֛v���b�ĸ{ҋ_$�C���GB\ }�?�}�)$���6�^=BEV�ie<8������-���J�lXzpj�0;.pHm��:C��t�l�A�a���b�n[���8)��.��%����~ ���՞'#ec��=?��>�XC���_�j��r��+3��ll�nq��iJ@NcqCt(���9��`\�J3�1	W��B����� S�tU�^jI�IL]�`�fص|
�k�"��d����f�M�u��\�q�;���L<�ߴ�s��C�p経؇!+��m:��)Mk4Wd�a#��?T����ģ��f�Ӆa��Z���G�9��x(�'�L��|э�´J�|��+MTT��<�����~b��5�d���j��=6�1DW���@��Fw��ӽ��!2����NO�?=[+�ydL�̐	����I���ad��X�z��h?�Y7Zo���T����_����[~��~�Gr�M��M����l���_c��:/�9�G�`� v�e�<p�ϥO����bZhA4<*���WՍrj>���L�hL����R�g'4�fQk��Q�6eÔ�@D�b[���Z��NyO*K��l�|�d���m�ĳ�4�H�T΋B�x�ͅH�Ӝ�/���p�k�b�@]��D����ֺ���ʙ�0H��Ć�,�yA���E��.�*��6!�~���ın�[x����ǫ�;ti�����ٲ~�Oɻ柗a�.+K�i�t9���)���$�i��o&��P�psN�`t��]�CD@!����^�W�ob�N���]��HGvb����ux�'yrF��[M�S�**�ꥉ7��} �
,B(P�_v����pj_��1����VD�L;|t� ���;ƘB�u�z5�f��B�桪`������U��5��":���'U(�~+z���r�)r��-��a�?7��@�"�ÍqԴ$x��U�ѐ@9L7�:�������z�T��	4|B&:�t3�3jB�&rUh��� �A-�����Ic��i+3O}Z�r��R����y"�@LD� qϝ�)�]��3�-��]d}lS_�3?
��j�v�e����HiJ{|KX4��~|y�<��%��X%9܉g{蝈��S;�E\����`�B�8g9�"��2���D>�?�t�0 �K���v���'���8��qp�8�6QʩA��3��T멮�NK&�h_���7
�`=C�3C5�D�CzG�cd��sU��,��_�`~��s��c����y)�-zLS``�أ��j�����u*����W��G�@vLC���
��P����]�Ï�X��W�S���ZB��}\�HIԮ��G�\,5~�F��N+���/��9����S��,˗���S[D���唨��`�/����4�[���;cx	@�~�wvy�o�r���B�����/�3z-�K6���}\x�J�mL��q_
����a�5�rD��p�.��X�Ie�}'Ԯtϡ�qGh�ߌ� Nc���o�B�%�D��i��&+FjD����Y�O�}���|�e�E�ٺ��n��"�p0[�����A#�"^asi�J��P�w+9�����@��1*�^G��T���&|2Y 2��1Րy�8Ȝէ�����T�UV�f�&�&��a�x"�{%~�&�Wnn���d��Y�wن�|@9� w�n��4��ܿ4��KN�ij�D!j�>VȢ0�o�8�[	0N�ĝ�x���0�9��N�8��/� �vJW�+��{�z����9]����P�(>HLW7�$&+�E��m���p������|�#�#�d
��FLj� [��~��P%>��9�mpgPچ�u+н�JT��T�>ZO��K��lgi�kO������M��Q�<�_h.@z9c�^���?��ޥ���ES3�e��B#��v�*J�ͨ�ҵ�i+ć�EVA���~��m8)��T,�q�B[�|h�(KAi/�����h�=���i��V�xS��L'v$ށ'iD�:᥻� -�{Ƭ�5Ȑ���E�8��-Y�e��r�K '�b"	3S^�0���n�É	��{�]t�����,�v��#�6��c�"<&z�}�k�3�o*�&ٗۛ~��#Z�Q��!���T�_��+Ͽ.�2��;�$/Q�.?g���ks���M�q�%jΓ�&ԧa���u0	�������=;�� γ��m�J+�o�
����a��p�S�h�2Z�&��`��=��ƥB�I�)*�K�;VbB��w7HG�F�*gb�w��e�=�3�:�G,	�d���[�-G�"xZ�a�ᖽl����ҲI�ۀ�&��t�A��Uxa^a}a�t���1��=jZ��C5ɒz0�F�jY N���j��������^X�1(]�$C9O8h��ǚT#%j��ƀ?�ddH��1��QU$����&w����(�6�K2Xr���}��X�	�ӳ�+��R�M_(_Y?\n��/*�ib���<U�*�ʰ��~�5���޵p�t ��4*���0K��{�c�xl�n�<�J��D�6j�[ۥ�\X�Bb����:�0�}��GVUG�HBL8v��}Tƶt� >��j�s��y��Va\.�UߗQ�������}%��O�c�f�I��^!_v����/0�!��`]�*�o��-z7z� <#͑s�  H�VAj��|0T�Ei«�3��6����<}_7J:�l���)!���<T���j��K"Ū�}@,t,\.�5�t?]���`��h1���(�3?�~���+2N���o�)���3��P6�F�9Z�GFY�����'�gt��3�>|�#Q#%������n]xK�풶5�����%9�D��e�OxnC��K2����f
''r�'�m��Ỵ��42�[����Gr[Y�~j��jY���fv�*�[Q�f�^f#��~B��H۠�`���I���4qP}$�h�i�舀�)_篐�c��T��YasȱB�(�	�F���J�!��h6�a�/$خ�5��1����|�&�Ìa|��(P.X*�x�����yX/��H:��X�YR���
�����
\z���X���k�<A�� �����i��z���*�K�Sw���CMZ�I<�VUl���[�V����%�i�*s������;?��Kl�ב���n��G����4<� z=��F��Y66���Ȣ�`�5������P6�b&~�κ�N���?�� i�ǲ�z ��� �ͫj@R�r��G�A��Nn�5�!�<��q���t������;�I���T��DAM�����f�F9��%˖/��6�����cl��tt�e����G�=6P��'�aJ�{$W=�0�̗BH�N�Ҫޟ�X&x��}�y�i�
2�q�59���,3,�k���hЪ�7Đaي����,>w�wjeT*9��Xˤ���{!�^��݄�
ݤ�9wɀu-�Wy����/M�Mv���pО�W��Z�9� �� ��ku|ጦ>��$@�'*K��T�6dCd���F:�N_�&��ip�=��벘�)]���DA��e�XyFf%&\qK�dOZ��R�7���D��U,��/�+��jz���]R�~7���5�x"Ǔ���З��`�m��ߖ��ʍ�?��onʭ��ɩ옉�"F]a�evJ>1T	ϡ��r;;�&CP�
I�@;�����nf#�k��ZO�N�r���$3J��K�8K
��o��,U�q!�o�/"_g�(&��'��+� 7=-�h�V�������3tr�R2���. i�K�3�/H�p���Ͳ`�U��x.z�/�e�����P#�\�a����B�����x l�z�Q%89����J��~.��OGpAa��<�{Ex���zI����5C��j5��D�KTk骈,&@rqf�W�&1�N�6��bh�2����F��U�8Zy�L��jm��b���U��y�{?%G��!�#h=��uQyXB�o\`@��u���f�lcwb��5)�{���fA�Д���Q{�ـ���Fv�$�ļRi��S��`�ą@�L�X1���ϸ�J���K�PwGK�vi�l�^k�$
�WY��!*�8B\s���(�y��`�Q�+1!ת�����	F�3n����j7���F��Y����m<��@S�mf+�\M#��M��ub�E�S}^��M�#/���\���W
��5Ro5醒�5�Ųv��V�Z�t�I~U@$QED߾��r�����R�8�n�oX=��F�q��n��iX���LȠE#ʾ@F�� _̽-��;�l�s|lle��,�ǱQ;q׵J��$Ï���u�V���	��#PYB�؞�tB��+�}�޳��P+^y%D�^yP����H�.����
�<�+M��TEݦV���u�������	�$_���">7 9�(C�n.���׹7�od�|[�U_�rZo��E&������B_m?�TC|yp�yǗ'�H�P-�/��c�Kmu��:�ۖ �;����$<��/���Ww�oRF��c{rH{���cD��%?��ݷ�����g@j�-vk�Y��J/W����s��a?�U"�G��9��@3��hg �1�Μr���N��Ы�U��"���|/}�bΈSA��3k�j������׳�����*CKPS��L��Xt$��z�ɢ��$�$;�����%Zg}�p�!i��m��X��w�uE��siz�Ԧ���^������rAG�F)������Ĝ*	�l|Pzf�sJ$�A�F4I�#��1�$�S���ӗS�V����e4�����w�v������\�o���T��U-�`=<E�h��('��KMCo��C�2U�3�8�wm�|�m���K��;?�����6�nLʹ��'�EawfO����d���h��x��}@b�3�LQ�O�"��b�:�(�T���nf�ugg�i�C�X5)~�L�3Bt�����N`B��:���Z��c�F /���W�yD�O���^���mۇ>r:�m��Mb,�ۮr2��6FX�L�26zS���ʓ��K��E9ڼ�n���s),	�0�-�E����jܘ�W���;����  �A0�y���*�帖c�i��-��`UF	���?����I2�
D7eJ^���"��Qk����{���}�=� �o��1b�8����O)��*����'h�����邉���\X��vDbN�k��O8�}wC�����͐�����D��	�Mdr���D?��� ���df����%�=�T�[��b�"ݸ�ձ��$����J���j�d�f�Q dư�V�	cG����ֶSm������0y�6e�%;�_MQ�R{��b��;�)鈪O��#�	��a�LV��:�`{\�gz��j=y�)F�R�+����g1�J����#Ou�=���cQ���+�������E�Ë�h�1Ğ1/�q�"�\m��V��Y&�uJ?���*���S�P0�͘�-�أ>@ ���A$����2���ę�(���S,6��ΰ����-f����y���uq�
I�۸�;9�}��43	���?�)�{*a`$Z&w�&�g[�u����~E�tj���Z�iAP#��J�&Ga��*oW�����)��8�_n*f�=K��&��P��e�˓&k<�'Od�Ÿ�s3���t��Fx9��5�i#S�%<>�0�a��;,6�'�,��+�(3�:l�Sی\\����1_e�0S�àT`�J�N� ���Vglƹ#�]t($Po[�՘���x:��셚Ys�`Y�ʕ�]�KNo�v�Le$`��-��ي���O��翷9��.�\6���ݬ�W=����UP��Io�ѡ�B���T��5rl܇���֠��!�Qrι��&�V���*�j�u�A�?���_h��N�P�� &���Q��9*��D��U�a��e2<�-�5d����
��#s�!`Y�fjCn������ gD����������n�	_ #!��p/t&0�E-R��_�K"��[�*��+� �
}��P�����z��2է��(�t�����0��Ejc�EW�wX�WF*�1,O�N��m��b��a�t>׆Wu����/⾫�����	������y��*&Z��fVT$o���ߴ�~>��r�#~�݊^��y��(��v�M�k���H��D���=��j�V�L㎓
�oM�j��8~�m��]W�%�;[�ŝ�c����~F(�ʸ�A�iC��K�th���;1�`q�Jҷg♡�9������(e �-��ZSx07br$p��ؐ4����3��=��yr&�s�d�4?�e�s���e�2��<�;��w­1��%-��Ԫ�w��� ��R�
�������B����~v��B��4o��l9�9]be��o+�{�3VP�!֥�1�_ �~[SP��F���$\�|*�������O�:1L�y�
��3������nrHq'k��D�_si,f���2DiJۊ�'0��Ӎ�Mq ف潡MvE6�qW��q�&z��}+5<Q/;��E�E:�~uݘ�1o��� ,�c⇿�����0�ڛ�A�B �&%�p�X�]x�<f������� ��7� ���҇�!V~��q�z ��'}��cǑ�AO�ӫ��DH:��<�}Yϲ���S���5w����n=o'������'37e���N_Qjɾ5dά��S��~	#�T}?K`P����k�zxt�a\3�0��.
"��,��������-��ab��=���!�9��eԎ�u�Xx��@4�g��`0]���vtA������|�s��*ȝ�1Kة�s� oO(�/k�� *R�p����̨�2&(E�j}Y/<�V�ƕ3h���B7���ǈ�i���3c]������iL�0�,r3߯5�jzKX� ���85�č��h%=�?k<lb�^2�/<?]'�ה��iL�`ֺ�s��۪a9�A��@.b�oM�n�q$Ƣ�qh��G�Ӌ=ȋ2���g�ň�g.~R+��r��8G|�x}bn�.���q�u�7ρ`nO=Ǧ�+��̟�Ɇ!�y�"[;� ��x��TV��Ls�g����&� ¾T�'aN�}����2E���98��c�^�O;JD+�Ļ�Ĝn�jF��c��\Q X�k3�8���I
���VR�܄�f�4�ͅ~7}ǭ�[J�� �`��m-U�DQ�vI�E�6~�~.�v���o"'�ʡ�d�2b�~a�pA҄{��"��s�}����?���qt:Z���׍p��Bck�X&�a"������d��u�b�2�tڕQ�����+���}�^b�仈ހ|(b���y���0�F�h*����"�#��}ڍr1TP�/�
�"W�=�"<Խ&�1�������Y�@��(I{�gc�υZ�����N���"g�l��p�5��qh���\� �s"?k{]��+�Y�@�Yu��3�p߃��P�4N����"�DbK����딩��I�z��@�ӛ5MQv5�fu����C�U��y~h�A��2d^��xl���d.�/��E���w�u�
r9�;Ӳ6N~g���Gmvm-$0cY���hP%m�$��Gdg2��eϺ�wX�`��]u�o�d�;�����A�x%G��=#���"ɔ��Y�p�]���Vs��fю
S��4�ȟ9���w�6�D�H����{�\��g�q�Ő>��ؾ&6%�y�.���zM(e�s3b�cQ@�HZ&|��S,�r�Õp%f�=�?3P+�ZP(LL�M3�_D.�h��5+���9��yƀ�;jk�o5_�x��Z�c��;< q�aJm��GÊ��&�ks�*?Ӂ.�L"%}AI졆�&T����[��!�e�ZLA�o�\odv7�̑�|W�T�u���14�T�o#���3d~)����OQǜ���.q�?��mZ�=�1�~@T.��`�7s��e�I�|�|6�[���8�l�e�DP�̕�"�� 'g$�wϡ�	 h%����=�Q��l�ՉT�A�^&�Ѕ�Q����HiFs�: �4Xl�,=��n �VCd��YR�˳+%�G�BB�_�%q��߉'.�g@U9j�0����+�u0�Y�A�X�E�Tw!��%���zK�X�8�Y���r!�"R����i�2}d3«# ������8V�W�&�L���:�:��;Y��s �'����
�`r�`SR�nE1��w'Z(��w�6�	n	t(���7-	�Uց[���̏�Z��2�f��\!��c ��D���ڬ>�  C�4Y�,]��LՕ^�<����L�R�huIֺ�S���p��(�z�u�b�>WF�n`+(v�`�pW���v��Q��) '�n|4i87�NO�	�,�2R�g�9���4:��@��^rq^�A7J�3��L�KDfܖW�j�
�1�V����bm�\٠L�_@1��7�v+�HzB�w�PFMw�6Q�Ŭ�'����D� ;p.*�
ћ訦��q��;)����`߳L"�3%V����u��`��tf%���\�rt��e�����֕x��i��˅�[�:?�m��*�~$'�#5L���d6���;䡋��
�|��B5��N�V@֛�;��ٓfO\�54�(�r/ dfڞ;��v�q��晍��6��D\�*(~o%y:�u�Q�o	�8|]�፬ߕP������<|�-O"0�����71L"75/�ay�F��D�yx��Jg���q�ѣ z�}���`WΞ}�TG�Ӕ~�X��T^^�@HM�jKzLEt�OPj ��!Vc}�`��:�����?�\��g�`����\x�w(?t��}���r�s2�����X��6�o�D���B4�h �@�PM�z���ڏ�>lI�(�Oy7BШ{p�O���O�[7B�	����*�b����_�O�Gq��aJx��ݣ����u|��]I��^�����������U�t��)��Quڮ:}�c2𲟶r�����7�oj���� d�o���\T��>�u�;/����<�=�@�J�v�ĂډK4*���.I�.���}u��n9Á[�f��Zl)�Op� �8�Z���RMb���+�gO&�C�fI@�-9��}t}�V�d�Br9��3���V�b�it��}����}�1�6g���Vʲ�2)r����	���;Z��a����(J�u�r��W+��Ć��Z�{{�6����g�k����K*S  �(�[����bh�ɪb��16�0EI8oCV��$�*�"dɡ0DI$~��f�EE��f�G���T�q�:l٬�	SW���s�h5�e1��>�&`YK���1�Mp�u�I���g�&�N��.�H!/�He��w����i�;1�ٽ�b5���f+Kl���JX(����u��IiC~q5�⪊���sL�6��P"i�^������
�����l�@eD��Q�W�kT�.��)�	�D����aZ%���侜�
�Zz���<���.+��%�B������=�q��p�4��I|p���`�+L\!u��
�Id㗒 ]l�~�ks��(e�tɟZM�Зe:L�ob Q�"<J�w`�h���ၳ��b�}p��'�0_�J��(M��mlo�	h��cO9�W��(g�l��|f�k�uG.��0�0z�[�%�@�n�0�����#�$���!9B�p������}M:����96u�!g��j����J<��̋3��bN�{>��Hz9P9��!��k>(�@����ߚas��%���&�o�"����p[#��:���ϻ��<�a�{�"���5�(1]̱�q�T�[#����`b4r�G�_�Y�A� )����f��ګœ4�h�z��3�SW$�:���E+<���ˀ�9�1 o�^�T6�'���R�G`��h��VB��Z�a�n�bhi&��G��O�=����mr���ޙ�o�5wP�,�dV�%x���S-F{�	�'��.�(������.�#�x~eǢ�>�B�=�d�����JRz98`O3NN�>^r��;�~�s�+�D�d�
��8��Vp�۟%�3y_��!8-M���Ƿ�e�TkoiU�w�J>���|
���o$����}�]��\wK��l$l	�h�i��o	f'����~?v��8{R���U�:k�6(�%/*�ZA̹�H��Ӱc�:Q�����@��̟�j~+��l�(��]~ܼB�~��������z0�{���Cn����D&'!���.���#K
,4���-���Mڭ<��Q�不¸O�ja��蜻�gI�@=��[�I�� H��]��0V +�����5&��<$x�C���٣�X�&�f��j�_3��Y����
Z��&dt	=����Z�����N�Y��ԕ���O�W��j�Ɋ���g��_�FU�(�����	��\�R����4��2
��Y'\�x!��y�F׿��>�{r�b4~'kQy%�I�He�\�C������(̾ap�830�g�ŤsPG݌!�Y늸O�}�'2v��!"�ϻ���-�V�j��<m"O�^�"�H@�DA�����g(Q�F�m��K����1���ؑ��j�H��0�X%bK�A���,ҳ8ح����B"��j3��cĭe��b��n��_�d�dJ�/�����	��+NO��cx���]J�?��t|�=�R�踚d"x��I4s�h3�����r0w�����Uy�l"bgZ��%֘��B�4�ۮ��c͂Bg���U#N�CX/�F���@Wne�%
�5�5�0�݉�]]*2n��E%s��=���m��`�;٪d�i����g7%���G����]�V��8.E]�����lM�gc{��ݪذ�6"{f���,�u{���=��(Ĕ4Vs�%�z�b�<~��|8?A���R���Om֑�y���>�����J��\�C����A����Fe��y!�KR��gzR�`n�m��\u�c�I�l.����l�X���<�����@���N�(5{n�;
eJ�]��I V�l��e��X������}jg�KJ]��7��{ 5��`���)����B�]Snk�t�lԁx{�]�
�E���?�9bY`�nO�Q��T#������a���b��ӞK�%$簸�QG��/�{�Щ��*I�qm�n;�h/nt���RYX>�M�����S��s_�u`���܁�����"B�lW�a�?I=�_ҕ��T22F���A����@��)˚��ϣ �Z�����U�d*���w���b��� ���(S�9?a9V���6��s[YT���`�f�lX=0�S�L��~z�è��S:���X�`��6�l��F=�.qR��^n�rCw����|�L�����$i�Rn��_䣉���)F_
p�9W�O1�lEb#��H�$��(�䰱�7��8�'��e#G�T�ݕ+�X��)׾�0����[�
R<��d��� g��J��8s��ȴҺ~H��m ETl���.���}N���}ȱ0�V1�^ε})�<Uj��V����1�ߝŮ��.r��-�ֿ�w5��R���!�2����I	�O�5�w�O�=N�c�4<�ac�<1!H�ޜjɪcʨ3���R#
��j�	�9Ly-R���%�p�>��	ѵ�g�>KЈ�0���~��q��O��jM�J�93U|v3/�p� ֎K��{�R�HKӇ�!27����G� d���k,�WM�:o��Z��(����*��W1.S ������$a�FRa��O�a
ƱԴA%P��L�М#��,eb�b�)`@�d�5�}`9-ۿ|Z"�@o#�Ɨ����g:�[��z���ȁ\8Z�"��Y襷d��(�*0�㷛_��1�E��=��w�U�Rީe�ʠð�ﵡ�2X�5M��|��w�|X�mn�?_����*( ���i�<���NW�{C����o&�h"���C����fE���Sf(�:W!�@����o�-�<�s����ɽ�\��t��`����-��Z��{h���2�P��S��)�4`^�I�L���
2�Ԏ8R��?�^�u.�F�E��XH&� d�_9og('X�j�gR�K%�9�����V�C������ZF������)���V3�7���1�q�eB��>֛���W~���i�ȕ&,�,� N�/�:�3��Ƴ~v(������*�YN8��U���\�w!�j�9 ������>�������z�>Yӵ&���&���f^�χ��cϬM��pO��@4��ል��{#Β���O�Wt|�f�O����J�q57�SY��s�z�$���Iٛ���B,:F�U�֘-�������tR��s��H�`���ػ+����;��*A*g�@�?�m��@��بX��8v���H���F��¹6�3]Ȟғpg��$��=$
��U���0��:���y�o� �~#�y��f�P�w�j�w&�b}��t��S»,�(�LNa�Ė-�r�4���!�������e2v�6:�������+;O-T��^�i1e�9�Z���R,�?�Ň�'7�p��!�0��%�7�k�����_n&��TR{�Wv��׸M��E�Dg��i���$����=�i�M�����f8�c����w���R��b��U�F�(e��h�y<�4�f#`�%?�~J͂�
��D< ��5���OQ}����Vƍ9�b��&�+�&�L��7���e��{�����U&3E���nhB�y��
���2�*�`ie���M�bz��E��.�j~�';�ޚ�+����Wf1���\B������cP(:��,�6dq����݁AB;�CѤbh�0����
S#M��]�����@�{�NqL�/�{w9������t<���2L���/#�끁��h=�^/���$�oz���v!��܂/ �虊��a��;rtc��R:�f}/zt������aQs)Vm��~O<5uQ�����q���X2�i�т�Y$�d-�t�`�z�w<�?jz����w���lp ����I9�����ǽ�BO1��<����1*���A��D+��o`R׹� }�2��ٳaL@�Yd�giU�#b�:V 7X�8�z��K����b�*s=���o��X��Φ^���nO�eN?��&�ث;��^Wͤ�6��☸��'�8~{�-�D����j`2��n˗��Gi?���?�@�L��mV)v�d'�aT� ����5z��l��s{sq�8��,�Pq!s�
��I1ri����w`e����������c�����Q{H���c�O���GF�0o�Ė�6�@��)������$3І;�l6*��M�����Ka(�g��,b����=��J�G�֕o��z���|���+D����nmH�n^��'t�>�85���nV(��*��d��	�c��dm^��9�<�<�0�Y�Xj���Ҡ�5���f�w�4̔�}Z�� i�R4��US��$���~���'ru���Ep:�%䣃�}l��/�ɦ������K9]�����_8{ ?s�U뀕��k�m�I2l)��] q���(T�8���PM���$�O�P� yr}���53��œi�,陞��v�I0�$��)�!N�
��J���_n�Nc*��hނ���T�}��� �qg�W��о�+BtT����܀�f��x6�-�
pD��+V�\'<��:����%xA��R2��-Y�D�7ׁ肓�w��[����qη���9�>ڋ�0���:�轹�'B^<s�	���Y�_��4��� Y�xJ�x^�䡞6�m�ɾ|��ǍS��N~�M�z�
��
]��3kg�n޺��o�No�|Fc���0@��6�ˊ��R�6\�{�U�eU$�����2�4��um�KO�%d�St#]N�)�9+ t��B3Ю6\��[���{�ԏw��B� �9yl����Bo�\�1���8Q�Q����?�?�O�Zn��`%u,A���1�
�߾u�����y�ʔ��MH�>0q)FΒF���� Z%��v<%Z��QU��FۆQ�ե
�"Jh���E���7���f��9���Ya<Ӑ�+7����_�W�aMƼ��*��%�⢁�vSȘ�������q�C��S@&��{�2_>dEw��ж~.ҍ����HR\�͖��,��E9|�q�ǲ 6�'$Q���I̓�a�b�"���/]P���u����^$���w��#<8ٹ"�T'�C[ՠ�#a�J��'`R���fΪKAt�v�Ic����9I��Q�7'U��!��P,���+�y�]���/����۠:�Aߡ�
w�]m��,�/Ͼe�5�naP��q�%��GJg�g0{��0Y=v'"��N1im��� � �*TZ(�N)SCy_��-���g��.f�����G��0h�Ld�k��tǉ|�/�=?	�b��+AY�9��CPq���@�S%�X����y��T�3BL;���>��~�X]I��It�,}k��%���#0�y���^�B���n}���bZ��P��?�ŷ	��\�/���r%YL�N�%v�7f�<��S����N٘�j}���OH�"��|��8�b`A:_4�m�Kr�d(])�|~u��w�	汫.i�;8�%�<{f�f2�.)HVXXY��ZK:��Ǡ��>gӉ�����vF��ykJ�U.6��醸��`C�{�A��-�(:�� ێAo�U�y�}n�ʒ�˶"��z:���.�]Yӯ�EKx�	blF��N��J%= y$�-�dL�8V����gl�s��k�R�����< /�$����f��s=��l'�W�!����Ԩ���3J���f\8%)ٔS��h�5c4$�4��e5�e��cU�|�Q$��!B>Ԣ"L���a���w�W�]�O�Q:L,�	C�y��e#
L\��q�e�"(�����Z�g���R-5��s�"�}bj��SIY�i%�#M�]�No_�|�y~��϶	�M�Ĭ���b=�N,�1�-~�� :�'��e o��V�*@e�-a�bɘ�45�A�f�WӦ�?����L���~d��c<������vF�'��ՙ���/-�_������=L�����ti���:��	������� ��x�T]���paE;$K�|���a�F���̄z��f�;'( ;X����Θ�;}ung�jb�V���^y��x�� E�&>7���@�����$����S�5-d�'�>�T�K_�E�i��Hh���4%�~B1s�n�2�Z�qi(1S�-����2�'P]�F����>�#���C���� �Ij��e����C�/������~�e:f�C���$�tf�Fp��~'�<�nՂ?����Q<�L1�x���@����e��N<�M����Q��(��w����v��{<�C!��?�~������Ϣ�#X����X��ӂ�wc�!�3kѩ +�}�V;�kd�	�ӃI�Fo�����ӟR����֣"ɨ��w�1a��j��֛�{I�f��0ٍ�KxZ���N4G������ϮX�M��Σ��M�zKhW�M@�*�Z��U_*�[.��G�mp`��ok�f3}x��3Z��f��| >���r���d����&�вW�8t�	�
P������> ź���xt�ڲF:���o�˸$�c_n�m8/��̨{z�0tIQe�>��;�\6Aiz��|��#z�'vTW��l�'�U���f'f4�]owT���<4���#.��Rhb<ήCd�D6t����q��;Օ����<���~r�;�v�>�����D�a�"�=|��?���Dci .����jMH�ޔl}�F�٧e5�oھ$�U�Z2��|H	�+HZM	R=Xszr�$ǂPp���bF��'�a����`8v�+;�"2�(��4
S����:%�6�,g:Ă�9�H�~��o�=�e�C-N���̲����v�{�����=�E�a>�&��G�S��ᔟ��;��`y�9�c)���;�3���iS��3/�4����MWVbtq\6X5�ٕ@����G�T'u	g4�zO#��ω�PC%O��&�>�qt<��P��wB���b D�#�����AkCvŀ�2)΢īB�uȟ'f��iM^]��iVX��'��n��
+���_��bW�Hn^�2�f� �C+�Uq�����P�4����$�J{��|*I O9H�vY`��`�e�Tv�}*�I��{y ���є� �����_�rْ�<)��;�rL�)�	�/w�Ŵ�6a��:�+wf*ȯ�� �FF]?�����@L�������i�#Z�~.�Q����bT������C�f���"e�[�BY
�c�����G j���)=�iVC���7Gf��]ZX�pkE����^P  ����ӣ��F��}䌽5�Up|j,�~�a��3����k*Y�q�o2Ւ�V�UT��௲��f^���ǙP�� ��y��,��L�ǹã}x�B��Aa������dX \�vl�F�ZDʄ��\�[���6l��٩;ϖ�us�W�O����o��4`�m.��p�tyo�{~;���=db:�J�L��ۤ_>U~㱵��!����������Zg[6����`�	6f�Ȍ�wF?U�M���d91�2��Y���bPMj�%z�q�䩡33�`��'��ۃG��}�(�ݶ;ʭY�,s�/7��]hr�M$���/K>Ҕ���d��E�T���w�p��M&<f�H�M���{(Ȕņ�cR�`:�|Nn����5����vX{;'���vl�=DY�.F�&:���C�i��/.KMN����v��JH��Ӛs��]U��	6��M�o.J<����8!dV�����C��|�*J"���(���-��g)�ᙇ�_���ǜ���ǃ`�"5r���k�0煝  E�= �k��ҜB��p�g��5�}��pKx=u�H˨�hf6�I��Z�9הv�Sԋ-,;�U���D��O���[Ud7�p��B�3Y���9|`���E1YB����
ͥ�Y�HK��X�5s,c�`���kkxw���֢���ozV��Ã�c��9���� a��"1��`1��H� �<.
]�-�B��	���g��bHj>��=�4�=0Na����Y�֭+��]��8�4���[ǋ_ +� �����Yʁ6����ѵ��L0#��v��AX{b�tH��s�,(df�)�T��Օ�����"=� rbhm��cU�\E�F���O���}X��<Yz�ֵh��n���7�
k-Y��ޖa�-�I��k�	>~�*�m�j�R�qS��Et\�%C������@���N@}$*�������h<���R	L3_�\a�?�Y��Iؑ�O\	M�bC �4������Ѽ��!�Ip5 �mO������i��״��  ���F�<F�d�������R��～$���'��߆�J,wza���o²c���	�n"O������ąc��ɾ�z��%�S6Jp-
���6!���'(Dw�$�P�����Na�{����m��<j-����I��%}�0��r�z� ,5� =
��Lx����UD�qC�1҉�_
"�b�&)��]LGFd��}��2���ə\˲�$t�������G ��P09�f��O�>��a������?��&(�ء�(�������D[|&��Ԥ샭�Z�� �e���m��!�CĶ�
�����%K7�ܵ�%�o�/*��m�Dր ��Pj�BZ)�����IM��?L����-�IV��c��P+l��W�ه������7H�&_c���7������T����	6�A�g/����;du�Cz)���y'�"]\}�g./~|<E�#u�e��~���?��k˞*�򹹣+	'�ĝ|_��w���˂�1��;%���q�D�7ݫ״"j������!�j�pn��n5��Ь�V��ƕ��{D�bJNC��eu[�� 'tRĶ­��1	H�4h���0ɠԯ�Fv0W%Ο�%����Q���u�� L:n�Y�nd�n<�d��� %xD�u���%����gO��㊆6��	�QUw�(Hr�p +�.5�_�`�#�� �仫�{B.�'����V�wZ~�T�$�Q<��c���e�bk�q�F-�(5��s�cp/�|�gS ��ɶV��8u�7}g[ǀ!�Ł�5��yG�Ha��휲��`�oa1J���:2`���@�enNK`?��>�:"'p���S����.޳*��g.�	�f� �3�t����=�3$�|���*УngAP8��'��� �nU�Z��^�ã�����/X�e����a�w�#kF�
�����.�,"M/F,"<!�>�+�)�+M�nta ��M�G�'��V���#ko�]s����������]�s���@�)�G�µ���d1�C��+�䍋�����M�a�����,�=E�Z1xx�������3!*=����K�VL'�.tW�4�'CPҀ�{��a7���%� �h����)�����q+;h�>��[f��&����!/����@�����S�c����y��F�z������_�^Uz0�ɖ0J�خ�ː�h1�yTZ���<wXhUUʴ�ǈ1-�[��� tì�����X�v��ڌ�Z��[}3���y	�|�p]�K��J�h���a� �4�O�"\�ɥe���6���s�AJ��ǳ�D�,gZ�> ��~�?jKl�g��ÄK� @S�-9�2��1��b���y�ԙ)s�c���ka���%��쌡�18�:E��A�A��J�q��h�����[��g�8��.p�T�^�Z���l��_� wDT}Tɟ��0b��r��J����!C����-[��=z�og��/�,l}�TU��Ak����a���ef��h�7u��XFhf��k���,aO^~�Ҿ<[���� ��Q��&�Tyc�Y3�N�mF/�pY>��.&đ�@��r�w��ui���ے�E��A�Cb�2S����1�R�W��G9�f�On�G3�W�uR���o$*�`(Ո.�e25I������@6>�r$�6�@b��ލk��@ �&��L��0`�ej�7���.�4����E�d.�m�e��0m;�S��!E$�'��_�x��ۅ}cE���&g����=����������3WI~p~���"�n��;o��ǯ���n�+�W�[ca /��k�?��:b�w6׆�JAc���AȳPן�>J�`�SC�dӤ6=f�~����Cp:[W��3��M��w�o���3�������-O��d�Z��ܯGس­��Z�eN��Db��$�J�=P�7f�68��d�/�
r�M��ME�M�*��z��IC���H�9��֮<Һ�];YU"����޲x�N��3-kr���(���+�Û��]�-����`(?�l\3|	��k�3І�rm�7��e�ν@޽Ǧ�� b�O�{�gn3�n�4G��Vg e��l2a�In*~��'O�9˳�c�\���Σ&�_���ߠ�Pc&�`�#�3*rc�_��Éz$�[����_q�)^��hmQ_z�khh-k^V�&X^�8uCςQ(�J񒲞D�;#@����K:2y�X�=b�r�PlJՕ�ז(	�����+o[��8������,����˛��w���I���XV*��55M��C� �]�³M@z�Ͼ��b!������$�x�e���9�����&�*y��^>�@��:& �>1���ٳ������r�ó6&��N�e�� ׶@g��@{�S��\���#�fi�T�2���gV�3x�/�����(�`�vB~��q���+��Q�X˷��ˮ7G����I�ᖆ�l�A<<�8�W���yi])?���&�B�z����Z�o����ѾȻ�`��;���L��*� 3��T�UEe��)�L{f�$�G��N���
^����trjՁK��%'���{�jf6��$?~knZݮ��zC��/X}k�0JÈE�\t�?��S˰�Cc

>I�	؁�R�42z�X�9�Q��ѹ �	��%��q�7�䧗�f]`*���c�^Xֽ��];l�O�E�"G��_"�?�̮E�xBr���O�6`�Kip�VK?���r�@��$��Dh�JPZ��.�I L��W���
���'��z) ��00��S��Nh�����p�gvEp�n�X��V_];l��e{�X��7�� I�i�p�T�"��*4��E���Z�?���l"����.�Y��f8G��l�9Sp4q�((��KB�ƴ���Fū(���3T�N9��*A��w��-��J/��6��O��|'\)�9�o�>��r�d���ةB�ƣ��U�]�TX�E�h'��F�c�L�W�[��[68��U�	�~���5Bá��P��q������F�نa#��X���o�[�m�&8P7�0��ڑʪ��C��J��%+�W�,@D��1̱��ڼ�������F�\&�I��󓺜�g��1�b�N�����(�'d�ʗO&y�Q��/�<2�nS���L+ʟ��j?�ɼ�n����䬨v	
KU&�6>{��N�NEٴm�W�7�흃m?0��㙰fF���D�����q��V�i�2[2bDN�7���H��^DV3�� ��"H��_ ݂6���#)E��j�潕���Oz� ~�;|�����)�'�aF�.S����������mm���M�F�@��rh9�нi���Ҙy̪x��y�%Zl'�r��=H�y�dS�(�rS=�e&/��+�J�?Ze\EU�.�t��:H���t
���\2�z �@ c������}�+lT�}~,���w�[�)�mx}����Va�d�k{3���',L�P�)X�A�=�+Y�����E�c�6�U����~��M�Մ�����`�`G�0�ψo�; �v�\��2�L?������~�q�R"UQ������
?�N�glD_�_�	cw�&7���K]�y8j�
0�G��z�cbU�ٕ���Yy��ˡ�M�:��1��y����pR���M>&@�7��LboA�U�g�A��>[�i@f�u�Ћ<T�"8�]A�+Ɂ�
�����{�)�`]_!|�a=e�R�T<OJ�G�jP�O�dx��5����,��� �aL���y�b�/�H���,K �mg$�x��
Y@�m����!�F(錫���p�n@��L�6���@/��Z��vH8����YT���ft\U��E]�, �f�����Z.�>Hց s����)�&ڗ%B��^���p�W%tO�:�0 m�K�䚁�g���鷞u[�˖]=A�+��C��2�}# ��2��' aZ�JY���2{�jF|���#{�^��[�	D���討�ehك�,�DEC�häX/6��$H0����yG�ix\HS>c"���A�7<yP�A���9ͥ�����d7��b%�l����T�������+��p�-@V��]�!HN��"�]I�#��3�
�{��OAc��k�VE{E����Af����9c&�z�:k��}C���f�]�f����>sb��C��ś}$�i������9�p_܊��׆k�TQ6���xI��p}�J�-L����B���ܴTr��#�g,B;e4�N�[�-���.s�JHdz����v�oyr֜ʚ��� �n�`J"���4{*�x���6�Al�G�XK8�Ŝ΄���+N���M����3M��W��p�DNf�#x=��l�7�TTĒ�{_��djc�g�q���@�m����	`*T�õd��_N�Sl���{�g@��}aG���J����YfN~�a-��恿��}T��r9��Xٽd�$�xtkw>KZ�/�U6��a���(H�l��I,@��N���m�U�6L÷�����J\���?F|Ě`������r�P�.��}40"�xǠ��^[9��.��4'����� �X��(�u6������ݍ��q��d+R���:��PX�.O}��s/a�R�C�%P�Ö�e��c�����U��f���w����A^�K#�E�0�rx�UL^���-}����?m�$���3�������.���;%Bt_x�m���C��r�h���F�@�G҆�_�?�-��I �Hß	��6�(��k��\����]�@�l}�O�R�__UZ1�������"
r�$̙`���T*7x\]+"���>O�2k��d+�0C/�S,L>�N���c�N$����\�o��Re�'��p;e[݆� ?,1�/��#�����WY��ƃ�j�{�5�6K��oD�e9�'e�3]��d$/n���3f&����z	���f� ẊHL,9��⸈��c�e痬�M������՗>��$���TKyUu%G��hNj��$������(W@�~�%-/���b���1�����~ȅ�S�̇-�]���/dT���W�`��&��yp���o$d�w��W�n�[Pi5���r0$/�-�����P?>V�.�r�Rs��6~*[�Α�-��k�J��̼��z樢��#�t��\�&��U�|�ym$��͡����Ӕ��ѭ��Žx��)�_���a�9�NΑ��O����n��;��i�k$2\�k��0É�r- C"���sl�/���XbJ;�|�P��0w�߰�$�-	P^G���� ��JH�}Nu�e�'1>����酖1���G���߂�*O�C?�p�=.�?��[~\WgHb>�1�@]�J'd����΀13��L��ݤD�b��`=��>��r��v%��'��k��J�X3�pf��`U��)�),�;�p��Uû�b���Ԡ�`�$��"x�/)�]u���$n~,�"wX��R�1i�Z��Iu�^n^���Ba
)��;S(�2�����|��1hF�V�{\������Ŷoq��`9����*� c���{W|܇wA�Y�8,x�g���*�&��Q��◅���~�)<5%M�o�{�?���P�[@N$:��^�</2�!Ǭ�[�[1Ef�)�T�o���W r<,��˽lا�u������봅�M�Hٰ��x{�<b�������G�|ϔ�.�L�#>T��J"!�]��Hv7�ll�p�>���*����͙w8%P�҈�.���Y�_�#S��Q�S ��Yp�Q�s%�B�Y%2s�/K��B�ԎRN`���	�z�Q�� �̕v�rf6�m�k�9���q�Miz��{P��2T��K��.O3*�`�4���͟�+@u�#�;��v���7D�}�C��/�F�i��;�3g�߹�� ��ZN Bo�^X��3��3�Nu[�έR[�<=#��`Ĺ�]*��d�\	���P�E�곭ww!5:!�;թ�+*����� ����2�WrKt���@W}�c�jAj��?�����Ҭ��RJ�9l-��n&�e�E��c�-57�q���`�1�4�G��H���Q&ꏧ[@u�h���2�*m�&�ۍ:�~5~<��|������:&����˲��@|x?�@#KG�zx�� 0�b�1D*9���f���@4��?���`M�j~�7:jU�Z��zt�|b_�A9��8D��N����ӉINu4 �7�j�%�B��f#� x�y�h���q/������"�N9-����@g�|>�����J�����Ug]qtY�NM�W�Y}OZ��T�Vb]_��H��Pu��U�'�_�+ ����9�,B���Ϥ%p�c�;,�s��,�a\���'dN���׎JwJ����8iK=����_SÚ��+�����p
�.�����+�*iMh|I�p�Y���X��i�����6�O�[rq����`Y�g�mi7�qC]2���Mn�!e�3��^�L4� qn�DJ;h�Dm��D
��/���DK�5����.���tņK̰�J׳��͙+HI*/����I�V�F"�kF�1�%J�r���X�������5]�*Ϗ{.����c~Q�vI��Y�ɀ�"�3�(/Ō�:�� �
����zYh��.Y;ds/P�i�B��~z�=Ŗ��몿&�&F-^�H���!8Å��A�ة��L?G�*T����bi��cq�6�"sۺ�Eb䴚���W���0|���դ>T��<�ѯ�/�������qݝ�Tj�����V1��{	�h|���\o:��m�>���q|�k�s��e�zPՊЗ��zp��z��F'����uCP�xZ-Zbq���j6��.�&�_z��Q(D�<1��o:?i�8��b_�o�l�`Fi_x�$�TNtD�N.9�3a� y���dX]ߡ��3��H�p{p�W�埵��0 D��ox�9���g{�i�Glu�I ؏1Ġ���e�]e�N�<�x�~*�Ka��0wS5�6Rr�Z�8{�����:�u��t*��.�_��T��
*�|�U�n/�e�{?�ƙ�g���p�j�0���U�"�_�h�iW0�C�F�-�5�#�ܶU�Y���G�UZ�(`#��h3I>	�G���x�c�I��_O��sZ���HB�H�kZ��/Ic��}�>aE�M ~��m�M�e��G����r�H���4maV�Ghwt{VΠ�7��'��AV�LF�'��c\�s��kƍ$՚�$./EW�+�
��Q �QAʶ/#�41]AD�ܝ>*P����Ӗ�����OE�m=��6��X4�q�@��$���x�e�ũ��؋��b8��]Z'��I鿵���t�u��-����{3$v}֏ϖE�v��ʬ�%{@ 28	y��[���b��S����C�5�v���͏V!J	�C�l2h��>���\�@�#u��\Y�E$�B��h��<�5B�0c�}�sW�e0��:;@*���)�7õhٚ�������c��\�[`=W�.�2�>¸F���Jݚ��U�I�E�'Q�����G��]����L5-9����ȡ���g*�1����7[з5�9�e,�ٵ{sI{^�e���w�hje��-�j�5����a��4d��h=G���b5�l=Km��aN\8=G��nҰ�����Ir��SX5��ѐ�`��J���� ���QK�A�z�`��&���{gxZt�^��Iz���tȅ�#\�aY"�Vu�ҿÑ6B4"e1��,�:5Ƈ�'QpU������T�H
WLq�t��;�W���e9��6�;�l(fD��H�������巅v��mR���c���Au�l�83�y}:�w��"d�pz�׈�k��{������!�@�8.��C�i�3/y���1�v��ȍ^k�˚48.&xONu�A��"�M�c��iFڂ��*,�R)0y�#���:�)�Bm�mEu���$Ϣ��b\�p�1{h���c��O�H��B.uJ�whǂ�a�oW�D�o�o�PC~��8fpI��8�41��g��-7�r��gSoF��K�&S�����q���a���`�m���0�r���Y�p,W��68���^2ggJ�!)Ogȣr�P٬� N4M��_�W���~k#j"�LCvϾR&R�6����$�h>��@� �0����O��=_WN���h7g@����U$T8����/G������]?Z �{��AW%�H��W��"�BrO�}������L�kߪ�MX^p��j��^C��vo��__�-k/Xȳ��Ǘ�3�����Pܼ%�N^�ijD��w����/�٧�H���.P��1F��^u�1��50����:o	��p����7[�b93�a��5�!�=�����ѐ
F}�zc9�	y�9��I��*�99��3���'ׁ��S;�:q�0��(�Tp�����@W՘
�!�b�|�k�6z�>ϐ�Q�[?�Ul���A�A����UGpܦ�+=�Ki͋��4���u�'l���&IV��%#�T	�ǹ�Mްށ��u�j87�"�G���\(���d1{��jG�4i([�A�CM���t���mp��:W�X�b� /���.&�1�kϴ;��Q1�QjM�(��la�H֙Q⸰.X�]�Ȕ���5�Ƙ���)V��$:���]L��P��[�פ�*�u�V�k�s�)��%��f��c`�����|���-��`k�QM�j��G����i��$�:.	�E���l��j~k2<uګ
	�����JCdn��b�.�����,�e�h���?Q��A_ȝ��}N�0z��I��nb��Z*lL�����|�,�mN��|�����	C��J΢&�F�#B �|��V!J�t�
��j����U����Ć�}����;h�A�ɽ7̣WN����%P
R��Sd�:%ܷm�눎��2�
��)�>ʔ�
u��S�����X��Y���^v�E�5��yj�Θ�H�s���8��[��~\���m��\P%1e�gWp9��>n����O�J�?A�ֻY.��_ jI
R琥q��܌x<Fs�	�v�+tX�Q U���<+��7�юo�G5a��m;����̴�?� ɘRO o�1��1�u+Beނ2�\�v*�B�A���Vdwa�`֐' ���#N�v��U�T|�n��s�R��S7�gd�,M�j}H����Mŷ����-�@�냾����O$����5��T!Xg��͍r��Qy
�of2H��^y䆂ta�$4��Ġ�j<x�U��#u�Y]f[�(j�_O��	Ip?I� ��%�n�Q��lk��T�?f0U�?挰�����|�Q�ľmo"���}�^A�0mm�أ�M�7%ݵbż�泛$l`�U)q�;�jz>�s���(���og�B����a�@�hl�I � �����n��.]��'�!]U�r���Z}B#4�t��綥ww�m�9��A�)�7��s]�zmt�;q9!���kb�z�*Lu���y�>���e�{S��U|k�=��t��:�9��_�4SqQ&�l���
��K��2g8"܂b�<��*a} kf�i��ì;M � ��μ-Q�[>��T��ؾ�z��°�C�h���
���ޛn4
g����0�v+���Ƴe�Hg�����rL�}B����*z~����X�����y�~�.���BIm7�#���q\c|�^���E`�$�h��(�)�i�C���Ű�-�J�wm-�n���ּ�>˲��;T@r�t+ҡA%\�����S�v
�ɿJ�|m����h7P��\O_��K�j�kWr^�09!ا��Y|�υ����-[����bxB[��N���_F) �uZp��L������}�8�����?�?6W�'L V^�3�X2Q髫qEbJ0��S�g�����>��{�ޣ�Y(��Ԣ\��eOcx�5�
,R�y��3�οƊ�iA�#��
�jP;�c ��E培:Z�c�c�=F��U�ho��ރ�ˎ��%���i�ѝ%q�,�~�>ٴ��eQ�۰�$�|�W�%<�<ׯPo�i2=��ݞZ�m�)�^=~���,�Jb+�o�N����B�9��<2ۉx�J%͟nR�q��a��1@]?FpB�_�x0�l��@rL*>ml�zQ��@�b��6��'*m�Ú�$V	��?��|*��:��d	����@�ް�?z�v0� ���0�L��}Ǌ��p�������TY����#<I�zˬ��=t�:�� ���1��lL��-�Z�@��}s�H6�a��k4���S_}�_�>OH�6�N�tÛX8th���B�T,/G`�Z[1L'l!�՞<r�$���ֽ����^�#��a�R4`H�a�����1�CA�y�1�@ ڿ�l���z�u9�%K�e=��Y�0��y��#�h�f�pJ��ٺB�T(�Gg�Zǵ�DRK�;г���4*�V|8����H�X�`��J֙���)�1k�~��Kה�(E �x�+��E�W&@Y�q�@��T��SCzW�%f���s�ˋD�=�O���J2j�`�TG����%6�'ΗSg�Ȫ��V��+��,:��݂���>� 4{iEU�;W��#fT��~���񇜒j�Ʋq��ŀ�ؿ��'�av�(�n�������%r�v�+�ε����]*#(�L�/(W��T�J�]HW���U�i�Ү!V�Q����$��O�_�J'���R��b���c��MGF���;�|�4XU
�}�&��g�h�3��	��ER���a����C߈i��:5���}+�/�^~������Y�f[�����&X��[�x�ؤ�ժz&$|A��q9�Hm�G{��:R�6|����⁧�W�Q8ی'���i�/�w������nrzW�?#9 �\q�B�O�?��w�0��;�"��+��D_k�R� �h����F<�΍�-�Y���A*`�?J{
���4����x��d��/�i>�v=��O��g	�)�^��2l��16�Y��[�#R\�,�/����8o0Yȴ�E��7�d��R`16�i"<�3��T1z��\��ʸ��?��vv��j�Jؑun�g�8t���t_���9o7����
�2A�J#�A�G��Q�#x@��cT�ID3�D�*�[�.��ծV�ZY���e�����[��1�|<g�<�'�\�dEZ6�K�ˢ���� r�s�aZ����Z��ٚ@��'�����f=�>��}G�z�
hy�nS��{![�-{v|��`l���r�B�I�	����;�:]#�O�6�LI�ʣ�I,,**Y�7��+Uya�Y��Kjr<jr�@>�dK�yީ�̪�u((Pc��y�J^C��A����
fL�VϜy?��Lj�>��P�}:?o�����lS�ҕ׳t���Cπs�6�5�|p�F�[E���5�A%-�u�"��G�L
{�Q*՟*�w���j[��%��w�w���e�}3���=��&C����Q=�Yr�O�����c��j=���s ����o�7���cA�k�׽n�U�������E�JZ]�5��i<�T�wu/�z�PV���Y����3*V0-d��fY�o��j�h��~�yu�:��֘�|�?��_��Rb��%��n���
P�!#��ͺ��ω�_��iqB3|\�S}��C��Q�)�(.K�*^�J˯���@L���/���&��f㢼s'O'1?�d�*Ӏm�sC����cT�%� l�c�`�,��9��D�4�g���GE�8�>3�1���3[��C	b�T�B��1��y���ພY�C_��^_rѰ�]]�z�v����͐��)��ė���2J/Tg�0�����4b�]�u�ooQ�M���
b����D��*XK��������DGC;MC�'�Dz���`�B-o�՗1���k����sl�{�����
��Њ[8�Q(�M_:I"� R��om��p̋JQY�X �[V*�F���-�M+�9l3��A�������BJ�a?A�H"�%�:���<A%H�}�!�S��&��_�cF[M�VwЌn�����eP��!�h�ߊ��E2��������|0!�0�s�٭M;9�-�j����{��h��l����8�4�r��~)v��lzTDO�#��a	�^,��Iz�Z%�*�-�*w�i[q"�[��%Xc1wq��D;yJ�`\5`~b��A�FL�Z���U	P+�D	�?yR�8NCjy>QP]�敬���Y�����Ec��1���q� ����� �Ft��S�i$z��T���)�v�dT�w�hA�/��Mm�
Y�(����<,�_ͮ�C���.���<�o7�2��o&�^�$�=]�M^��co��C8WjF�&�����T�	�~��6�*,I ��K�l���)#���Jح�Gx�i�P"��en^0�9�%k6�G&�+��5�����h(�M��2>Y�%36��'u�D/M��Ό�C9Y�˻C�_��qw��L���;�E*[��<���3��L��5�{�~�S"^\/�kC�(����z��D��iK������7��b)0D (�"�(Lmԃ�k�Α.j|m�Z
e�Q�ި�	doU���a!�c�c�E�o�	X���\$��!�ۮJ�g������a΀�Gr�VCm䯺[�F�5�r&�m��C�WǵW�v��� ���<m�[G}��G@Ŭ���i�ࣧt|vL<�oh�~rb���� 6�;@�f[�	,��
S�p]�4S�2�mGƝ�C^C`��7�_4�Hg��;��0�����(��jo����n�C
��ʠ)s�_���)�y���P�r(��X�����gk�"WpM�����e+��hA ��(���¯T�(i��Y�����{Q3$�Q�Q[���+�j�ք�=�d����8�$9�D�حn-��o;WL��U��Xj��c�N�R��+��ː��!@&0����.�
��y��4�fa۲�bk�z���M� F�F��!^	��U��L<U�&x\70�P��H��2����9D��a��?OQ���5�6�{Q�}�/�u�	d�ߠO,TD-�M{Nf9��h�w���rs��Ʌ��<%�¤ھ�_��AR�X+�����`"�6wR�:�~�!��ϛ׋9Ip�&����W̲+�0"ڰnT�`�P��S��_�XK�Q��7J�����L�A����CB�ܗD�bO�⻺��=�U=^�ѳ)D��?��w���7��o��:�)�7�G[��c"e��u/b˙ �WȂ6�0��($��Ǻs�8���¶c&@elM(ky�ͧ���q�Yn('Y�����C���3�P�~	#��D�Ss $|�?�w\F��"�~,��3��� ������|M<���WM cV�����T��!�$��AчҧѠ�b�m3&x���e﯎�L��]�C��&��yI>��Ӗ	�yѥ7tbQ���u���F^rT���87����Nm*%���G.oO����������!g�lN��Q�m��S)�#��	�O�{Z��c�S[�*򒐫lz�8Tz����q-+!�:�B�\�M8�&!VH��?g�U$�	7���e�o���1��B���Su�{ଆ:���֣xs}��k���@
�2�ߖ��f����S��C����O�ƔOT�R�2��Uc�5�=��G5�o��r��_��wϞ�LW4�8��(T]A�3Iv��`h_��ٷ����eexaX%%��T�;�c �t+�Ӡ�t]�ȍ��5n�I�n�������6�6�_�5���2�,x�/5/D�N�;�T؜%1�����Ī�*,�g�&��k�Q��V������)!���i�(G.E�x����~w�|U��\"���YD�����ǟ�G�	�E<�ʮ6�mH���=P��H��`7�ʰY���1$*����:� �1@��O��?(��y��Ɛxj��lHA#R�Ax��n_����yH���Ƀ�XN�S����c5�oHc��ۅ�/��פ{�?�,�PO�ժOvz̔^��W,�t�0���Ӽ\�D�@~5��C?���ٶ��yKl��}0-���]�f%�
h�*�z�p4 �~�(WG���C����^d@>f'\��?�3��CE�:�ʖ���#�8�X��,-�԰y(��D��Oئ��v�(M(|�����!����4)��NW�#*��v\���/G��R��O#���n�FAM�@�y` �-4��8��Y�7($�W�YOM!�3˥h�^��?�Uj�s�!EQ]=� DR"<��A�� ��H��D1���E��'���?޼�A�'��5(T�ł�(�������t��irY-O�ryn���J�Ջ�uS)��JS@W^@S��lYh�L��g�,Ц�y���ﶈ�Gҋ��:��c����9GOWy%��vy��+���Ui����������SE>5Q�
[�C_L�?ۭwi�����!�g�p��In����+0 6���!�఻G3˻V�h}��阨D�l"�b��=[�S�g��tL�C��P)q3����� S�"y�8I�+�/.��2��jl	A)�e�m�|E2���݈][Z�`�Z>@%�5�{1�)�AQ�,V;��s�mx�;Kb�in�d�=F���?ਰ�vw��L]�O^�̝�|��1&����C��(�

s ����w<o�X�~�'Xu�No:Q���Ki�(�Ak`!z^�	ka�?�g����O���k�ʖ�B��̤Gߕ�ǋn�u������V*�~��;k�B���~�>p���a��Q��,��:}]�0J���ˬy���	��1�A�8����YS�Ļ;����<�FCB!�8�˩��T�({+tt3-H�$5=�A�ھ�P�Ap��_��j�d�d,���f�z���f�����Ն�DYH�S�=��ִ��_T4��~�&���r,�f�w�K�@C㮲/��(��o�,�P�r�CT�����:�/ʀ�S3u��zT[������'f���PB*p�~�A��� 3`�=����6Mx���$,���Lp�W�?�\�� ��Uچ,�dϐ��o�e~�U�P���?7��^����=�b�����0V��3�/����8��N���
ꟹƫ�>A���֢`��O$���Z?�U�DeXC�CO]�y��9����|7�fkd��-�v@g��i��>�ڪ�$Sc��f��7�1���I(�m:�{�����{��N����ȷ��-w�D/�i�!TK@��nC���������|T������Q�G����㈯�.:iM��/J;��$4"Qc麝����}��g8r��'���P�n1�<�|�؋��2���D3T]�|�>�'�;���$jqeT�(�o F���.�2z0K��[���c*�a��"�\,���+�-:�hj�YB��4��Q���!�����?e�$9..�x ��ND�v�=�WΓi
\|7
1�$%E;��O-g�"�̰��i�1��Ъw1"�s�Vj=�3�@w愿��z�G��W�@og�ǫHmd�(6Y)fKcQ�Fq�O�a{�+�dX��􋏔?�}��V b0��d<"�l������)����ܒ��o��d�#L��ƣ�y�*���d�Zb6d��@|��6YG[Uz�4b�@��p��e��!gG#�t?e?8h);�o[K-7��h3n����^ �h6�;gn�j��"�!�hQ��[\i�ѻ�؛fM���4V�%�uUA_����,��!$����Kٕ�N��|�k�ehn�	���A����٥���ED)��kmr���4���XF(Lі�=�AY����<�8����.'�@��$5C!๮M���|ȫ�����D5V�%
��3@)�ud�����b��@���Z���"N;	��2W�U+ƨ�������Tߗ_!���*��Š��u���"�[]�4|��#u0>5��:��2@�ج���@���"�ѫ��-������¥�l�T�"�����LT��&���q\���q�`h�HN�y
r6s���ϣYmͥ�x�oU��f��H�D���瑢�`a2\%?�f�B�"��X�~��&���O�[@���c����W���kj	���t>��]��Et��'-q(t���#΀#�q�ƴ�rdOw);W}o&���Q!�`�#NOd�x��UEWO���kt�=�Ň�,��b�,�	e����!�̂���=˦u�����.�:���l��[z�O���۠�� o�B!���86l�a.�L�P�����5<�1�|��A��d�����`	�ט�n��*Ȉ�u���N��5�l�(>"�>C�G��ӡh:��QF�ګ��#��T�3�3������ �b����:�5���a=�zY
E.�K�_$	 X���\���*
�%ƺ���|o�m6�%�	"��NBC��g:�v�� 8ٶj*��fQ���F�ƫ?n#�i�x�K�1����b��!X�|�h&	̭�Oz,TO�����(`V���eӄ��ЉY���D��+���VM�ai���<�K����㏉��q��̷)�6沜�O�������<��2[���b�O̓$/#(RS^��������YUB�v:�㕶����ks�
�&��;n�B���[���}�1U8��l��ö�����!-Z�>�%��)Q��57!k��3��J�~�v �Nt����T"���љ������L	�F-��7�Y�B.�A'�'g)���ں�9�t咳.>��b�{�ģw�ܺ �f�k�]�~��D��� "a@�+����FO����S+�XQ��ٶ�i<�_�E�PmB�\�SWD�OY�����GҨZ&��d�������
���Hy�y���jhP'*�>_*�ײqG�u�Y�Pt�v��=8�Hr����0�_}��j�f]rMX����s�~�Ia�9KAw�;��>�Ĉ�EG�ִ����G�U��1:�_f��O�v�ߩ��m$%�r����e�fA1���P��;G�J���݊TYd��ݣ���!+}��g��<����M��!���T��$Z&�p�r5�������,6���Q?u^��1OIlP�U>��$vUb��U�
9��d2X�vʣl�*�P�Od��'S:������I֓�V�m��c �KI��%5g�ҕ6+�-��g������<S>����٬���~r{m��|���b��d�ʠ��p��~Rt��1͋.]����?��O=���г�X�ʄB(��z��cތ�X?��8xWT����߱��c�d��o�~q����}* �	Վ1��ہ����)����[O~|2���C����^�v�zVO}i�XQ���t���lb���J*�f)�
�qK�tt,��]�6p�bM.��کl�w�q��^�,{�$\� �3[Ҍ�#̷����h�E��47Ge3_ƇA�kԄ��v~ʍ�C�Ź�%�Z9pW�Rpn���:F��|0�]�g(��k+�)[6)��OL�7;�tH����M� Y�c3��p�p��5ֲ�.�P�5ڕ�5<�Zݍ5d9��2��s��;�pC6}���3���j"�sVɗ��m\UD�;{�,�>���#���6��a>o!�Y�Y<6^�F_#N�?�YD�g��E�p�;f_5q��ъ�]m�}����OS���*���G����u٫�񆛳�]2��+0�-��8���[�e>�A�ig�<�y�& ���.���j��"y+�>7�Q���R3�,*����.^s�Q6}�{�%�`r��n�����]3�H9B?�Y��AP��a�<C�r��s8+{Kwgl߈)��;m:��^^�ՠ�-�S�������?�H��gQ"�ͥk�c;�V�A��0�g�v�..>���D�h_`r|72��;,��h�����g���2'q�`-5?���N/ �a�4f�tL+��y5o?���gDަ�-���~�,4�Y�X���%��28�4����u~v�P�Ǳ�/�D�4F�)3$�@�zx�#�׺S4i�d�$Dı�)1ԙ��6i����Gu�Q�z%�rOMj�'I�M�����=��&�ћ��Kg@�s,M����>Yz�J�k|VX*J�����nC5�uHP��'�vZO������y�,�ޑ��Ƞ1��Xɶt� �r%(1����LeHs����i���W4�DO>ٺ<�"D0썭�g:�[����W.���l����D_Jf���ASQc0l���8E�y����ώ+@�Jד)��٫l��-�y�S=���8�ng����I��J�N� m����Y��c;0J��n���4Cpꛑ�D�G�Dū���ܓ�V?�mcfs�3:I6���[JG���uU�ĭa�5ջ&�)���o�Xb��X���\�{~�pI ��eԠ�28K�S�����[j;�,R����X�=H��	�U���~���MW��՘���繄��n��c�H����ڡA{+�a�TVjǖv�68$��p�W˱�=�
I(�<�� �l���BC�>XqOm�M�A-���p��������x��J�Gq�~�0��vS7���e�ֻ"&�E���Ʊ~`pTH?�������s�&!��Na��~���0'~J�ӎc{|@}t'��mkT��1:��V�}��[�q�T���7��p,�UC�2p/�-H���'=��Y�S@>\B�,�����3	�*Y=����������⣾X��'<Jr�ͨm^^�K|��h����	X��=�����#�ò!��V�h���&v��h�n3��j>�@�z"�7n�_�!�G�!�a	�!�C^2� -$1����6���F����XM��EpF8�qo cY_x�#6HG;K����7/2����������v��/�u��x�?��/��do�;
, ��K8w�)w����r1��<GS?����U�X)�����f�Ƶ ��y"�A:v
�nh`&Rj�Ϻ����_K]x�"�\ڰ����K�/�T���~����tH��!�5�&����M�@���+v�@u�Rǵ�*��}f�?��LS����@z���8�ˑ�h:s
���}�wul�T������+*�,N�n;�T��������y�5O�����󟒹.��K|u\�&�F�~t�����ss��r��g�����w�����n��p����cŔÊV,H�f����5Q�э��Ѫ2Shs9��R9���ř�2/������7sA�y�֥<�z(~�!��KM= ��m�ZGH��Zp��.f��K�Qq�(L~����W�"�v��z��~�[�2��L���T9����Z��2���o��1�'�х���g
ή�ȩ8[��� ���X+��"�g�`�	rQ���?D��w�b!����� �/"E�m:��{
��ɵ#u���u����"�����^��}aui�ʹ�HHՠ~��:tJ��+���a$����#�ũ�o��+�L>Sz���%#�Ua��"I���SZ�����m�ћ��6�M�`'W�*V�ϛ��N2Z2x���l|6"�8�Rwj�mms�;�8ոC�ŧ�:�6��D�L!!���K�ե��O_eL&�r?E�G@vz��*k>1e��Κ����v�Uc�RB�����Ě���]������W}?^J*´\�h�0` Z��e���TM9s�}������ƙ�p�!�|�]����aed��!H��, ;�[������R}�e���-�>��&�q�݌���o`U�)0m�x�%^�>���,�
�(sȼs���;�Jq�Q��#8YJϜW�y�)��A��?؋A�0i����C�e�w�t���~˞�|�UY����c���)�k�������G�:��B�Z�ƍ���O@�y�w�T6�ֹW�zWx�x��j]y<?������2������5 ]˟\+s�D0��|'uz�f!�;ϻ�C:��k�؅9x'��Q��tP�m}'oE-��U����,��a!c�'�����#�����;�Ur���%�#���F}�mV�Nɔ嚱�ʔ�xh,�\�[�Dl�-�<E2�N�}�����(Ha&vnq�J�S6�2�����1��������|�v���ȳ3f��'#7�F`��nD*5���ڌFzU��	ԓ�N2�_?���,t]�I���-Rri���ń��-������8y�؃Vϒ_Z�a�bd�����i�y�K��\;�a�4L���?�~�C1�����E�2�P¦��� l���8�ɛ�o�&м�c���u5+|����FVc�|f�g2'��"9քu�)>�DE��f�gC�9�tD��v6��&?s���^�k�f�ˋGaPBl�k)]���z
#�Y�V����g1)�RL��C�$���C2tv��0���{���h�࣡��k:~[�ǡ��h����7�D���֋1����O����CN����x����d���hZ��)�peYڪ��h�r�e����TVs���yGӜNp�w}ls�2xW5Q��>�g�d�������ʠ��� �n\4܋��~��r�=��f� �0��	�P�����͞����w�摡��?�����1���n'Tϭ����>�rC8�m��;� ���O���]%pD��
��^?���[wJ��`�b]lP���uz�X��Mx���������i��2}�S�p�dQC���6��RLk:�T�!�+%c��5گF�9޳��9���k�o*��^���
���m��&E���ɸ���	��S�wS��qp�^l�=�tO�f�6�0�nP��Z���ɑc[bT�y�x����,)���5�����9YP.�=YƐ�Q�o�}ˊ�v�4�I��b�����o���
�`�(�[t�C�������/"�)�[�>�֬k��B�,�Dש�"m]fʪ]G��˃��\a� ���s��3�B�P-��L��0���l:�~�(a��L3���()̽�Dk����Ԛ�9z�/k��a̓��X�o����fL��� �B�t��X�++n� ְ�S��L�P�k^��Z�x���$����Ǘb��Rc3F3%/rr�	b�h��x�K
�.:��������)�hH@�*�6�|$<}��+�DO�� f����a��P�`�����3�0���Q�{��a�[y�eJ�/u!����i����!�dh���,ʳ���^��|��݀uj��!$�̓���@{���	d� i�y�g��R�{-N��J{%��f�+�:��8�3DYsadJ.D��z��<�D���@�p��v|%h�Δ�m�J#�C�Ms�y�
@��X�"͕^�iSD��amv�E/�/��!���v%hē8LL�=���Lkͺ�"�����L3d@�ʯ/�nR��x{:<�>IK�K�������� րB��C	��e?nčSEP�9m}��]���2n�L���W�����7���H��̮�����ea���[��E�T�t�qv����M����{��Aꡔ����"5�3��4?�qk��[�䘰ۻ�s��t�ᔳ�,��񱐔�3>V>�z;K�!���4��  ٨l�3m�.��
mO��t��qH�)�b4o�_�w�8AoWi��tʭ�7Do|]%A���^{;k���.[���Xv
/��H�����߇�c�:���#q�+4R��p��@���E(9v��Ŕ��yג��~lx���nr7++��r��^��7��R�Wa�Pݷ>�ǚi��Ү	 ���(���%�f�յ�%F`�������VK�9R'Y�ȬO�� �ؿ�7����=� ��;��K��Ķ2Ӻ͖/�#[�e,��,�gDH+E��������V��Z捁_��5+�Q�ll���S��PD����D�TX����ξ�vJ����l�R{��[+F	|��N}<+�S��uB������{�c��a���g�Dz�kW�}�O/t�bw�'n��(Yj����t2B��G}@-��I�zqG���"��'%&��������y��s!�T�R��1�a�pGY(����d1
hB"f�B����k�9&���$�U8Vsl?�6��}1H҅K��
=�q�
:�d��wE5���a���qRSqnq���W_od��~�%�f�׿�����=U�e�jF&�[��Vk��zD���kO��b�zu琻Ġ�6xD4Rsʢ]�
�H�q�SHm�Q;�8-�G�E(~��_�����P��^n����iof�f~"�E��͕G�A�F�u���<ݜ��NK4z�H魥:kя_*o�;CP����m��G7����;3������Nz�ta�<��<E?�@�m}��,��jl*�^wd����n=�8��C +mvG�ó�~.jk��W�F8N���J�|����8�~t�S��m�<�!9��4�K_����#��o�.8j��c��	����h���H���v����*��Z`�s��д����?"m�iǸw�>Hsn'�f�N�8_���?�N/I��0��!��z�x��#�b:��tp~ؓ��=npCs0���v\���"9ZuRS��s� Jj���l����vO)�Y�'����!�m@��/�:��p� gb7W�+9P��G��&Rm[��$S�(U3/�7)�������FAn�E��T?-eĺ^ ����u���}8�n0]P�px�2�#ė���W9١�qm�1{�l�<�yV<X���N�,X������v�~������CK'.�O[
0�rW{o��(c"��~��6/3^���g�����Z��cY�8���[�ДU��xA�y"��O�j�u��� v���C��Q,��-��f��"�j��hJ�����P2�~��
g
HI����(v;��,��߻�w��#g�:U�90r�J�}�<��t��V�Dȟ��|�KE��Xԑ����r@-���х��I��}���j�$ �#&�ǰf(s(�_4hź�i����K�#���T�L��R[!�r@j����]�"�h԰;��S86���>uҩ!����1��Ŕ?�_i��@��$v�����&��w?'�ȝ�X�	�G&��ꏉ����̙e�6O�	�^�p��G�ό��������%^O�'GPO6Q�q�+겔�P��Sm��Z�.�wp����h��"�<
�[t��c�"�����Q�*@Ӕ��O�m�{z�i��}�O��z5���Y�t��y�f�v~����-�Ͱ�K�˓*[SZ�G�DC���}������ޞ`^��"����%�CC�+ɪ���3��* ���r�&*y����)h@�M���aXOg>���
|t0�`�_-/�&a�TQ�E����b�c�җ�g9nW�(+T��]_�]�"{����S��D���/z�g�o6b)ûII/�Z�uf��;��M�i��;p�D����M#s��^Kߖ�c<�<p��p�,�!A_ƏT�*���m62������	�b�Jǰ�����U+�9B�Vb�NP���o�ʌf|́�&��g��7 V��>������ś�5��!�[���*D�Ƌy�͋��ۥ���Ihu��Nc+�<�$��^e��%6��G���0�Ą��5��~mt�0���2-��я؊:������|�7-�\���l4z�<�������Ft��ܠ+՞L�kU�| &��a
W1�۟��� ��;�~)J�&�5O�8�*2����ɔf��u����jdl&�(5�ʊ-� Fg���h�x��@UO��u�T�5t���7M4g��n��x��]��	M�4ۭ&"g�0|T/_�_N�O��j��$oX{+ �Ưm���i8R�E[.�����v�G�B?Jw�<ʋ3$�T�ޚ���H�u#�YLL�S�n�JDߨbS[�YLzdt.�o"Z�}�֕;h�k45��TI8�A�Q�������88Gdr�g��Y��S��:���\~�~��qET{X߀4�x'�~��`�8��Q�/�u�;vKb88c{Z� *W7tو�N�J��^�;��fajl�5��W�<uk~�s�#|������Ra�Zꫂ9V|#N8J҈�.�`!!�L6{�i�H��.�x�p��?�Y�K	�r]�-ފ.b`P��z����^��8vm�2@��W�_Y ?fL�w�p�E� ��؛�/
����^y*�#-2����Ͻ���F�m7M��L��AeZ4���Q��$m҉�^$�:��Y���D�c��,\z����G7��V�2R<@H]��n���%}X��O��� ���d�lX�;�]�؄�P�o$���K���*:f�sS�P.f�X1�����Fe���R�@\�#¥~���w	a�	>�a��A�`��-�33Ϸy��Պ�ը�j�u����4{���L����V a��A���|���a?�ĕP�K��ܙ}ŭE�[l$Nkq/Xw;fG8q!}�.[♿�Z�n�S;-�H��/���)������#.(KJp\�͡�|�XC���D�dK���5��Xa�b���|��`Kԕ>bm�6�}x����ە�)`-Ļ'*�_�fr�K��duR4�<S�����%������<5��6u$��wlCљ/���Hq2]�k�$���#��M=O����Ϯ��|\��NvN�C$�:1G�����J1��Ũ7zܧ��j�n���ub�Q$�����4ͽ#G������:�p�@3Bj�zYZO�\/�	�eG]Y��]��K�j@7���8��zo�8ͮ`U;��K�7�zSQ���"}�����&��N���}���V�*-'lR�x֭�qJ��g�o֗�6�Nu{r̜W��67�Q;��w}�/p��D�8&��e+o\�Ef�u�K����2��6��l���~��ߒx�[)O��ob���nVU�\ �DC��G�z�_ �KP�إ_�;Ho~���`��t�a��n�v���'ׄ'��x�G;�ۢ��{E����_���]��uՂ��\qݐ?~𜅉��M��!}:5����h1�:��J`�̬L��_�UkW��V5�#�S��q�d.���\��N��i�����T�BF�tt���0�3ŪYq�R�X<�U
���آ�O�X�Q��}�2�[rS�l�tq?�G��I����]t���B�����p4s<08��U}�zT�z���y�n�����FM+?Ӣ^�'��D�c�e<B@�B��fEQ�t^��a�H��Fuӎ<"�e�
"F�f#T���VM��]�΁l�"�=�vZr�G�����O�a�۔ �a�D�i�vz�Z����������ʣ����ɢS�#4�ȃA�i�B������tI����s�=,����\�M�����=P�J�QC:��Z
���Oԟ��e�b>���њ�$���+��g�. !�%���޳��e��:m+�o��{�=���_��-���wG�7�����R�/"v�����+D|�|��x����P��#z�FaA�Q���ͮ0Y
[�2���5���A�n$�D����X3JxK��mRU��0
�a�&��ە'���)��g+5���G���IS����PŜc��(�B�y	}^�"%�VۆV�_�=VV�?U�����Ί"!�Dd$��T���T:�]��������5y�R��1r,}s��t٪��},�A�����Aǐ�W��B�.�M��ԫ��ӫ~���ȷ?1�GD	m��xU/6e	���X��pd��Ԩfj�j�W�&�Bt��0�<�_���\�Y�Y���Ys/Q)N�q�~iHU�� )?�0:p*��\���he-�-d��&�;yP�������?�8JBC����\8��!�uVw�h������9��!��w6>��-��������O���%����	��2`�&U�1�F��(SE�YϹ^����hC��}���u�����l�}�>P��H^�Ƹ^W7�4X��rX�U'��� >8;�o�;����3IF-�v�G� h4�Jq�+�oc��]Fu���e�3��J%�ȮO?��p�9��G'�)��!�����mP�����>g�ˬ~nqi�儀1:��/d���ϛ�:e�a�Vi�2��T}��Ƀ����0���<�ս]��%��<�O�/S�1-FaO��a�ᐂ�6����\�W#tQ��}��E�e���d=Lf��Z6R	>�k�m�:uM�yМ����JMq��]Y����7��e��?�O-�jҲ����f1���N�!�E�$e%�z$��֙Y`qp�r��v�
�����6*w�m�����6��7A��}��i+hQh�x���"��\+B��'ކY��<>f<(Z��豼�5��`iE�z�RaW$�f�a�<���3�j|�:
��o�aM��gi���t(��1L:��|���%��]E
Oߛ\F�Z��N�.ܴ�:�@�d6��d��p$�p6�8���윙�u~�J�<�C�FnE��BM�7Y�6�b��6g��ax���.�����E��Y_�*�M� ���%�76>���E׺�'�P��w�Z��7Jn�ϔ%� ��ٵd�?�~�<�p>���yL"=��nD�O�YCUj������ ���O ��GX��q���� ���n�G��W��=]��.�5	Oj{�!��lr�Y��;�&7�*��K:��8^���j4�p=�\g�.�������}Ж�r�g�3ON�xl|�W��;�A`*FuU*������1_J�����UX�To���h��#
�@2͇�����f'wű-�t~z�
���<��o�Ӟsê:CsN{��d����=��.��]�YW0բu�T�ʡMY��]�WKg�>������K�5(�u���O�{F�E�&�8@����	�Xk&^�R�'��O=�#PG�&Ni�@��"Ƙvz� �"
��P��x��,_gl'B�f�Λ�u:��M&�>����[)v�r��}���~A*����n;��92��L��hY�uz�Qr��7����9���'�5�%��f�J��P�����Z�$�lLI�p٢�7�ɋ�h}�"���c���ވ��ܲ<l�DiV�à��(�m.�2�mPG�t�[�/��1/��m����*`��Ėߜ�g��AG zD�h�}T�V�&����QV�@�|e3��,�$�Ŗ�N>� ��D��b����v���V�vX��ԩH.I����{:��(J������ɂj������`�bی�n����[ۧ���+c@mɆW��͒3�H�zt�F���.��dY�a�5t| �3q��cN�Q�I	1i���}��m�������7vcK�9����AE�]��qD Jy�7�P����VF0�� )R5=1�E�fm�OoxPh�d)���%���UUl�NPE��1�?!���������?�b����UB��YD��[!�7�R�uQ��mR�f��uĉWqb�C�O��pu(�y�{c*�AQ�ݩ͢�_��q�q��I8A�s�{��4��u:|����}�ä�^�1a�t���A9ׅM��,v[%�3��cI�(���3=�s�u.]:��%�
))K�_�u^�9�ؕ��Q�'|4PN��}$��B�5�P�������	�Q"d>-Ti�0��aσ ���r�*�n����ab_�HC,e�bX|�x����&�����mi���1�	��j�ո
��c��D�� ��9�#4#�'����@M�o�Cg�����!blW[;V�Ҽ:m4����<]4󒖢f<��V1W+��`X �w���f��=�N��k?ޏ��t/J7��~�"����ȡ0Q����z��F,fh�ms#���ܖ�8!�����,Cz���á棚E��ݣ5S�&����Y��9M([ݺ��BX^�	�2��C9@�K�$�FZ�t���u1�XY��8�A4)��#0�1��Լb>���3]K��%8��,5hz'�g,�/�呼 ��e�p&��#I|~VMj�1ƉJJB�0qRt<�=�2`���{�M��):qی��+�f�?!$��"A6�d�3iթ[d��9��N�Zx]��u�Cb�����4�Z�'�[���a �VHf�m���0�����������f,����������|������g6��8�F�歡��{{�F7��O�(�+$�Z{�֮[��	wt[A��G��q 1#2�i��JA�,��N������W��/�#�李a����s�$M0t[T�}�x���M]~�c�<����/�%̘3T��r٫;��9~+ns�_O�����%�k���|��s����z��eMI�8L�$'M���.�6Y����_l�	)�����説ܮ��m���%�ٵe�F�h�:�C-��?�l_lH��l�#O�ϵ��iݛ46��0�mH�� Y-=,ө$�
��K^�ŰUE#��!�I�z��6k��)^���`1��=��p�߇
d�ә3"����̟�[T��c-�|c��`�]�C�G����v��i��TGM�K{�N�_o{��b�� [�~T��ߤ�N�G��O)��f���}�g�ٿ���t��"�K�մ�]	^�}���έ��6�G*���C�\C��v�D���ڍ���=g:��R\$Ϙ(���'��cK�:![�)���3����ߧ�N�7b��I�/�K�Sh��5� �u�c�#���Ҝ��o��#����L��wL59��׻;i����9�H
(D��'�B0�����4��0����cE�R�j��f%�ˋ5sAp�z��SZ�HL�)F�-ͪ��ޯ��C`VǘɌD���!)8g���O�OZ�lȓ��o��8�Xx�,��E{NռC,�����7����Kq�������Aq�vɵO����)s�v�xG�i�Vfm�|�B��LJ(U�5�Z��:��X�z��G��RN��>��F�s��J��Z�����k����(k5;�QL]��DY[AdS��m��k�'�"��k�ڌ�\q�g�rn�#$p��6�������[8^|9;h2_��Q�ߪ�I��f(QD��kb,gVc�I��,y�U��Xj�,|���Z:k~^�!k�}�pr�
��Cq�����R&�{�%��q���ZUR�lM`�q�L��S�&����|J��A���J���h��\av�v�$Oܽ��RjF�p*���5g"w"*ؼZ��t����煟�7V�x�����?�t��)�Iy-h�Y�|�@!�t��:�p�WJ���Q�|̨K�luMR�2���g�C6�ӹvË��;���G&�ʟe�P?���Nۗo����������"�"XW ��C��jL	*U�M}KjZsG6�6�@l�X��+�M��6o�vH[�wߊ,�R72�\98�-��+��c�4�q�]V����6Hv*B1y�f��u�̗�x�<#X��\"� L�NF�:��3�@W����{Q7_1V߉��'~��{�����me3�u)r8�&o��2�=��{�F��Kz8��b"�8)2�Qd6-��c"ĭ�H�{����6Pvݩ?�L�s®9�ZFB㑜��Éz���s��N�|9��g1؇��F����&�D$^���/�|ҺD��_�l�esL�U�f|~$����c ^���y��~g{�ex#�7��=���|��A��x9�pոI�<�,mS�-!cr��CHL������9-JG:����J*-�R#�=k3嘛���A���������V ��V6gp��Ԝ!�w6��t0���͙/7��]�?�J��FX��dj-�v))��@�K��|�q�[9Y/~�$x3>�Q��m�7�~�-�/�N��v����
K�Ep���L�	痒�t�/�R�	l^^�k�ś�|h�f*�������������!��"�������S�4Z���z�T���"^T�	9������� f�A�7��9R��1�{c�;!�Fc��a���O#��V�꽥�'�yp6�6����׀jq��[o0��*��ՙ\�G���+�d��Kb�[�K[y�f��CKw�F��BX����o!l;�|T����O<vr�&Qii9g�\��_����A>�W���aPwuح����U��?��LyO����(���6D�?�7/+%�`*+y��x��_� ��bճӘ�Z-��v
�����T��j��{sJE�m�=DٺbpA;��.��G�gI�i�5D����r�ϒojvP�����ZF�t��UeF��2�jFK��G��"��0����x�j =�D!��X姟�p��q#(,�.o�r�e������Z?��0�4��(G��;Ȥ�p<s:�t���rfɹ�	OM��=Rp֒V�:�f�L�EXf�:]��4��a8C��>J�ީ����r�%�s�r*ޑW�!� �6O�qfHa��D�=}F�o�yꜶu�~l��i����l���r�qX
#��G*�l+��U7�O���#2��2{܃�T��1�):��+��8�4�z�r��.���*�z�!I�n��<�<�^B�Bq09�Ph��Q�=sd�v���[���Ʀ��LtMU4u,ێ}բ)?v�rќ�
%+4���-�LA;�a�<��a��J�l�~J@���\��U�>h��a���W��p�F����F��e7��z�&aO�l,c?r�!#�0m���!�������-:��=���9�k���O��
���֦@.���8�K.�N�/��g��+#`��y/=�h�6,��6��T����Wx�fL��B���-�}�w��jP�������o 8��v@�����d� u
$���>��!�T����:��sSڠ�f�1��w,[ɒ�EŌ���_o�c�{��E�!m��I��8@�C*��gi2�t���'��|�3�.�|�HM�u#\��Aǔ�?/��0�� �.h��0lz��6
j;�Ԥa�h��d��riz|!~�G�k�Y�j���V�*�ew�B�ފ4�-7�>�y	��V�7WK(��0�6%�9N<X�n���w
�b�<~��hm՛Nd�B	�-0��ϓΑ�)����SD�c1NY�o2*RZ��^rf}I��P�fM������^d2V�����[����Ο�{G�� v|����w�bkH�XNT �b`4���!q��-'C���cgT0���B��lߏݸn�X�T�](��i�O
��Ÿ��59���V(q��09��I�S���l"�<a?�AX���"`B�h�ДU������/��	^gr1<�Z��ZC�0���]E����M�0�]�x��I�:��Άev�������;����P7����i�<c�)WӼ|��f�
�m��*`�"��*���,3#�,G�=nU�{VN��a;��wCW�Z\�6;�b��#_�����%��v2����.YUh{1�*&$W�����O��k����*QǢG3�MV��[���T
�j�]AB����,���j����l}�=^���-A%��<t�-��Hx���P�敇�h�ׯ�ᚐ�$��3��G]�5�+��W�\ �߮@s����S�V�m���-�X#����;��Oc`���#����+.�Ӗq4��f�EF� �v2��\ɑꞠ<�6Uvy"�K_�κ�C����|�x�ąA�c�RJ���+�O9��l"�e$O1e��͌�䌏yt^�c,�U|�v���C�����rft/|d�8����m*|^�ެ�q��
�.��<N����ߝ��&~��D	�S��_�"MI}ӣ����H�ٞm4����@o��"��$�oF/�	���;�� �=�~�W�聡A�v��)	c�i~��B �D{}�4�llc��Z���!��X�ܙ@�wo������6Jj0��$}@^IG��A�瓍˱���s3fa�*������쒪K���akW4�+��ٹ0�8�ZB 	�ո o��Q���e�ӌ/�k{`�]N�[J�Դ(���1g��'[ڷs`2�$�&����Ph�#d���G�WWdP�$B��1��Xد��1��w�Ź
�����S�P�3;�݅ t���(ʷ
�W&
Vw����%���F;.?�9K�V&�в��B��m�c1�Y������V���7}7\�TYb�$nrT��HJ�W	�C��фn~k�]�I!�ř��#M�tE�@�2��i�i`��;$�t�<�S��tbe�l05�ѽ�2���	�Kg8iDV^U<��U"�<JB	����%�3�+bOK�Ze����fd{6}M���79>Wb��9/xf���uBjs��˻�丆�/*�WYng�RmG�]y�Ba�u�	��P���N�B��L���b��N�=�R����������'���[6��]ӿ�i�:'�Qs���ր��;ۛb�u�.C������@��礋�1���?�6���
52����W��H��gs0<(�䘦��KfZWʅ��e��4��e��wM�Rh���n���`'F
Mӓ� Pj������
��@���z��A�7��w��V�qNl�� �zl���B�-%{a�d��	���*ǧɜ��-:��\.�dM2D��00��Y�K��ֻ�Kt�:0&��V��N��K��R��<&@h,
�k5�]� �1m�Y�b.�v~�_�/"���4/U��ŷN���E���>��BQ��l�47FUV04�)�9*�M�@�����F�����3��Ǩ�Ii�Z�c.IǺ]�{�H.��յ>����ߠ��k���ܙ�rBkنI�C�e[�����P���h�rN���:/�Ty���f'��GU~�I���ֶG�O�*￪�P��l��$�f�5�b�T\����ح �1�咧�&��m��oj>d�1[M�"��U���2R�I��V0���GYO��wr1p6?9V��4)6�V0ׁ�����7Z�g6�W��.k�RZ�L�nc���/���7j@Y�k����M���,�w��8�GW�#JV}M��n��0�m�c)�������n>�U1P�ZFu~ժ?,25� 7���H-̍���)8뒾F�ʉ\.w:�L"FAו�l�,)����s���m�?_�q;v��dl<�D�oCx5!�M�ȨâV�P7�9����i���w��QE���dPK�D�!��E@�E�*��^�`)��	b4rʻ/��3N�ѩ�q��"�G�ePYh/�޺�΁�9R��z���<?�u�%��'Uc!��P�s��5�S�3s߫�携H0E8:��� ;�+0T*NN`_�+ѯÀ��U2��ʲ �R�Z84Gi����w����pcߞ[�Љc�.N�*7�(14��?H�@h�9�V�R->I�?l,��2�{�-��1M�ۯ�<U�,�X!Q1����@ o��I�b�ai�j�P-JԀ�Crc�Czke"�f��BK�yq]�lb�k�r��G�)�dL���Պ9���x8`yP�l����ɠ��v�R��N���R|�b�1�_�����\������#SK���ʭ}zi��Z�����|�(Q'Lv)Jm���+|d���uZĖ9 �Ǘ0� �H~[���B��ǿ�$��Lp�so�k	�֑X�:��
J+�~�j�͟}�࠯-���1�x�d��;�����7�fΪ"Ҫ��iGTƙhpѿY��ec��
YC�-<܊�X��I�bq����ݩ���w��[�{Z �δٌ=�e�Q!o�Ia�C���F,.�C[��Y]��L�|I\\�.���Y��:���rٳnK�(W��0���\9lN��X���c��#�����p�KR��w|��0����f��<V!3j��:��M�c|��������˥��� d����8�e](���p����[6DZg�H�km�N���k�^iޕtީ!���-L����h�X}�΢r(GI�֖3p
5�!�O�ǌB���"�G���l[��>�ѵ*�8H���Z���u����N��M}�Z0�P�cJ@��w��Q/��\�h;���w���K-H �@Y�^�΍@p'ȼn���J8`��BV�<e� d4��] �,���������8�q�B�I�]TRgňv����P����,j�<�գ�#�*�������7&?|�k3�������J�B����&U�Y��w*��G�\��ַ�Ca�O�]�)��E�7t�Ԙ�?|�j�J-��<��!זxͬT�"^�d�m����G���Ѐ��<��v�I?���P�T��Po$��α���~���T&�mJ�q�}�dH�=�֦��t10Km*����k�E�S��g���E�/�� `q$�Lre캂����t����k��� 7���,�=sH��Eݤ�Sv�ֽ����\������-i^��-�����j%�U%�Y^~�٩7�^:��lW4P�C�������@�X�G�9�Vm(7��d���K�6���h-��K����_u�k�9���A�595X�a�v�&"�l�}`8�c�����F$S??A�Q5�ス(e����5��4/��rS��H�Y�6񚦿��	��*O1,��q���=���P��g(ƨ�c��D)��S� X>���6{���˙���.σ� �zHg�"݌(����:��r�S�ơ~s3�a�8�]��� ���9�WzxtcD���K��Y�{�KvE5���5�⼁�7��9�ga���+��n�a�qқ�&��ի����*�)��L�^{��D�l�h �1�).�7����W�m\�?��O���e >�pݢ�񖍣�*&�����,����� �3g_�/�]a ��E�����¤fj�H.ZDP��Pg����M�D�?���h�F�Y�si~ai��G�cHy)	�V 9{�?� Yx/�{,��"k�_�'�hi��a4ι�[
�6��^�bWGY��S?c��J�)�}3�PEz����Yw4E�Տ�Ȓ�v�K�;s�LͤڠHLue�{7�j]���Z��=����?�Y�=�-v��O�o�IR��ߨ��+��/h��G�ܺ�Ȇ��N��*�	�?�%�����۫[�F�����t�&�̬�3^�@�]dZp:5??��S��~���Zf��=<��u'Ҭ��_�;��U�|��~����� 1Zi�2B��y��`�HA�=M�%,mS�*��E̐JF����`щ5��3�LM[7�^y 0㙻�7���ɉ��~'Rبǖ�jෳ
�+�|�Ox��I�w^� �~�Y}�e%�+y
��_x�z��X&�f��,a�X����ҿM��}Cb�rڿn��ANp�Lpj��ً�r�Y��]��~���4�^�6�p��3d?�H����T�t�m<�t�0��-��C�bܲz�b�tdΕڙ�-J���˦����!)u����FlԐc�]v�x� �J�%��R��%P.�%�J�7y�t�baJ���=.C�<Ϩ���W%���rظ�Wn�)��$�7�'��܎�������㉺z�@Ď/zP�u2rk�%��-q#6�tda��7Y�{���6`WՔ�r��8�D��D)x�������mR�\*Q}(�~Xh���P�����5���I7	�����!�8<�l���O�B��(�̳o�
W�<ZWZ����0w��s�=�]f.AA�m+]�K�l�7C���uRB�/��\w����flcqSp�,�Exe=�:�pd�w����7|y���S|��T�#\4]�p���n���l���ҙK���?��&Uf�LO��:a7a��l��.Ǆ��'H$�8�^��6�M�d3��A�ab	5f���k$B���/�8���� _���a3�s�ON$� 'J�.A�B���5)����N�y9��n۲�y(ē��ba(U�DvĘ��0����x��T����;��~F������)^�E�C��]cܡJ�lR��=��{l&���qIhv�Y�2^�M,X&`$)�>��/;<�����8m�f�zo>m0�K���c�l���?~�Pk���$%h�A���c�����Vt���>TUݲAN�@�0�ܓ�ꢞ�ۻƦ�W�5�H�(�T$�	=�Xu� �F����d3�D$ ��y��T�גW9�����m�p�%!�ꋔ���������������	���������G�(z.��:�����L�BIP_��z�čo-�:kM�R��X�X�089� �07R82���4��_t��x��v+�4ʼ���G��FS�*9�%�3;]�^�E�[�G�3i<�>鐾�Ƿ����1+gn���3u�Z0�#���Cp5tn,g��PQх�rr����1L��ϕ0o;]h5���;�0t�74�BӃ����� 5}Ĭ~)���2X�0ĝ>A�_����4g��Yɾ{�;����ߝ�Q�e�A6���QB���B9FL�1>���A��9��8T�h��g��c3ł��$��R�����EG�S%zvt"����x�͓������<Rq'�G�$��P����u��y�f�<+c�ж^ʥ�� ����������+������m�N�g�B��,w2���lM�!�rȪG����e4�C���˻��v�#���yx7Z���n5%@�Ch�ZI}Z�٘��k��4��38�9d5��8�F>(����'T�u��Ԉ,����Ԑ�B�S��-[3$�W�@0{��$��U��C�G�%+C�c�T�y���������M[�yR�*<<���!Q��fD��9LL��
���� ���O��?���7�1 GJ�@GN�JJ�R��&��i�_0�n�f,N8�*d{�w�` *bD�9���B~g¼���0O S�<揜��5��+�D����/��x��'>x���7�s'c5�͊�����F�/�zrt!5�&�$>R�a�H�_��	��
�/v���ߠ|�� <Ǥ��v���еf��Z��!)$��	#W!O��R>���ٝ�@,5KKV��?^Io&��y���#�l ީ�v*�}fK���ЋuY�$�'��C�1��0/�>��B��2����
�`܈�=y�	Z� jF2�Nm����sZlZ�}L�d ��� ��~E♬qz����Mt�~r�?uc�e�y�'����J��p�3ۯ>� b��,v5k@��ah�{"l|M�%��0^��k�$FG$ ���8o� �E}Һ	����t��퓐���:2+X��E���X�[��P��bH�}H,�u��#�vuz��!/���w�ar<̦;\�.a�j��to����pP�	����Z��-xh N,�6P�R���Z�G��'kNsL�k,�v�W�y�����ϳ��3�r��Ҹ�H����o�1��F�>~�%l��'#��n����Xc���^ON������s-(����o0ߗ_"�#!�C�!I˘�g޾@^ng'm�7�8K����Rr��4�6M�+�������6�V���$����Q3H�۳����~�9�Y��g&��q�;}X�2����uZ�0����ű��P���É�aYVņ链��T����-M��̉�c�*��ŰpΨAzc�*���8J�8X<4�2��iH2�TW1f��K�82��LOc����ݘ���<vJ��C=�d3b���{̲�Dd$��?�G�A��Z��������rE����ѕ��`ZP'����W��JZ4^���?�7Y.�D���!�\$Z���9����sӾx� fv�+t�L�d;i2u$�zu��Q=��'�Ȁ{��ߒ�N�1�9(��EyV	�E�mw�d�{��_�#�)�cv)NO�$�Hdu
0	����4�>�����
O�n��q���=zE�nWg�^�DJ��mל���2��Fo*k�Y��i��C���8⸬��3Q���Rǻ22W,��8x�5� n�ԕ�yi���@\��}y��d�6.�*#C1�Cz/����d��u��3yo�8D��Ʋ�n�T/�L�%�(��CRy��)�!���}5��hZ|�(�Z��n�{ǩ����+<�!�O[�T"Zc%e���r��B�P�f�`Z urW�C����[�J���g/t�=_yK�V�O1]�{�P��'�~o�I>s�<8}΋wxg[�s�y�GK�A�S��/�6j˩f���|���l.b0�a�A����ե��C%���GK�*l�/��s��
�녶J�u���;��/���,�U�W8o���7�y��2�*3�����P��H6]��=�9�E4z &h�})�D6�P�?����؇I!j/2�;�Cw����������9eM�	��*��5ep���AS�f
n$?#��-�J��e��ԻQX��Ų��!M�L���#15�#r�liB��ߴ�E�Hl��v�g��䢞	��`��0Ϛ������gbZ��M����N��k��h9-�A D[^���O��S.�.���>fN��(�M�B��`,��kց�m�����&�4,�1>�[�W�D�(��E��lD�>�A4$"2��!'�%X|��}����e���Ô��I�E�t7���6�0{��6��LE ZD�\(����[\��[F�I�6r��!�KLK1�[ *<�T�{Ҥgwh��R���^�L�!a{�΄.���u�G�C��x��[��)��Gu%�t����Ҳ�pd�#�8���~��JՌ������vߒ���w8R����
-��=}4!�y�´]enNA�3͔�/v`�@�lg#''�gԤK���>&�5<؎M�3�"JG��C9�k����[#�a���a%Mu�K���0�瓴ݧ�xțAo�4��ɺ=Ĕ�:��l��C������4S5���u�W�'e��G��Uk�վ�Qu`�^��\`&�\�5�Ԣ�����+��y�����3�M=�V���p���y^�b���ԶVyj��'\���`����v�9دD``�t�&�䧎!n����4��>����g�{����	����W��f�nD�SJ"G|P�͍���#�).������W��1����6���qP�4ɋ�n�OI�����Ȳ�h�e��Ir瞹?�y����)sf\�n�)�X��p�'�yx$9�A���b�^��=�]N=zΣ+V��c��X1��Y |y�RnC1�����p�^� �n#�+�Q�q
�)_�\T_��w�=�j����ˬ�$
���p��)��I)0'��:-j��a��A�����B�{N?���iĂB�����2,�}F��U�z!���xgY;�|7Xt�斐lY͏:��K�����GM<A���^=��J�~L�Q[F�M_ζbOQ�@������7(��jfZ��GM��S�>}	��B�,k� t�gM�ibR�B��?���*g����O!���+["p�澢D�����>ݗ:����i0�H=�+FfD�S�"�t(��/h�R����:'����ЇY2��j���"v�
��E>3Z��JY�� ������ �,�D�?e3��y��w�i ���5�?���:�^{���	����dq5��#�-�JsXྮ^jѰ&N0xXh<���ܥ��Ih�;)v2��9�x�,�bjWA������{�U�N[��+�=������xE`e�lD ߩr*�tȗ,����f�lw��#�a��8��C
/t&��/��X����^y{�����HD�¢��K��M*_a�*˯J^�
�W�.���8z�k!�U�:ǣ/[�{�~��k��V��f�%�!g&SVT�r&��*��*OV�|�=8�yk���s&�F0�3��KHq�-�5�>�W�����S
E�>����q1����F��CS՝5&�M�ɵGvN2���=�g�a�8@(?<c�qv���5\�#]���*���t�
PT&�h��4�-t�:�g1v�����<��1h�l�����SH�F�U�K���f&,��V���8����r!-���œ��0"�!@Ԙ��a�N��v����Z���~���)��F�-�h�]����?��~����o���9�O�W��J��"���syG�]�
.�h5 b��}?ԑR���6��L���ݭ�����R�=	ل�6%+@�y��dK��1�Ly� ���ɹe��6�R�3�4�I)g�zR�rI*��<��b�>*��)XK���Jc�^:��1�[���Ф��[�0���쳩	�~$�tO��� 
y(����{.A��#��H����(@����(	� ���7��ϻ�^�W��<�|<,J�
�s�P�5.�g;W��ȫ����48Z�˰-p�t��4������7��!����N�ݼ#?uFxHs�P�]����oc1�$����'A�q�1r��G�O� ��N�`��!���纮���S�A�Ȕ�Ԏ��'�h[�nC�����u�/�sE@�X���v��<ߥ��yĥjtøO��ɫCCՅ�ljԫ���%X�'�,`��zl�ڲ���]*�S�p��������p��%,������3F��U��Lߛ@�Z�>��_����-�9���'sS�����[�Ae:��ξ���>2`���B��EC��>�!�(ɡӐz�7�l��D�([�E�y �v�b��\cv��i'��A0|h*(�@f���O"_�N2�#i�1��E��{���V�<�Y�4�=z ͘4�]��wQi��)FA� ��ꚞ�W�?�	��hǬO�ZL���Bb^������U���F\�A5����xi/��Ohj踾�	W�����)ky�ŖC����pJZ����c�����{�H퐞0nwP��<�14+�Pw�Τ�D���+� K*28�k�X`�
��'O�4��Pu��Rf�o����@{�D���W؇��!�>���>uz�L\5C�*���[�h1-�/��-	��O2���PJ;D�H�����Xk���IٿmN%F��.:��̄����C>��d�����y���<��@s�d��<�[�ƨ'��wC_��3�ԑ+#�7�Ǔo��	,KG�hܹ���60�Y�p6��g�|�Do�u?جV�c�k�ӏ�,��j�%��v��9(vD���G蘝��<�[J��XG�3�O����0({��6�7b!�Oqȓ9,;rG�̇k�����M��=P�$�JG���B?r�}`*�����F{�N@��ٯ\�?̸��a~nyZس*4�@���j,��j$�Ɛ��ư�G�h���*s~24�� ��dL(s�y"Is38w�� iz@�8^���Р�ua-o�հX�OWލ���D�)���)!�b�d	����������6�uBm�<�(A�����UH*�2mw�&]� ;Eɐ�Y�b��5j�LD�C�C�}@Ƅ���H��A����0�ȩs9� _cP�53J6T�{G���L��֯=9��Gީ��iS0"o\e���$<��K�,V���;uOk.'��t^=����F��ż^��o��q�f�Z�YC'Ń��S���5�N����	s䳧Up?M|&zjf�zŎ��>9jF'MǷ<�s+�K��bΣ\�%:=�`d��G�}~m�lK@P�vw5���gH�~������v�s�]�
jQ۫C-�G^"���B0��m��b��.L�4�L&_�iGs��Z�s�f���O/
�H�*\sk��{a����GN]��H�=���G�z"e�Wc��9 �c�P[�p7n����-Hʹ;��w� ��~;��Ys��0ڀ��� �\��3eѾƽ�s3�+5hz:
�N9��NJ�,:�&X N������.e�e1��A��S6[���P���[�� ���s����
����,�*I<׸�XJA�"��ݯ�q���p�y��>q��tٽ�9�&4�ɬ�q�Y�r̿ZR����p�ZpC<�*Ϭ�F�)�e��n�M�>�3ơ�*��P��٤�U�e]mDL�&:�'��^ �g�s�3��Y�g��=qeaKG�. �|ya�\o_���ں|S��,x�th��B`�#�b�?��E*� R�ug�PX���â�����&;X��g�e��,/K�`��5��k��ݬ�����A�hJ]:��	nҴ!�}�77�`�OH�r\젎7�Sc=)3�FI���Q��R�L^x���j[��A�ëb#5MTw&��R�[S��vRD1&j9��bQ"��"4ۼR��*� �i_����2!`���nZ�
@,�D�B��������}�[@+�L���5����$���Tm�~L�� �d�Ձ���~eZZ�%��!>���
J`��O=<w���L&�x�����b���'^��� �4��Ņ�HMÆ�0f�����i�s�E.)U"������|���&�K8�T�+z�3~�$\a���"���A&v�ŷ�n�z+�[ԍ���"��pH�C���"�`v�eH��R_5&�R����'7u����+���w�v�M��8�!�1i�0)�1o��W%��?B�"R"����U��d8W,eJ��<�'����(qo���n"����]�C1~�?������%D9
��7�a.�{��O��;�,���2G%7�A���ԈԙB�e�7Ï��������������̓�=������&���`N;�g�{���3I���$!�.`�I������9���WT����V�</���u�t3,���7ma�p�O���C+��|���1�/I
b�[�	�T����z��\�ׅH,�p��s��C0�7������:�J�MBJP��n�@C�&�c9���|alɌ?��D*9�p���q�����Zt�y�G�\0��iY2���3�T�Y�P�����@��E\��㝯�;.詊~�6nrT�ݟz�����w���ǽ���'
�]�#�ɢ]I���5�Z�15�
��w�Diĉ���U�E�L�d|����"%/�
�d*9���#h��=�捸ᴸ��j�`b(��گ䟻F��2�?}F���7i.�w�cR���fsj�Y�vB	�7*��@9ЮT��ꛡe�s�L�E�����{��7���$+�g�І�D�S�G�z\�Qt:K.{m~�SN�Z��]�v��NM�j/� �EiQ3Q��/��J(;s@yA��2o/�t,x���h�#�u�� Ja7�e�k�+n\ LGR�W���K���M�{+<��C�,�/�a[w�����(����U�o�f���=0�T�%��[N�`����m�V�J�F�{M���/$�_�Y�˗ ��𽂁)��1��n�Bu���7���^3]r,O�C��n�cՑ^R{Z�52�ꌩ%�j;��
{��m Q��Ou���F���b���M�MC;�mD=�N~
��1£�&.QH�%1��*V�qc0Ȯy���!L?��F�$ex=�I����A��ҽ��xTZ�)���2gW�MB�AS]T�TN�ȃ�*6�>���YGBt���k����C}�/�WbS7yo���<C+<#Řř���D��rc�;�RS�) �x��|j3�=q�T�^�dA�	�ґ�`�C��f�˾>0:!���ﶛ�'6}�󥯙^3!�9�/[���u>�4����S+�!t�	C}�c��3t������h�r@�f}(x�i�9G敏�*���3�q�<b�w����t|�bN�\ޢ�*��Nt�E�t�0�!��9jC:m��x�Ӳ�DL��Z�M�·��S80D�"â>�"t(6���híʁS9�ʅp�R)�C��l�WbM�ީ��H��i�?{N��ƙt�=��P7u��eX2��v�F3�G�<줂i
EZ�x�X;�����v_�Be�/�Y�}ȼ5W�J
*����+��ƒ\dSg�8�f���э	a��^Č6'\q�4��D���|�I��2�h��"�pWG�h�L%���,��09C�U��{��	�6Jv��?��`� �O���?L�1:�h�N���~��hAd-'��WQ�F�!�<_;�r���C��lx�L�Ӓd6��XH��9z14`��4@� �/�m����0�բF>9}�n4�lor}Z,��߸T�דgt)�	��pYL�?���eG�u�����]H�J�,j�F��JV��үiy��dA�9^�b?�̤���@��`�i�o�#�"N�ТA�����N��^������['(G�7��uܔ`ь\]�z'�jj"LY������K?��I
e�&�b	�՟@Aİ�r�قp��Ghn�Ou}�ٙ�/,q�)��#��HIgс-�I�Z��wS\C�_#J�����B��ϊ�J+�>�M=��A��Qzd 5��ˑ6��<O�=�L{�!�3��;MH�G�)Ւ'����F
���E�H�E6Z�F�+�C��)Jn�����p���ݞ�B�5/�=�!�g3�U8<ı�Tr5:&3��"صr�$гdF���:��;lՋ�uΧh��	=���R$wlWDz��U�M���C��j��迂r'�.�l�� ����`�"�4���ʋ;Iq��s�v��P��@k�]���^R�������h3(6���\q>K#m�����{M]�þ��o�D$��/���Azr��S �#�j���;�]J�%E�zn�:��l匙�"L1��ٵ�x���I���얪����F�,���
i��^�=�^F�TKᬧC�������(f�1�n]�{HLde#|��f���>�v�E��I�P���*d�~�7j�j�{iŔ����'�IC����v�����_����f2��l���`��	�f����gy$=p��S�x6HH�;�Ղ)#�2�>�*�����8P}���(�e�6���$�_[$���]�y�ۋb����K��9�'](3v��,5s�x�Z��s!t�%`$A��:��0��hlWU�(�FՖ9t�$�x}�V�A	@���W=��ڃB&�%=��N�-k�TF�P<j�Ưr�Ol;.e�Q�z4u��-bIX6��$��Nŝ�`A�r����T�V?�-���CN�Uv�d�w;ʈCh+8���3��Q2� �:#DkC�uyөK�\�j�t_K��{O<������&,N� UpBK�Y��HR�0o��`[Z#D�r`�1?�qk_;A��Dy��|l���	���-�牞�F�nf�ò��{3��t#�<Eqy�.A����f��@������4��k���'1�eɥ1��|Uk��T?�]�������M=0kO�y��R?���j�L�y-�ƻv�qp�lwǝҗ�d�gjo���x�ZNg�	�|������L�A�U$)�>��1�+#�~��'�/m_�xFAO:VR�U/�P��)t�g��L�.��-�'L�j��K��j�\�9�)��SF��cG�ɳ�6�I��@h%�hr���% W)�����-���~Xv��'(��K������]z*�~�-��c�zU�":��؆����y��Z�u=�Q�q�8���)CÂ�JcP����tօ�&j�ә]C :B�����O-�����w�掗�ўk�j8{��!�3D(�CUV���F�F�Ɲf�B��5�	�qf��~�U}�D�_О�&o
��
�Vmd�r�����v�G�R1�=eO&���E���I���7����]
r��;J��ũ
\���6�ʼ*^Rc{��t9�I�s�EY�7QW��Y���ch�0V���¯)�����F��ָ0�]��$����s��x�VL�h4D���;M�T1e87~5j; ��
��&�Jdłe�\�-3 X�K_����z�� ������PSDV2�
�O[ `���U���[�DIyR�ͯp
���?��,�B@q~ԗt��e��,Q`*��>yF`�նӭ�}l}w���]18�Ϙ�R� ܑؼjo�4l�~�nk$�X@��̽�,���&c<��j�+m��kʜshz�9mU�,��q;�'�@W˿r|��i`��� �Z���ͬ\�����x�m&	��T�F���;�'#_���{L^V2��I+��E�"�(9g���US��}���/<[��.�7����oeq�na�͝�zGȋ���;i/u�n���a��}�0�X�l����SF�$�1�	���+�b�����L�-�Լg�E��}�l��H��cfO�"ؒǵVńle�����ҕpg��4(2=��6�i��e��z��\=�U#�Z�)����b�%ۙ>�K��5B���hRNA��u���T��譸�r�5Y�m_x�V�-�艣�̹]S��֏�@4�]��1�1~}Po�S�!�P��[1�r�'"˃�w�ON���~PC��Rb��i�"��,��T����fu��@-�Y���k�G��WG��2�����YDXd��!w�t0��*�kD��fI 4�S������N>?��b餹L�0��m�F���9|�C��[³��Ȇ{�ΟU�_�ҙ\V2��2�;Rh<�xII}U�U����^�Us[{�n͗�~����+X�D�wj��Ԏ�����65�q�C���O��4=�>=+2G�
�GFj���l��W��m����H?K������z�޵��Y`β�t[]�~��̟��D�J�����4S4�D�s�"�ߴd���ʶ{4s�Z㋏@j?�'2��e�9y�����[�-HJ��ِ�%|��:,1��FY�D!&���.Qr31%y\� aWF~6O^��Z����zi{*��5gꀔ��f�v!��Y���a_� �1H����AL�q99$��@�6�����J�z�w�=-��y����^bY^er���{���%c����`�ަ����o�˓�����բV�ñ"v~��D��������IF�%�ֱƕ:�+��֟�����e4�	}����������C_Sa�Dl״�6��	��~OCR�"	��q�/׽d"���6���4���\9���J��V�]\Z���,���}G��@���(	5�1�T�����Ph��`Sΰt;�P�SU��i��Eu���������#��{�j�%�#�����S�E�f�����q^J��+�}����ܛ��*|���:U�
�_�^�	qD$�gէ��Y���<	3eY��>ྯ�ɫ�Y��2 �V��a�bJ<�;��?��s��b7R��؃E���h��y�Q\�Xh�F�K��A���^�U���^����{�e��{���{�%r���b]��`��0Ns���i��I�w6Z<jV��&y���'t�C^�5�mKc1���؟�Z�9��K�(��;����P���Ñ�)�d�S��*�Y&���٬3&�|�ݎ4�"/�ua�՛m�%9rFr������$Pe�������`�a�W�vU]�2��r�i)ՅcH�C�C\DM�-��ܦq\:DP���*$,7�Y�x�S�#D��f��C�{/�=I��^�8�����_#Ǥ\�e���l�/z�R F��f����Û��V:��2����!_�'�աꢢm/ ,2%��m�^ڹ�,��0xb�Q(��߽|�eב����g�fd�Ɠ\R l�L*-
zB$5nc�wʅHT��M�Ec�f9�pc�'M�	N�VE`���	c��e���?����W��m:R�Bͷ�^g"(N�3R""��ib�Z?O��Py �ѧ�J��(� MY-�-!��|&�����
捎A��X�Q#m��x^u��>�;�	�#��f��^�P%X��B����ؽ�)[�E	4Q.on��A���)�mo�n�� ��|��{�wtx���$���!2	�AP&�FM�m�[���L�����@�9=럵����L�0��z�Cp0Xw�goO�?��y�0yh���-~ـPk~ǖ�����6��1�N�}�-�����:N��^G�Sķ��/3�V($�;zD�+��R�?s��j02����;�6��S��B�i@��1��>n����/"�'�m=GS�����^Dɦ%����T�_i��������qM�Ra5�(�	1٭s&1�8�
T�����ֶA ��Qk��V����lDJ{6��sH��i�RA��I8��.��̔�e�G�{�"�˲��+�>[+t7�5�
S��rK`�F]��(*�n/��H��{��Ȭ�|ׯ� [���_�Ӿrgt��=/��.�/H������N��[�s����z�?��~�P�� ��vKO�^�['W�e����Ҟ��{V�7�|��k��&(t���,�g8F~�w~�!��������� �K\q1���nBGo?fJ^߇ �G��U�� n�����A>�����C%�g�{h1�EǸr��rqXY$���ŕʝ��n���A`��Dv���<��51�X�����E�tM�=�q�{ȕ��Dm+�׽�G#9�w68��r�N�c�A�RA�c �,��t�{eC��C`S�j��y����ѵ*Qp�3"aj��I��Mh�
�
S���)�1%5t��k���I��L`���o5�A�N_�<N���ܯ���w�h�R��l�/l�Y�1�U%yB���Dl}@�C�#���?��=W��6jL�t٠(M���2�m��͆�I���]��y�W�</��&/]o�QUn$�T�}T+Y�hEDQT/���*b�Ru`�
2�$�{��v�GHDV0*Q�n|_2Rq_>F7���;'p#�X9��"�4J%� \UA��ǒ��׎��:4�a�D㤠�4�
۾u��]VA�Q;���Zjx�_����2i�����;BuW?��K��V��ҩ���ͩ�))2����)�n��i鬆j	%�6ߕ�5�g����4)k�rr1�[`S ���ÅB��i�/N������ɔ���зI*�����d���g�%�`�M؟��j�IأB��>V�D%v�?F�Fk_R4�X.�T$�Ϛˢ=sl�iP��$|����6vM�k&MO={"��S��I}�.ϯFܹ8z)U[����>�e��f��������$.hEl��ϛ���XRr�O�C�@�кZ�	�h���;Gܵ�~̳�Z`��\�ߌ%'r�������%�(����<�oKV.3�
��Ϣ�is��ͥZɳs�k��F梀 �d��ޥ8�)����:M�Q�k�;�z��{2��vG���W{��7|������.��)�#�fZ�$�BI��!q\p;���
�-�p��^����Ї4��*J`Q��#c�%9ٹ#iJ^K�ڈ$��.?���f���w�_��z�ʈtBH{�����6��~����U)n���pFKs�`� c�R��K��dm0E�{��'�g0��Ӊ��q�D(q�O_��F�� P$����t�f*B!A���F!���,���{[\�M�ʸX�R�VK@4cSIN�/�l��z���Z	G4�k��lE��n�S�G�g�b�������	u"�����#2/�e��,����-�roNnT3��Q�� ���,�I�����I�Bܨ�X�S���I�6M:�\)sKP5���V��_�XĿ
�S���n��'������0��kᓄ50�K|�e)*?�w����;T|���Š�w�#(�B�4�E��5+G*G@��y]�e7sJal>w׏�����v_��Ԏ�웉������v�c)K3���(滖����H������D0�`��ɫ�N� ��E�e��3z�����g�U�v�(�	��t���D�J�����d�����#a�ۦ�M�sb��M19y�#� toȕ~�F3NKH�|%߈\�_�߽\A��}���Ah�%*���,%����uC���^��l�}������T����Q��{6�uLR�h��١���uʫ[X<J��'mĆ�����LleaD�VӤ6: K�|Et��b��� � qQ�W��J��+c�ٿ����aVcV���V�R�����s1��O�q�DH��o�:&~�}܄'#�����8�_-a)�0Q���@*\*aK�%fG�&P�RF�Q$�Q7�W���հ �01�|�<~w�n��3�D���o���$���Ot�Mh�C�أ�Xšگc{v���7�E������I8y��CԳ�Ȝ�����q���<���`�RƢh<�#i��6l�v�);���Wl�qAr�K�a_�yh+�VF���]��B`9�f�S\�s�����lGTfT��$��>'~���o�6�n��~\���ڸ�4���K,�$�[E���&rМ���(�\��5>�+�~��;8b�Es�:�|�D�|<�Xڎe�����Y��+�~��,����u��8�P����n��]N���AqW;��;<�	�V���ȼ�pٶ&Q�lx$gp�w��G�����tP�Ϛ���\F�����"8������+3)m��ڦޜAC�9�}���D��Z������*��(�57�$w2YJ��ηV(����ՙ����+p �0�[|a#�q�e����yf�XV����9A0�Ҁ��H�/r��^֡3�]�)�ئ88@��u�|��Q��ف|m<��6�P -[h��'O�� �kA������C-՞�B8�����-�eQ���L~��,�2�R��h�G��Y�r�N��\f�ՐM��߹z�%p+���E�W��������:�8T�����1����wv3���'T��>�yl=e���a���9�lQV�,�?�9Oj`��l�AvM=�ZI];>\�打�H�
��%�*
뢬��@�sp�d��=d��Z��G۳�U~kE�F�C����
xВǐUvzŎ�0��K}ZS��y'�4��0��������I� ��������9r����X��V-ZP^_�y]��S
��i
1��
�N�	>�Z��n=�R7|� +��s�B�[�q��F��爄���]�Cا��*2�5#���<s��&��%��K���!2{W�mܮ���xv9j�C�4�lf#��L�Y ��c�(>�j�gu�e?�Ze*6�%�iyP
7�&mIbB�D_4�b5�:�/֒
7��֟jZe�L��U���zD4���O<y5�msD����s�A^UdN��-��|�EX���"���]��_�\����@�Xk�F���.��P�*�_T7�����9N#`���,4�?<F����,��C ;f��I��:�E��ѣ<�媅j�o߯,�7.y�Wq���/R�/�f��r�Y��{��3���#��f����~"�IEYH�'(��|G,��`̣�X��z���°�
0�*�sWs���7W7�$��v������1����_d���@wN�1�P<j�P�8�䬌�/�+�㽷⽮q�7��袴Qq�]�%�w��g�,��K$えz�	q����CQ��bM[g~��w�ˈ:���k�p�W�q۞V�����ϣ"�C��H��w��#q/���q�M�YH����0�	[�������E�ю��g ��(�;2ǲ�"y��O���_�uiy�#;���n`	�ig���z�>�T�]���~��o���#�;�f6
��dF(S�����7^�q��׻B�E�q���8��9�|78F�3���4+���p&��"��qJ��J����5��HZ�[߬=K��{����'a��n�oh�F�}9���k�&+�W4��ڶ-z�{e���|3��b�-��B,���{x1�m�t��|�Zo�h�IC�� ����"�j�tֱ�.��ff��GhE�P6�ûn�9(������m��v3�}���<MT:��<�l%� "�4�1��[�A�򂃝�x��7N|W����18I+!`�8~ʒ_84H�:�q��ۏ�i��}��aE¹�>���;:��38'�&2�� M����%��5r��p\�A�2����섯�yv��YR ,:�kfH�8*���K�"p>���*솽�q��U.Z嫼'*��ʓC lS�wq�~˾���;�F��DV�>wy���\�틐�X������R&k�礥�DH��b�}o���$��@W��;�d�hs�	78j���$QR��Yd�4�.y�P���#�?zu�,��ɹ}D2 5���m}��?S���=����k��jO���Z����]dX�)ˀ�ԢܷG�<��	�DpPf�̟5������*���n���}o@���𩁢�BAj;M 
%�Ct
3�ї��dwR!0�]�-]�����Gدus�-@e{��l�4��e4Ǿ�挅�/FF�t��hb�z��egmߩA�Z�y���n`��w�M���㣊}�g�D��I���s9?�Q-�&��ݳ&�L'ٰqĄ�?p��]e�C�'Py͙��`��6�꒸��/�UC��Qxe��1>1sn�N^�9m����T�n���Vjy;#��nӲz�8���-`���+C,����8XګF(�fDh�\OSw�)���ԯ{���cO��^qY�%�w��2K:x�t�?"4���[��!9�i=F�(�@�m�E�`ɝ��Fv�+����ADA�\�H�@#a/�f���.3;?e��4�>�d^�ݼMm���·��Ln��gg�j?ie��VS�o�V�Hu�,%͞ﭓ�K�vj�ʧA<��\�Ejݞ��Zx��P�U9��Smˈ>҇a�׼:= PY�����-��k��G�$ۼ���!��N;��
�K�=�m��a!��R��ȑ�̨��lL۵ge�y��w���i	c�<�i�wOP����p�vhϝ��D�/���
S�ߊj�Ft���rAX�O�y���-Q���j��A����d�Wv
,��q1v���=/oz*��� _�Π�;}��z���X$��?�t4�ļ�9���
6O���J�p�-����v6��&�K���ź�RM3���f;>D�a��Ӆ7y	��[�r�}���d�$S��| �z ��[QX�lO��<A��W)*M��X����U�8!���荇���X������ɷ��ʮ�@�j;M���.,"g�"���i��q/��T���H1��G�o_�����N�u�ȱ���2O����z��q����h21��z�U-ܤtA��j���Ňz^hDZ�<�k��!�������I�kY���v��o������"�qӂ��9'W������¾���<o��� �������J��FU@�K��_8�V5��Ni-�vy�W��܇t�5���훽��8��g��PA�{��qk0�!�����s���\mq�@��/�s�[!�%��-��D���Mm9>���������J��9kd���Z���@�l@s2VsAS)i��iM���n�K~��7Уd�tO-������� g�DH�c@�E�ԕ]�q���/�0w�\b�`�H�>���OŮ.w�.ڠ��ImO��ݏ�6pa�l��j|��1���GID�)��Lk�Y�D	������6K
ֆ+����fPw���h��q�����(�
�jɩ�kG��(���p�y��h�:�˕��p� ���[#�=�7I�c�~Q�����	7ym�L6<���BI)1+��6�vr�]�1�fo��1W
Hd�?}:�CuW�"Q�+X/�W>MG�r��D��x@�d�3��A���H��J���B��3A웩U�ʦF��@s!���\0�R�����碛QM51"�Q�
���kg�8^��T�x�N��^���@��)'d�q�4;�#�g�!��������!�m��2����p=|Q�L�IU�/\�&a��S�\ug��2O$˒���.�T�`�����7S�l��M�ޮD�gt�g�<�7��*R6)U���-�Z�W����B[�l^�UOxؾLY�xg?�5Oz
��uZ��E�)����"��G�I^��Td��h0u[�E�A��b�ڟ'G����bV�t=�g@��G.��1l+vl�8��?w��o���yqj��4�����e9,�2Ƶ�ӺS�������@�Mv4>X��3W�O�=0DC��q-��|3�C�^8V) �8!x61�ބ;�z��
�a�&;(ϻtK�[����������\�$E|��,��?�|��wH�R�#~cD��+�M���xu&!�5f�N`ƹ'���uuӕ8��>钋��o�=s�m	L�C�<c�vi,�j݇�À4w��/LQ�������a�CC�e����@����/:=C�7��O<��_Qz��^�C�����!py�����
/�A� �f��k���U��l9�����j�-�\|ʃ��Z~��=L���&h�~��P=�Z�^����8Pgg��"��6G�
s6q7bN/b�>�����6B�}���Sr�&r�yv!���FpP*���_k�X�&� �twW��K6Isn
r���>�%��H�FGEN*�Q������=ZH������A��!�F�;%�R=�qe�N�����]�ΫC/�On�L��j��p3����w2�hD��z��Q��լ�ɑ��<e���r9둨I�t,��e5D��KJȐ$�I�_Nu��.���IϚ.H2wR�G�V�U��� s�fs����-����s atzc�Ϝ��b�%@~�8�Ê���f�x��x -��?4
���0AWk+|�l=n��ք�XBI�Ppp*�{Jv�}{4�����3��m2�	k�E�ѭ!bPG�6n�jO
ة��B���l�����y�e��H7�z�<�K(KZ��O�N��k�[�����ػ%W���m�Xо5�ty�6РXل�lh�ע�������X�9���_/�e=��ҵ���K�q�4�Z[m��Y1x؅niD�̚�_1_!�۫�i8"	�8��+#IY"����*#�t����Hͣ��j�,����U�u����[i�f�H6�Ki?q�8c�O�K�7�8Z�k���6�juoH�he�b����Lf����U�;s�(�-$}�m�~I�!qX�z���$9��g*��p�wZJ5��Je����}<jN~��D��/�|[��"�\����(����.���Wh���G�p:d���A4����<1��zV�Wr�9��ɨz�LW4��_1��v�Vב;�KgU%���4r����O��ZzD����|r��G�E�Ugq�����3~(cq��qI>lʊW�y#7�ǔ��'`�4�ɞe�Ӣ}0"��H7�q�? ˘��炧#�?���F||��K_�8`�"�e��2���/>��%C�I��v�G�-Q��A�I�su�/]���Od�H���-$`���̫���o��$$P�]�+dcV1����nU����G�ؙǵ��y�Q��,0�P
&F5%a����_�rRK��Ah�wD�F��9_¾%����]���H-���P0Nj�C{[A�a'�F��7��
���I��%��%�.ٿ.i�n�u{8�?���\<�����1���h�a"�Fw�(��oV�`|����;�0�=ѻ��%���l���}MIc0֜G�r%#5q��x�s��&�W���/�׋�TQ�0�U���yRj�W�T쪘�Yۀ�w����@��v��4;&plfm����b]��f!�����)&�E�W�U�p��Y�ͣESś�&��D��Lܡ����<eH�+���4>�#P2U�2A����T�Ks���I�q������a�*|�L�:U�jɸ��-�>á�K�=|�g�����:Y���	._r^�Oa�r_�C{Ӭ��,�0�k4��iw-n�>�>���>���0f��P{�|�� ��ȁH�~J� ǿ����l
�)t��0���W�2��d3Y9�\���b��p� |r���/_�V,$Z�u��W��\Ѫ\�jC]10��@�V�����(�D5��g�N� 0���6�T���mr(��D�BѺ����*��|�JA.���� �V3B��)�|���'��u�&�I꒚P�  _��h�j�^C�D�c�J��I���pNC�=��(F �-8��<�'�iVtH�[�rM��Q�-O�� �[��^ԸC%h3�o�=tE0�J��bx�&��Qm3G���:S��ik��;�i��UDa(۴A�
��7H�;3C�✉�CM��[!ɍ-�W��D3"��f���}٦X�qI�@ɍ&�{ �q28g��~8]VP��$qd�R1mbs��3����/׳�D3g�����i�{�%_mn
�#5��Z(�)z��pjC��0�MsS�i��ee�z���0�ݩ��kx�I��V�,�V �:�M�^1���@Rk��Cb9+���]L��4s\�>����(��!����Y�K���Ή)ε�lP�{բ��B&��q�-oU��.�/�O+��^�^ZJ�,��'z�����W?�k���o���ٳ�Z����)�\�w����i�,�*,����^�}�����U�_{4�d5 x)sd>v��RY�s���w3q$V�t�7�\M���`����#�-1����AȍX"��y�房s?�pn>��^�g�ÿ!1?y��Z8MC*�;����w=_���H��E�Q�����Oj�1���^��?���.x��K�lɾ��9��w�}�#p�E$0R2C�l���)�ќ���P�Y�7�J��A�����p�*Cﳨ�%0���h6�c?�K���ʖ � ]TF��z��xNlʜW�_nTI�D����Q�gj�>��i(�˅�'��gdׇC7F��󗷸�M���I3����WOiՔ��S�D�
�:�O$C�����%A)B�F�+�*������l�ナ4T�.(R4����������ެ_G�/<y�<�!C�d)b�L��PwH��#��_Z�������l� |��a��Zz�� �}r��y��p�%�
}��"���ҷQ�{@`T!�5	4�MAES�z�2z���a���L����9E�NI��$8t�������m��6��~ܫL�W,Y�ɤ����9�n��#�Z� ���+"R������c@<Rj�m���࿐�#���ӡVg��wz�R�s{n��sL;؝6�Ȇ&P/��!��W=�i�4��|A~ȗ]�R1�BO�5x��� qk�=�]��*
�]�1��[�)���$e
�&���|�\Iu��[�aE��*O6����� ��
-�f���+�T���ЌlY��`s*�*�0t�v`P9���(���t(�u�QL��3m�?���z���C��5]����p�ݸWY�\4�0M:�0�ظ�Ѕp,Z�_��0Xˉ��i��{�������ߝ��!_O��K+`��́{�3�*�n�^�
�E��F���ے�r���A�Nr�� C� �f%�%�3��,��9�f�<��E*���>'���Q��IR��hL.EP�g���oZJ7t�����z�G85���	�	٥Au�����T��  ������hOS��3�oڳ;h���uiȏ�2οcG���F�p^��~%��rf���-ǧ�?C ��(y�ܟ�,�F��s@)���������h�]��Vf��f@b�����Ȍa���������+ozGҦ�S:ş��0�74�W�c1����D!���r�9�}��1KmW�$�ܶ���p]��ͯ.��Gg�l܀V��(2fsx\��'B��(	��� {s��x}7�b�p�sά�:��J�x����p[iU.4e��T}j2υ	d��;�.���d�O�h��%���� !�j+��nőplﻑz������dq@RfD��!u���~u� ޱ�>�L_�_�\�<OjT0Id5\&���-<�f��.K���s�|��� ��<�h��y��klB�x.Մ���	�(b��n����U�}����%�)����&F��4�|f�v��M_f)�+�a��w�J��F���v��?�PNȎY��9:
�]��M�?[�>`�W=(���}�>ǰ������#&l�/"v���4�>J"W�!H�X�)J��ϥH��.�m'���D���I����H^��t�Zd�|��Mn'��dG���[}�p����&z���B@xm:�Oǟ-	,k�7�P��C�=&V�g��|9�$�r4�W���"<��N&O'p�9'R�B������2��}�`OZ�}0v�ed��7&��C���1D�gQg-����K���L��3d
��a�(�b���R�@�x:�:ɬ.���v��õ�.'J4@����'p?ؓ��8rٙ�m�������0Xu4��7f���{�Sk �� DE\"H���y�Nq��)�r�����/��Hhh�<tR嶰�`��d��`�s��{�����}�p�JC����v Z��& �ܳ��H�|�د3l[�\P����� �R��Y}s���?8��D�h��!
�p��b�����"H"����H����{h��C�����0vu17����~wv���B'�����4���IV1l�U�jPؔ㹗�\݂�����Z2�'���jn��-8�7���<�'���U^�p��f�<���� B}E��`��#D�N2�rV���Zi*�܅Z�p:N�����Q�v�X��A[��a����$����Ɓ��q�O�1���T�ڲ�K#��Gֆ֣7�?D2忶w,-wo��xoYw����s�פ6�dw���v'w�߈�>([Jە��I_�#��6k��YM�7����v|�LҴV�L������Q7���r�s��Z�fr�\~����N'P��������y� ;`���^�t�JV�D/R�p��ͮ'�36�u�[c3��~,� 1c:Fϳ��(�h���Z���J#�4�L^�{�h$z�n�?K��� Q9R�]�&^�8(0��Ȋ�}�W��r��7���$�i4ǵJ�٠ظ�bC���|��jv=�'r����URH���B`�8;{K��9R$��?��ΰG���m��V���R���{�/��
K3.1��$Ї�I���`��F�K��(���0M2�%��];>ʞ ��Ʃ%Lk���Y��*��
m�7	k)�j�kEǈr�6\��,����:�����fn)"(���5S@`M�c��d��d�9ĉ�302�7nj��ӭ>a,��P�}��U���6OVi��874��}*�uT@x���+l��S&8�H$if��2{S�3~������'��k �-�ϯ�:���� ��1q!�D�Hw���v/��3���~ xX62J�����
�7���:h�ܻ7�ei���z�%���-��`^
=J��?8(�-�ɽS�<��M��\�W���Mk�SH�3���Qh;ƀ�Ga�F��5����D,vp������d���|q_!��z�Fڌ#�3�%Sǜ*��:��D��
^����	��s:�A�`W4\D"FbR\�A��Ӥ���	%X���7MhĢ�l� �5z]����I��Gl���k�J��8e�pcB��
8��?u�"]����؜)g~�C��Is��Y��*�'��7��5�k]����)7����,d�����2s'�B3��n�V�QU敼�J��3O��9�;�y���=U�>��T-f�V`/<��t���&q}/�Q�]u��Ֆ���'�aU��h��C�{�FւR���E9�u�(W�F�Z_��	��f(�n<_V�*@��z?�m�	�Hn�^��q;��-�T�ʥ�쓡�᠌��@��I��;I�k_dƠ���h��5XQ-�zH��3X�em�b5~����D�ۗ��:(VAȯC��� 5�xc>�KG��|�6�H��:��-H�	�,6y�#'O��7n_�O�fb�3�����˙c�uA(�#����>Ӂ�'j�&I�k��:�%6 u�d��o�ʏ����(UA����q?�h�v�@�dX���6(�^���R�i�ؾ��w��+'�q�$*U��,��v���p��4�C�]�lFn�m���u�A{�����q�*���s���.-|ul��ݏ�rt1�Ώ+j���6�[�+�G����R͔�����<��s$� lB|<|V�oۖ��?Wڤ� ��`K���	��y��A���<�SL@$葧Q�bq9+a�g�{D9U?�f���鸔����$��$膫��t.�ny���I�q'�{#����l����])�%�.vI�+�EB�#'�ԁ�y�i6�ɱ�sx7�[h�/�&eRŃ������/����)���������/y2$T_��у��cl��
�9E.��ZY)*?���?��:�.�*k�>c�OW��q��sFⳈOk\�����y�8�\����&
��T󑨲v�
�fϟG���1*b��Dϋ�j�Ѩe�^��䒘�	���܌��N��2�;\�鐹�̧8���[{����Ё*�wi�L)��?�u�Gv"�P�T��Q������@%>-����!�sɨ%��b��A����Hpn�G��LL%�Sp�lE'=Ħ�#Z��R]�*d�y/��,5*:]�*Sԕ*[Pȗ�?�IA#Q�JAЃ����B�ͧ�(�G��i�,o!sM�w� A���i����L���^��ߎ5���j���f��Q~�Z	N�B�v���q���b������<+~��K�;A�
�+N&[��;(>	�?:!(�d�6ȷ�y�v^�$򶥱���v5�`l<*�D_�	H��o�3.'�^B�-~׶��![mo��AC4�����I�J)�����)�=�j� !�(M��zj���t�P��mE����l!I*>^�������G^Jz��q�,�{��w��kEֹs�d�p1R��Ҫң��OV&y�2�&�H�V�^�"�"�gI	��Zf=��q"���XVNl�kg���Pf{5�>�P��A���Ѕn݉jG����1d���3g���,����~K����bP7l
۸r\}�~w�~[&x����p�����R�(�8{#*�n�)���n7��}ln�S'�[��@�%L�YbX�r����MJ��G��9�w|δ�_�!"��ɓ���q���/�S�KV�`v�!fܵ���1����)�ʃ{�=HGKg%0�ƃQp@�
��G!�+WZ��	��t�W>�L���1m�9�c)��=R�t�	8mM��o0�J�Q+^�YkX_1EpY�'�J(������8*�򷚯-���<�Z����	���Y�dL���)w��1]��@��j�#Vm��:2sۤ��
��#.��gU�V�d�2r�+Y�m���ߍIrH|�=6�P��@]`<_���b���o�$�:Fy��X^�	�%�X̌J�o�?�J^o��!�}�j�"4���F��"���9ہx���Gm�Ib�6F���-4�T��x�"��]�M_��u���]�KTy?�'3���N#8h��7�nrrm]�� �H,�2�i�T���Pb�^���3�e�8Y�g�4]����ǋWmj��:�`���c��!���r���gl#J꼷t$���кX������:�;,��P"�P�M�
����@R�� k���z��4�ɼ��{;9�i�e���n�/�i���i���o̽��ť�$�v��S'�4��`ζ�K�W�Ah�?}=�A>������s*(�Z�6���V��NH}�pl ��$߭��$�z���� � �(�$Ku�*�ey'�B�s�}:�����Z�C�����Z�}�4�q��A�T���kw�l��|�6-�+g�}��wu��&N^��G�]E��gs���Թʨ�-PG��#�V��<���7��3�-�0q���h?&�������)3ڙc./4|;��l�om��p*He��>���0�A�D]�h��Fw���x�$"�$��7�O��_����Y�.�;>g� 4.<ȭ���1��Wav���b|�w�o�)]K�]�a�"�;�a�^[ջ(�߮ -J:�s��?���u�����%z�=(_�蟫:
���6]�^t���S�@[Č>���c��F`u�Gc�k���q�N_ ��H����L����e �������x3��R�I�?4|�v�7(�0{�����j!�b��b\Gm��A�S���k��	X��c�~�`m똥	�)�"ɖ��~�.&\n�~���6�ZS\��n��a&~�2M�t�����7^5}���������T"�D�pv/oW����EVٱK7�����Zc(��n�i�ZG r/���D����x��gP����~�_��B��E���(,�|�m�5)��]`'W�Ig�\e���k�\��T��8}b_˼�}�v�a,n��垍t=@��t��N�.��|�z=�")^�G�%'�&.[�|8�]L	�f�ry�E���G���Q�)}(�p�$zh��W�%�^�E�ߌ-�ڠ�l"�p'�d)j�cS���8~�6��{�����{��U�V����ɋ�]iű���۾b$֝�6	P���A$L=� ���J5!��C�����:�K��K>��G2�B�%��E���]}�
�����d� ���(���/�4��夤x�
.9E�ql�c]���z�%��S\`�oIhy<�X���WE�k|�Q���vZ�%�~��_=�Fԏ���4�;�m\���8	�.ȷ�GbU�G~!� �.ߧ���$���|�#8��žk��h�su��ٳl��GI?T)�\E�J�u��7�p����w�zm��E��]�O��k�{:�R�:.+*J�
_,u��,l_2 �i�R�� !��񾿿�ږ��q����Wv�@R��4�k�������E��
�N�Q7Vn�F��v��_��O�Ƿ#+��i ���=�j`ӗ�޼4�n�nZK/�kV�3��~[vP��r���p^�/~��
5�[_i�)�i�w�g�Ѭp7�=��̙Η�u����+r�n�ڏ!֪:� 8�}`C�6�.K��$����,a�Ӱ�:�e؀�:V ��F������(>��`G�A��T�����	��҈`�\*0p^�kd=.Ǵ_[+_�,�����Mw����Q��`���Ջ�R����ԢM��"U��Ë*�޵<��
��!-f�tmP�l��.�{�.��"��؏y�O6d�8,PW����h��ᒽR�z�彁��B<U4��-�eӖ�͋K��[xM�-���ݵQ�+�/e04ѷ�P��F�����֨d�^�f��K7j���rD��uZ2�O��Q�J`�Y״'.]�L� W���a���m�x~<Gn?E�^��j&��aN�pW'Y��m�m�g?�J� ����mp�HN[�	��M����_g���kF����w��1�]���,Ƀ泐��[O%��?Mh��T>39���A�Z�E�t᭗�"݉��,�!;�����lV��Cz[�������g�\���%1P}��(�����YfH�o�9&����R� �����T��C��78�Q�Q�R�`�>�IH|�dU�e�'�����:u<JV�Y	K��<�����#��v�jUU�����_F�+��KM[.i�"��J���=�t7��ʢ�_67��d>�(������!�`��&�_Vŏ��,�I�!�.Ep��I05���$�	���U�^2l�[���2�Tǲ�B�sBu'���r͓n�_w"0�Ahj7�S��D7#�6D�yC�w Yp'����C��zeA2�A6+D���<�[ӽw�mX����I�sz�JW-N}�����}��{���/�w�w�JiOXM;��� �
��ˋv�,��ǥ<��C��mU�����9@�qt�v��=;,�և�-߹�x~YzȽ����":��|�n�؋���7��ѣGd�#)��y�����؞�	�9k2+6�Z��dQ��-\;� �N��MW�Aۛ�#Q�č�d1�[�$�H� }��mVtf���D� �e �FD'
�9-�&���6��ߵ�(<��,��m�W��9����(J
CO���D��mYg�f���.o��N�X�1����v\?��D�� � tC�}��l�@�`���:�͍�&lL�����K�:�9%t�����¨����1~N��F��4�yl�.��M!zNQ金��&Zڗ1��4ƣ	��<U�ȤA�y}1�Z,1�/���6+�k\yUXW��+9�a�K^���Rv�,L��O�� (�	�-|�a�7QbT'L�����������f�Z�l&�,q�K4r?��.ò���h���AF�N׶�7�}����۫ -�d�{���jf��H,��*L�c���y���������j9���Ά�K⚼�|Ƚ��@f��_�(��5g?+�N�
���(��Q4G@Vx���{e�!��j��:��:��{*t,`���Ъ�.M��0�9Q�!߆#��.!+��k��H��aU)�woё���n�N>� �@|�}[pT�z9FT�'��2,j����k���J�S�
�P;�f�H�����U���d5��z���*�]�Pe-n��  ?iM)�%c������C�.�8m���������ZR�G�cm�*����ݳ�?�z�ž��.�a�n����+��0�:/�l����O�����٢k..FƧ������p��-+=rH��߁�F����kB����-�AdS�ڿ��iōT�`Up�������<��w uP�A<�8^��2�`�np�f&�բ��$����R�p���_�{��)pF�h�E�4��Q���U��ٗ��k�Q'˝:��3%��Es�c�xf�i"w0z#�8xL�ik|M$�Ka�+m�G="T{����9�]8�墕#�&B���ߠ �i�+��Ê����( ���u�U��p�2�V"#S��;Pj��ʹH&�=x1\��X5v��܃iw������]���Jb�t� ��b��[��b��`~�E��F��/'){���/Tԕ���r�޻�#��Gg�C_1'���,��|3'͉�v�͸�OS0�/�of%���n�������Y$��Q��>h��6F�cY��f*X)"&�r���5�b>��������������+��P�3��Vqi�fZ��\+��r�-�5�?LN�A-�_q6S��[M��:Ff�.{�=��w�b��`F�gk4�-�\�����M�I���=����B�.��xN���26Ҽ�c��bl��!-�"C\\d�E�4]�&����C���Y��b�N��O�����U�j�t��:3�oW�1��t+!��pLvR�j�n�/�1\�3=�0T?�~b,I�h&3�f7J�z���,�!�²�ho�d{Z��0�1b�h=�T�0���D�N��N�70-�?6��R^��?P_�i�l���FQ�	q8�4ֲ����
l�l4�)�Ǹ4������[*���������+Pqsh��f�z�[� ��;YnWɆ�O��sV}Y�Ч�����/�t���o�uF�e��]��i�dM_y���apo���:٭ޒ=~5)Q͘�����p�����g�=���jw�nl4]*�"�K��1�6�3�p�؆)*φ��f�D||��lϳ�! ����cl�`��VO�G0݌�N�wm��,Rl������Q�ձ�m�����B�1=؂�L� V����	��]������;���r�F"D�$,!�o�Hc���b�'<|�o H*i��"-��� �Gu&���w0S�:篰��ˆ���j��#��_���v��X�x�/4-�V�Sg�� 5��!�7����)��K�l)E"�1���I����J\_�yn��)�e��o,��O���f�p,Pwwpr�8w��= �$b'����_�zA<\�]�'?*���,C��;���Գ>�~M�-���S�������K�������`X��cVuX���}���$5k�bĽ���X(t�?��G�(A%e�����%<�Yyl�w{�ix>�Y���W�C�S҈���!M�,�wo�(^�h)���$+��A��7�
��O�;6=�:{�B���vp��A�~h1�[�ʖ���-t ���ئ\=�3$-`Dr�e��Ǔ��s�����C�#s��4�`�jY�*�h��y��g]����kj�C��邽t$����00E� �i�LCbPf���U��{����ޕ|/�u1z�0n�N� ,<\�GZi��yXD��{��ρ�@�Ztp^�	V��Se�u�dd[`Cg����֑޽�����L
�Gެ��f�p\�������N3�e�ڂ2
��R+m(�?R�U��*�$�B(��� "�����G��}v~�p'+���f��l�X� ��r��8�4��D���	I5(��/Z����і�z*�@�Rz�@����b���9Z7�y|����2�)(�]��c�?d�ɟ��LPa4CA7���bqn�.�y���h��4�G�L�7$�y������By�s7��U�n���[��u[�?���dMd�靺�AD��.���N�N����z��tf j��o�+T
���/��iu��l�Ch �1��U��
6o�(u-���9�r�E1�'����N���c�o��QM��l�$͟ ��U�Fc\��w�0y=n����n`GR#��ǜ2w�l�hD�����p�=[].WF��.&&�l�Rڎ�q=Bl�ga�E���Tj�++���2��d����q.%<K�;|W=I�	F13�Ί����բ3aIms�&ц��27G��$Bݩ���n�q���.�'��h��Ů��և&D_��E|u�v�;Y�Ty8���tC�����H�H!��Ƿv�ʖ�zh�M�BI�J�����������f�u�[��j��ŀ�Ht�|��,�����٩m��8�����d� :�c{$�������q{$)�o� /F�5XG��K��^�x��*|R��	���bq�x؋Ct�nW��:�n�@�'�Kſ@6�#�߫�kPn��#�� ���Ë���1t(5�`�:�ӉH����K2�^�?w J߇]��5?&���H� O�4�S�LE�`��ґ��JG���_7����~��FB����Ռ�I��`אQ[� PJ�r���bV�f�e6 h@�=�'��8��*�L�8U�ӡ
�C,:Vρ
\�9��L�J �0
��M�Hi6��s{
}x<�{�j6��E+���:J��;=ȳ;�XL�sə��,n�_zЧ򥃹}m�2H T(o	�X,�5�q�\3F�i]�;>2�~�V����Ե��_Lk�9?3�x�# O����l��	_-7����z�os�<}�` 'm;(}UZ�T���<>�s���*�Rn�/����M]u'r�����&�����Ɛޢu#	�l����d��Q��r�X`#���tt�Lt�t��W�.��<X�-jsc��6cB6�*����yw�֚��J^�I*^*Ҵ����=�U���V�&%ʪ/Ƀ�vb�n�2�!�-mn�����P��v{��x�B��ޒ�V���I�_Mryǆ����-)~|d9l��y�¦��a.>/�i�56�T�;�|���Z_?<�ix�nּ�����[��g��p�D���zs�q���$ss����?��a������0�HL

+y'��Ic.��׶������VOڐ��B�m��l�\mUT�f�syig,�	0�Qg���wj��TX"�7��t]�%���\��g�T(�,�{Se%��G�*������Q@%B��RU�qCNb����򸴢�A���`�ɴ1��<Aó���K��U�d����U-HS��{ � �M/����^P����-G=�{�J�W�S�V��07���Иg�R� 8�D� ��&�m���^�ಋ��_a���4�����V?���H��˞>YL
�{��[��̆��C�N-�/�+���͖�b&���1�N Zk�ぜ@�G�����ٹh�|+ê��v��j#����w��bn1Z]�Ϝ7���^����0�!��݃�|�1ѵ%{��A�9�]8��#����V��ϛܓ% ݁�u(�D莵9(%�l�!S:�T��5=U-l����J-�=���N�����Qwدq��KИ/�*7���g�_1L�����tİ%X�v s�`?��͏��C�����2���t@�ȫ��1K�6�z<��Z^;Ʋi�+��t���=���h�g�66҈ns�o�Uy4��n�}�_�9��so�ӯE�1Ѧ`�0�!.�rQ7s6��B/�!�����c��3?FhJk#T�&P��a��k�?f��r	(�qE��>�[A�O�|������K�xl��a��N��� ̶Ag�#xL�f �TM��Fa�+�o&1�i�-xU����tu>SZq��]�i���N�r�޲y霉�~2�p��Ek��Y�A*�/S�ۃ�.����<?J�oX����C�?�,*���^q'���B
>�B���F7���$�s�͵��>/T�<��բ�<Ȭ+�y�G��誖-Gh:^����j����9!M�_2��9�Xt�sG/�9N!�s�o�&�`�"�/�@�-��t;7��_�y�b���$X�\��jǩ��}jl�s1#���VԹI����1�4���Rsq�������Zw�%��-v>���~h��/b��h���p��v*�����#���l�%A[,������sغf�[���E��3:7�A���5��;��J���Wr疩��R39���R�V }�f����zlp�����);�3�����.��Ţ_V�j8a�ԗ.��C]�D�����~dlF��S�}Q��ȯ�/�dW���/>�t_�t��4��*�\��ʹM���_<��|%#�R��L�	���"S��úIO�&@M���FL�'��=<�9U�=�0}���w����kC.���`p"������q���ʏА����/��;�9�]*� e2םx=y.�/1�c�du�vDG�ŦxQcB��稵>��9Q �G�/ �+6�SC9%>��ME,�`k�� tv��?M�蠧ݎ���B*�͙��~F~ۆK����{�t�W�����>N�3#�L=1�s�������MJ���w�s$�I�Bs3~�a��P�I�hs]����kc���6D	���Ja�Ojn�0L#��2�`p��v��)���;�a)
��N�7�5|��H������
��7�^��l������>�bN53N?w<��w�N��N��W��+6�"�J
Ks|�ԃ����cY@4L2�!�Wx�tSo�a����4:�~�n���W�Y=Qo�C5�;`>PZ�c�h�/�M������߱IkꚒi)�F�P$����{r��g���>t��NiV*��䲨'�d�:Xot0!��A 6
6M�Ff�!��m$�c-�&��kgp��ɨ=]�� 0�Oe�8T���t5�������9��캵}��k��V���D~|�kQ��)��$y�s���z㍥�?�[xK+�q�ml��m�֓�lK�X��i#BQ��ֹ-Bk���-v�[9��S� ��
)���}YC�/ǫ�srs�4�Y,���h-b�-:�۰`!^5p`��3�*4u�ONKE*�3�&���vm���X���ۉ��M�6/����� �I���p�fw�(QR���E�{g�rD?鵡r�rBߟ��V���ś�}�f(���!x^k��"�g���	�
{�L{�#���Kߒ��e�۸����윿"��� �.�(��-���p��eڵ$��t�_Ǭ2O��%��|,���r�i�gB9n�f��z�x�y�'W�*m�#�PS��J��?o�;�����&�F=3�ƹ�w�+<����Ȓ��1�?�w@EpZ�m�6��ea�����pj��*�P ]��WOi�;��K�H������kxkva��ME������G�Vw�/N��p�{��r��֯��e�gm7��kȹs����t-lP�t�pQ%���8C~�	u�b��y�6��s��]���(+W;���g��"�ѯW&�tz���F��*N��i�1�^��H-$�9��9����F1t8����%R�����!�9h��2o8���0����7�vPu���V�9�n��� SOY���Fq�"s���$�-s4���e�4g28z���o�l9�ĭ�Ȏ7�Lr�~s���zg�suZ:�U)-��2 �������yƛ��7E�њ���x�|��������i�(�H=�"J����7NY�O��o^`3�-�>R5��̑�?�K ��lyI���a[��Y7t�e�a�>�} NR��ض��EM��b�K�6��è��B'r���3�o��f?���j�������̸�9�,��c%�Q�߇��Q�Ǟ��<���A��# j�&���g�c"�������q�tt<TV��_ UJ�������ӂ� '�DM����ʟ��f����m�-6窖�0hͫ������=�c�Yأ@XH��5�ģ����%�d�R��p�h�N�j(�y�'Ϗg��T���Q�%/.3Г|16 ��3zs�=w�҂���8e�vTF2��ҙ[@���RL*�ݍ/��c�w�bpD�/tґ�=2jՋ�>AV�d�ϚԎ�	:`p���rzi��2���/&��Բ_;�i�}�|��MRW��Y�=2眇٘���Hō(fh�����\;n�i��&���N�� WwB�FX�N26�k߱h`��[=�L��X�����R��� ¿�b��ݢG�@-=B{)r��VZrD 7�:-.�]���M���d��*��o��:KJ�;-�ǲ�v��	��4cO���I���6���Ƨ��Ȭ��^yLe.���u9 Ը���e(�*#��Iv��8��l-�<]�]��.��}WW��U���R�K�m�2���1M�Eq$���?����_����H-LP�M�!�<�/߁Aa Z�?V�U�u&i[צ�={ 3"!��s��d��J-�=S�����Q<n���ϻ��`�`�(�4���X�3C(y��N$^�/)�Hn�(�d�=�̥�\�Y�:Ƙ��#R�&*����y���v�7��.0��h_�^����a�%-�W,��f��(�`���gO�-��/i�����X"BO|�_@Z��B�����ղ9FvƉ�����
��]}g�B��̮t���j?�-[��~.�!�Ļ!ъ� ̮�5`��8������xm���1��&�p~S��J��G��a��e \�a��U��T%�Ř�,�y-CX���Yn��;���50��HR��R�P���ЫV�^�����jW`�0;VNz�u)->��V�Z��FJ���^V���S��A��g0.����uZ�b����i�o%���Xr���Ħ2�����{z��&¼ҍ"�󟅲���L���҈�'}�7Y���睙֥�h���\��e�������8�wfX�Rv�'��O<��!h�-�'EEZ[Y�]GV��x�l�0ӈa˅� ��
@�_���.o�5ț�sE�f�Cn����({�U0�G1��ʗ�=#)#�Y��b�T�?Α���|��$n�w����'��źh�>L��a,zb�Urp�?�d����wD#�[��y�
������3E��D��VF>X~mg�xz4nOk1�¨�1���=�����\c��3�� �E`,�R'��F$2�ED��6L�`r���v��n�_�4+;l�Ҿk{�:O�q]�YY�$!bhbW�=�$�eG��?ސ�����cl��"^cpG�Kz.��9Bz	�.�+}Myh���+��,|u++�9��V���ہ�	�Ô!�T<�����1��ɱ�ѾK4Vb�~�DX��Ȭ�1�|�5�f�	���������:��V�U|���s1]�[�5%�m�d��6�ƶӏ$�(q�9w��f����z�ø�ęܧ�8j�����U���<m��2%���j���
�vLw���g�t3��{��J��|��6��Ց^�T��E���^�?Y���*�9r�L2�/�� T�s=U2�`�S<c�Y��>�FrZqC���*f��^��:`����nL��2.,�jn^�>:��ߞS>:�~4Ȃz���S59h��߬�C�lK؟j;(o]o�>+�HS>`sX��BJ��5��'��`N�8��Os$��w�`�dtu �.��~��y�N��D4t�Η^�d~t�>�/N��@G����>"	��?Q������0�>9���,xǭޕp"r�iI���ɻ���w�<����E|�%�a�ex�\J���D^'��x�B��7{��Ӷ]���L�^�"f�����\=t�l�n1�-��z���/��&� $�����{A˥cΆ�7K�S$�阮K��\�
��S��gbطܞv����R�uvئ��%�n`Y��U�8#C���-��u5��9f
مH	�{���O�T0Qi���0@���v��N׸��I���H}����O��y�o�c }l,v���K28ꛥ޿���ւ҆}�������\��1�@��a�{��L~;�m�j@��䕟�����s�GHh��X��ᩣi4��_1s���7P�(��d�׿r�`~���s�ė�V{����$��[79|T%�I�� �D3��/xF�`�܏i�P�Ok�fڄ��z̛O�f���OmMY��Z�`��̆���ƅ�ٓ5�FrWR���U����~�Aۃ�6�IK��4f8��b���p=��8Gj����;7ɲ'~l�f������Ɂ?�30��4=�]�3����fk�=;#�V�M��A���ݝ��C]rp�,�oޜ�h�4(�|�ɒ`�v-�����V���5�zg6��uU���:��Ú��3��	�C�'=j��!��!d�5֙�{�Ŵ�B��엦���Ԉ\������y�*�vND�'=fO/5C������C�}��Ok3f9��Yl���s5v�QV,����zC�f.����gd(���R䀅��M�a�*�X�5����d�*�ڦ�৘�#�?��`�t�bZ���fYƖ�\�}�?ڹ3<Oʅ#_h��4ͭ��;}�H$�2�� �
���W�y!�D6��#����Q�$ְ�U�Y�d�T��O��>���k�5\U�$���4�$�,[�| Iذ,�
J�&X_ � �
u���G�V�vF�u(b�����Xoʉ@]��4���Z�&ׇ�XQذc���	����E�)w�)Mya�O�Ew|_�0���³.�ā*��RǦ�J7]ڡd�i�>;S࿌��-y��*�/ȚP�	��?�5�I��_�<��ݖ�~��?��H��X��̕�����m�a뤽1���C�R�+�>:u'o?F¾n5�evD�|Xg����@���J�)��޻bw���ZC���)���,&?���ԥ�V�x��A��+���I��m��:kh�ӝ��?���ͳ�Ϥi�$����ι���AN��_�Q���s��]�%���%��)A�S�Kq@ͦ���)�B��%��o��o`���<zv�s��h������
Ȭ*�_{(rī���^��u"v���_#{�b���E�S�T��!
��b��y���7K����Ŕ�@��xu�U�+ّ�ҁ�.7�K�����Y��=)Z���A�g�����˓g"�%c�����bj�yw����	�o]�����;��n���d�6w.N���Y+gT�Ka���;d܇O�o����9�*���1�fqy,�)AD���T�c"��f�ܬ`Y쌈� G��:��ݐc�n���fJ�!1�?�U<pg����'3���b��*dCV�_���u"�}݋��q��FR�_5���)kr> �`I+~:��<���s�����l��G,��ꀣH�>�V�=SN�(R��4ˤ� �M��z�W�B�ܺ�6Yi�k�� 'V�|��˯�^��;i���Ш��1��R��^�9-��s�Cg�2d6)�.*���"�i��n���7�1�I�cp�4>���Xh�ܚV���o�4[������9�{����`�����M�\��t
V	��9)�i�g��Y�@�����8	 5Z�m�����-���4o	&�"͈�[2�[���,s���1�~�6��,����J���@��C�I�q˾xiYD�?J��B�ޓ�A.!H.eÂG��m����n@~]Da ����W�"Jj��W�N�r�G$�1îxsIU*h�p^D�^&�DNA�]�Ѫ;���'�5���Uۿ@�UC��Z�an�&��rlp�Ÿ��v��Q�c1�k�C�}e�bƶl��X��LI*N!"�ޤ�� ϡ��r��S�<���W`ޠ7 �	3�;�8Ӟ��ʂR+}X�	�4��w !�D+�������i�Tz�~+U�H�?�:#��3�
W��K��Bd���Q��+��z�Y<{�o�6J���}������&4'L�Q�ҙ~3�WΨY�����X^�e�����n1JA�<x�$�b�egU$������}�
�k� G��F㓿����NZc%�}n0 "i��[�ϲ1k�#9{
�s���F�M���P�3^�������
�!��K/��hg��'�UR�9�RӒO�%uAgO���%�/q�Q|�����!��e "�D)���%���o�Z�2��-�5���3��3_D�ʝ�u��Of$�S\��'���P��&g $�g��/=�*��������v�S�? |���Gus&�Q�>��{$��S�P��X�Td��d��Qxg���A���y��嵱�VB�,����X9F��sS�p�R�4�9�L-W��*�u�~�4I?E�@��{�^�2)���41 �� ���		M��=hE�٤z��YB��HB\)�����iT����zxhi�!e@�d	����Nuq��B��B��]W{W!�*6|��
d��r�d�d}������s(b�-��RBq�t�*� 
tV��"�;��� �VgN�w�8�L*��u�Qg@�� �g2|��Jm��k���m�ɫ�'zb�Z�V~P8����o��#D:7U�Hܹ,%3�J��H���;�Sw��A����ǩd�80m28\y��`��9�OXX�,�RNUj���9�W>~�c��'�D~��m-��o�,1�D����X@+G����ȕ�y�o|��Ų���({���k@J�DK�IR)���AC�}�P��F�W3&�8�ZEu�a��w�"�	}Vˏ44��)���r���r��F�{���ʟ�MEE-�>P6N�^�����דu�{�g\nW�Y�n/��� ~MW��3�k�Nz�K�1�{c2,3℣L�����'�!e�m \��ZX1'���Dʬ�	dc?d��a�ӯ�3�]�_�:��B8�g��y��ߘ
c�G:i�2�s��7a͉>���w|F�y(��#�Bt��tWF��K5��[|���p<B���D�"�/ɶ�Y�^�'iy�%�;���A�f�۾
�S	Z�=�~lp����W�p�hk?����������J���u�7��	nwBf�Ǵ����d�ɩ��٨�����!�(1%t���Ĕ���9���r��^]=��+���Ӳ�&U��75C���*�����ǣ���u �\�7�Y@Y�Gbs�=��ai��f�ܿ]�"�t�X*`�X|0ߒ�Z��Bj}�'n��vZ����[�,mL[�F�]�0�̆Za�%�?J�����mQz���Dc-���,��i����.��c��	�e��J^0�If��.~!�B�L��n~΂1~�[͍�XO&P;����!�O�&j0RĶ���߂�䒽���;_u�Ֆ�|4A��4��:�|-����1q�9
�q�n�CG���:��.�P��:����]T�K��.�c�W>��Z��1uQ�P��<,E���2G�bj�R�y]$�,`� ̴�*��]������Ԇ��l��a~<�s{��Ɏl`�#��O�^4�,>(F}���_�G�xS��s,�K07F�F�R=OW���؈,P>������cU��>Y���j�}�R?��N�Tr���`,��-2]j�w&|/҉��kB؝�p��������!ƺ���*m��
�)�Y�L&!�v�:�c�,��]�)��]��G%�ޝ��m���c�S���<�@b�ӿ����2��/�L�����RDuG�����;d�9�"�?5�3ǘI;˖����I�2�(>�O������>���m����:��G��UV~l���9ލ݈U�R�<�J7%�J� �r��4d��j��Ƕ���g���;������P�^|���=ZB�~ �f�Ѡ�X�|9� �2��Qh�+Y��:�+}��b���»���p�f��
��s{������=��~jս���x�������ԭ}��j��쩘��Pa��H8���w�� ���HLQ����{��o��k�g�8�ۚ�"��u��85����i�I���$�Ӟ����:���������S��hY,��ΑV^�ǐ\�tB�@ �� �&U���
v�X�f*"Ǧ�Y�ވ�$��Q��)ӝ#<�\��aP
d��V#OE���h�f��s�/�ᕯV���@����m�Ng�Z�!l���E["�S|�����1��Vs�ڤ6��4V���J�t�������0ߠ�
�+��F0�а���5n\�#k:����^i@�^Pg-o�.(��p��Z8��YkQЫ.�� �**���-"�Z�W5�i���R�ڟC��T����W��#^2:6�4�\8�Bst@q��(Q�7P�gX��D�-�2��n׽:J�Q�ƸpYn�����\������U�W��2�k�>'~���c��$3�O̩=�x��M�7/.���~GRMG>���z�pӝiz��Kϻz�y��
�K�R�x��/Fu�!�	�/�ȫo=Y���Nn���F߸�����^"��}8u��ԗ$����~��P#�PG����z��O�AN���`yT%o飏M:�r
G�t@��2fyM��K�������wT�w�w��Q�4�>��1VF��eςם�ށ�x�2��IUA�=�Fi@?�ɼ�������3h*��ׄ1h���MU~��/����*��uJ���b����`�K$�d���k���d�`�L}��tU$�ˈ:�� �v[2�?T����rQ�RN�4��lޢ3gW�u�d%;.�Iml�_(g��S5�/�b�.���!��%p�⟸�㽸�y��w�-�sB�R�f�ΟI���G�� ���%��.B�
)��1�YNA逺`�L���M�/n�~�-��4� �\nu��Mċ��_Od��6^�����(�BVb� ��>ס;�d�:٭�Ҷ��kY�:�\<'��O�1���ދ&-,GH��^�R�lQ���Q�k�]�@��Y{�/�|c��lt��	g�t��{��9�����q�Қ��X���v�R�,0��D{XƳ+զjZ���t��l�DYn4��RM���]�w|@��Am��נ=uD�vc�\]�6�^�|�m�Q��m�m7c��O\Q���C�T!�0Q�j�kl����}�b#������B��ߎ�����H/$�qh�['�w�K��M�o�Ȫ��1�ԊI�QK\�׾���y�sh�(�0��Hp�5W��E��l,|uّ�ng��`��u��p�nP6�~�!����S�?�,_��x��,��e�m�]^�S�q�
�rjK�<��Xt�n��`����
�v2.%-�=0=����YP�U-{)Q�Q�AfN`�)q%�NǙ��ni���y(W��P���nhX�w��h}�<|;`dr�/@��������ֈ���|���q��uf�U�:Ƿ��4�I�u����<k�G�f��[�Q<�#�q�2���ăɐ؅�k%v-x�<�?B��9�7 doj����[`����O
�*�A��F��>�Y�VB�s������c�{GU*�k�$�.|>�;rW��v�@(��ˀ��W;�qoMwT�zy���1��~�����gz����c+#<
���vu� vs��׻C�m�}ŋ�[�[�`���|�FvJ��Y�k��6+�Y-��,N�,��jl�x}���+��~L��[���a��r�/�mW-5sT��RPp:�"����!B����u��T�Q�h�w�>�����*pM�K���G�b#�g�M��d�\�P$#�J��h=o���Q	�%�j����-Bs�5�2�m�[ˢ�1��
K)����RFL���4�u��?v` ���.��>�q���m}��r�q�`�d��6J�<GJB�y����4�s���϶�=�o�$��@N��+��O��|I�������%�
�2&�� R34���z��S2���0I$U$�l��ٵ��]��?���.�b}���9���ئ4n�:��>�=���cFm�g4j�[Y.j��ɘ�����M����\q'�I��鑡�QK�Q�`����.T�lHYw��򜱂�&�p�7�~A*�_�^<���<y�G�؎,������F3�V�D�Ln�ᎎ�5-dgр��/|��y�P)�tӷ��߉Yd��G��?�Ʈ0�. WZu�/��ۺ�{���:���!"�0��.8aA5�|*?�ټ�Ĉ)�N;�Ҁ�
�l��,c-��.����R�W�Np�{�sڿN����&@)��ԛԺqGh���յ��i���-j<��<:N	r[�RH�^!���6P`a�4����@�/%	6��@&]�e��p�ގ�X=_����-��@��/�[�����Ҿ�����C�p�s|^Tu�Sz���4�i�B�7�&���Px+��J�6�� &Ek���s�������C��W%�� �@l�eժ��n���V�Z�6�1y�$C�?��c�7�j|z���Y���/�_�9�F�k�71����������Jq43���DK��������!	�ͩ+�xAcr����Ý����ʹI� ?�vm��K*�-���c�Ě��B~���]|��˳�D���z�]�lC���Z�?	� 3��e��6[��3i��/ר[�m��6I�V:	L���%_8�9k��3Z0�ntG�=�y�9ͅ�j��* �iҠh�E8��_{t�x�����q#���)����pC/���P:I�rv�+����h�������&64}P�V��U�
���a�?E�2`�'��%Ʃ�T�$�2I��䰦IL���2�Ty=���k��)Fk�3c��Q�w�g��c��є���f�0g XC5^ڝº7�ư��������3Oy7��E7�RU���w}�OpVc�ИsU?~���[k~uJ:��X�_g����F\�y��1��Da���c>�J9xƎɟ6��WQ$�%��.h�s��1y��������;��*�ұ��C�UF홶������Cb�zz(�o��+���TVB	�I[��K���E�"��/��M���1r��Qݎ�Q�0A�5>��q{�K˴�`~�W��*f�?`�[vF?�OY�뜵�����B�z���c���-<z/�	9r❘�K�-��@�u��ᾘ��/\?Q�D/�$KT�{��i��_��a.�{(��r8�����ۥ���z�y�;tó��䟁�w5�!	Q{�s�N�x=�Y)� 4m�˓��̩��ݶP������@����<��-9�Z�p�-�����=noګ�x�`R ����	�UE���(�H{��|rдN�muYi���p�{{��$��îDTc_���3���9�_PȆ�<�{�Ǐ�����#CT�ə ��|\A��B�M�}5�b#Av�� 	�S���6n#���n�U5i���eW;`5{#A�*��O��c�&�96�mӹB�7�h�!�"�I�˸!I`���6�79�rA��j�s�^$�ظ,eW���19��� '��������j���AN>��r�aV��Ċ,}���u��U��$.��ptNS!�b�:��(��1�Nu�c�#��27f|�*�T�᪄԰��M��V8���O���5uhSoQ��Z/��	�ˢ��ŴG?�&9阐�����~UJ@��� �j"M;f��&�U7,U�[�����	&�{���μ4u@�^{s�h�{n)��c$VF\^��DI?�b��6��T8.����E%f���ҝ��4C��M�F��5�nt���{�����d��ְ�j���2��1�$���(�k"�,Y:r �!R�X�)?8A��XMD���s��1I��P�����G���B�a/ ��]1��,@B���@�l�&���-wAjߍT8�P�$�HzM���R����0���k�q�<�L��-�v,Y6�*���	�X�~��x\��H���X������� `'~b��й���dyd�{������w��-��)�1d���
�Z�%1����\�H�(�!*���R�K�q#VpH+a$���rAej喱!��hT����\k�;������t�i��75fiӄ�����	-аJ�]��^{�q��H%*��R7	s���A� `�^�.aO�إk��T��M뢮���`�~�Ъ(U^����n��s���dj��sg��+u���p�5DomNͿTZ�v�'�N�FS�-;(P~қ�\�â�uzU��Ee+pt��:�
{4V<ia�rdf�쾞e�|ӗL���"�<�iT�	rەb!� x��O�YNBr*k5)d�t9Ү�2/��vcܸ���f`E{*�29H��8���8�
��.oa�W�<1=�B��G ��Go����*����5�Ie�.�]���J���\Ht{nsV)����DS�`�y�Q�N��=������D4�F^9���#����xq��/g؉�s��*�T�7˄2�A�o�I��+,�)iݿ|�!a�J�����mghm�b�:�6��p���^сg"����6��O6AH�[�[Q;[�l&�h����F�>�)�/}��e�[�c�+���B�$��_���2p�{O��q
�����8p(�	�au��4-L�;�U~}q�,�Z`����8����E�2ɯ:c��+$@�-P�/�EP޺��N�@���P�+�퓐���8xp�4&�B¯�O�D9����^1�	;TJar���tN�W���.�j����;I�D�w�)��]�G�x*�nfH�+����P�����ˠ��� [1y) �q˸G��� �<��j)�dFB�B6�/p�f_��}�q�.��Es)�Ns�*��.7�$v��0�������Ϝ^Ym����:;�5#�;'�1%	������;�F*Z� +P��.�l�($,��������7�Ҵ����9������ǧA�+<�z�aߴ��Ē���r��GɡH�H23���ҖX��{�L�Y�v!G����\|K��.x.�|D�t���,�C����^O%�������y��שּׁ�MY@!�f�M�!B�_O۴2��>�!	{��Z�%�j%��Q�_������;�p�L�]�c)����rH�7Ϛ	��eb�ù��T��j�5%�iV������(���EVv�J6�w���zd7�`X0�GY2�J��v�-(�tC���;���-bA_�6��-���$ؙ6�a󄻦eH�D�f=#��b6W)b�{�FY�p2rǝ3�o<�k�'�"����eCc�ѪdF,d�G����_S��W���#�2����[R%��.��}4	�f��?O,�'u�µ��<v��V���>E�2E��둥˪52��νF]�<_�J�!����C�<��*:��R��Hp4�|��yf���1���$9���_��h�:���&�K����PR��/U��ֺ�[�����Yղ�A_��.+��eR��� �S�D6g�;2hU�O�6D��iPl�����o�wS'=p�7�F����k�8���>WnGʛ3���� ����v�ò�[����̱\�m��S �����$��b�)TB�v�7�������|�8��K�Z������Xr�ɑ7�-P��wͨ@e0|H,&�h��`"�OA�, (��|���u�k�5�J�~��OF�E�,�� a��Y�����,�'��y7�/���*�`�a�3}V��ġ�Ŏ��]�sm��]D��+���Rnn�hۓb���q�γ�Es��Җ����l���ْ�y;�׀�^"���(	$�ʹ�kR^�ZǧU�!{���u����R���X���G���ˮ\�S/�%:E�&^�O�nW��0mk-���O94;�;Dn5�nn��w��'􌴭3�'��l|%$�u��/�G������̹����?
SvY@ "I"a"� C����E���{��@���I�~���q��p���N��&"��#s�0g��YKd�A ����_�C
O�n	(i�Wql�����J2V�'��me�b(�o�±>e�p�Z"J�>��S�clZ� %JӘ�X�a���4b7���"�7�#��<Bs��:���҆��ar�r�^����Qt;Rs�"\V6?����*m�[�W;B?#E��n�7F�ŬɎм��]k���A�TND�D*3k�:��i�<=�gqb��j���]��'Ԕ�bl�ȇ�H&�ǜ��P'!�<��T�j>߶ĴŨ�
g���xP+Y �k�f�%�I3����/C(6+^U}T�B���
����x�hT�f=h����8�cyf\2�`�*��M�Wؚa��!���Ã��rz���
i�6�.�u�MW)��zCƫ�W���w����-!��p�Վ\�Z�8�Տ�f���;/��)_l,����O'�3WÐۿ��U����,B���0��;�Bw�!���1�m�:5;"G�Y�x�#��FLׅPc��6���pSCNش�����^:=���t��uW��.���BD�S�&��u��vk��C.\I,N	n�|�j-������t}�r�� ?���)%�:Vb*���~�J�>�%�&�4��ZN����ȑ�(�A��<pȌ0�y��X`�^�m���i-k�!�ګ~��(w��R
�IV�vA��Q��%��g�"���Wܬ	��2�9�)zGIqª��m��eq�
[��Qͻ����n�/���R�D, 1�Z�C2Թ(UD�稝A��;9����7�s�%*	h:p���136��n���z+�@_��6��C���0ۨ|��x"_A�����B���2s(i��C��RB�(�`��I^� "��Mz������s�X��טOM�0��o��5���x�̲'�v%��Y�������6A����oDJ'��S�A��q�&���.ZO
��}9bIt5"����ߋ�y4��l�����r(�|��P�M.-�<�ȭ�n35f�
A
l?��T15�>�K �m� �/��J�L�
.�ż�χ�B�~mx��'�dp /3� HT9E����8��l�t]��ʞ��}$�U�4��AM��������;�AY�b.�27p�G�V��^��鋦��rL�dqʑ'{8���\wf���s���쾪+~@�]Rv���Z;f�03�����}��`i��	;�)0�F	�3�t%����z1��M�mI�
tg;$ߎ-�t���m��g��E.o{2���jv��M�)�����v�*� ��
됀B��_���e��܁f�S��⏺��_zi[�%�k"���3j���/O�j'|�z6�/p8������S�}��dpͿ���f�>� ��/qx��y}�s���6��5"9Ju6���f�8�o!�c�Ѻ�G�ސ⤬ ����z�gͪ�S\B��%5s1�q�dQ�ľ!cx�{�G�<̂�(OT0y�?Z8;����{���X�`P<��-0��@���d��^�������Ӏ_c�r�k�1H~���%���M��f7�\*e���R���[tlӖ����s�Fc���se1�v@�!��� wy[p�zt�8wc��,�!%�7ߩm�FC����v�EOq�������g�����w��i���|��gZ����s2ӥ�vP�����t��*�	�a�{��̇<"����F�9�${5����O�.�*)}q�RՐ��Mrk�@�a�,��?�(��
I$[�I��Ry%W��6��a=�ݳI�p盃��|��b����qN~D�̕1ִ]y�
S>�#E6ȭˈ7ޙq}���	 �mL�U>x\mjU�}Գ�ш����t���M�Ȥ<��iJ��ū+���W��G5��r9�V�O��b^\�D�� �:�s��Q6��dt�R��y��K�M�Ƹt0�kj��4Y�P/{{��rP�a\�D3���y�Dlc ��ϯ�.���L��᫓"z���S|J�X�YF�1�1K|��$C�v�%X1�Oe��{#+�5p,9%ꢇj�>�9�*Y��w����f�k����x�Y�8{u��o����&��������[eS�a��F�1���71>�؀0�5�T1!��4�k2p[���(�r�e�z8��^�m�Z�ĒQ,�cx��c��Qi�.�Kq%��|�r�O�Z��Ov�N�[�5'���]=���PZ��=m�f��k���Ѫ�\��XǖDZ���"�!k���X��X�X���2�e�餟"<��t�3�J��kfҎ��x��ķ��wҊO�:k@��[!'P���k���Iqk5÷�)�+B���_r�N&dNT��\��#��S��3	G�=�;y�-6���ua
\��E��������l.��H�6��;�F{�K)��4P\�B�{�V�\��yvK�)��n�0�m�O绡���k��Ei���+��$�\�(����8�>��čdP�����2A
��2)jp�Ew����ۄt?:4c��1f��J���L�J"���7gv`�QlwwP�6Sj�78@9E!hc��I�wf��r	�uL�i�l�-��q��i1�<�d�?�h�ڼ�{�7�����G��L	���,�*��C��,�Ŋ3���9���b�.� ��P�5��T��mp���V���a������6����4�J�yy�K���eZ�cnLV.�E(���`{���\<{'Ø��#X�{�7�g�=�)��t�xn]�2}����>��z�^@�,L��Z�6?B�l�	OE�wH�Nh"O�Є8�X��ZF��ȭS�, ��1ֆ8������O��9hl�Dh�>vx=±-��ǳ%��6���m ��9q{��%���Z�RD�����)i4�1Pk{��i�:��\���[nM�̆ �b���}��"�C8R0"A�g��#h��R�/��dVO�Q�q�wi���W�#DH����\ ��ؠJ�PŁ�āޛ	��bh
F�/u���@ۥ0B;�ٝb�z5�(k�j'7"aC�@������ ��u�m���/��3��
�UQh~������ʍlj��rR��uA�C+�
�0��j`n�C-W�iT��V��ڂ�
��-�,^���xE���~�F�w��)�D�y;���3:V�����L�����̟��?�j������Y���<ڞ�,"�� ��3�ӽ�y�ʮDɋ����` :R����mB=B � ��N�m.� ��W�٨g��Q��ٞ��S��]�|����cP-��]�9���b��|x�m���?�s���72�n���D�8T��u��tZ|�b�g	�0�	��I\��
�V�?�>�?* `I�8�4nT�zДpS�1��R�K�dU���K�s��av������T�j�'�	�Î<��ـ>6x����B�|�,:U�N�V����ǐP��|�I�n�P�q�eTd��q$�%������2�D�yl{.ϰ�`L2�H{��.;O�@϶��ۀ�Dd�8��'G����c�-�$�y1H�����^�m4�w����}2��VC���~*w���,�B&:L�|�Q� u��Wl�Q?�$"� ��Q!���?���+�r@�[S]�zI!%UN�i��o�_����g�ӟ܊���
������q>̶�XZ1}����zk�"� �{:����6aU�ԣ�a��x�ɯ�w�< ���gi8�DOj^�c&S�Ԉ=�E<�fa:Zj�M}r�PnF������U?{��D%jo���~U)B�{��	 �Hj�����fbec����֞�N�d���{��-A~�
�]�A��I��@Z)%}���������á�l���*�{�?pH W�jj�,8"ȏ�K�ℽЧ#T%Ǽ��%��H��i�������E���6�|�oeФ�L���m�p�����������Ƈ9�g(��;��b�5����	�$������
�a�]8H��wxy�:��f�#����?�ke�f/`�G��
 w洪ݑ���:���0+�aب���D�4��2CY�4�p����[��Hy�`�W����^<纩	,�Ͷf�DU�r��M�l���Y�y1.�G�<~�Ħ���~٨|�0��_���Bַo�^Dd�g��{*[!����K��`O9A����H�w���U��!NOV[m!�*��C߰�J�m�kN�mm�$��2V[����.6�G��d�[�0s�A����O}x�����?��A���&�CIR�����?\	��oV������v���?��ta�K1fa�Du ����v��2�0��Ҥҋ�܂�ٍrh�8�s�2�6up�f:b�#uo?,H�����fΙcZ����9bc�m f߁�����ɖ�������/��� 9���L�ONa�o�I����XP���'��㲦��}H�a1�x��}����(��$��"�p�RY�]#�鞡r��{��i;��'�		��*�i>3S��ޙ
�����a��R��[_	�6a��j��#=u��-�2b�|��d�*0.6<��XIv�ȣW����t�����lI�!J|��!�=����(-��+X��zH�a6����$�jF�����29�W��R���>�!�>�eD���I�� �UO��'ޙ�O�S�H�)5�y�k�~cr��
-���{�xiMvĀކLvS��K��� ���a�j��Rj:���
W�U��0}��)���>L"^&Bq���`K݇��Â��PsW ����yD�e}	ٕ�)	oPz�˿nѯY7K�§o�� ���b�_� ��,���Fy���R~����2���"M�Y�v���$
�Eg����	�Mx�a�E�^9�7E�⎳u�'��1�s������ɏT����o�ƛ���V���f��y<�^~ ���Р�'"Ggka��~orr�@��[�Χ�e2���Ǧ�����?�aO�-�(��NsP-���c��~ȿL$�0�]��_�`��@d0��C��o�������r6m4P�ws���^n��4CP�����%�� wL�9B���C䬃`���;��a�	e��0�\.Z�1Z�#��`�R ���bA7���`�}R.^VF��ʶkI��3"�
	��(-^��v��)̇r��%y��g�趦��8���;�����}8�,4����T]7�x�|��d.7|�3͉�nE�G��%�.x���'�}�֑iA��{%3(Q����t�q�M��)v�%���(�je�u8��g�::?�e�4PbO7V{�;���*����.�(,rJ��W���Jc�8�G��ּ�V��M����r�X�x<�VRGD>H:�I��~ �I\��A���*�|��+�!+�����8Z��[$�6@G��ψ�q����8R� 8m�σֆD	�ķF��6�W&� �S�+�����"�;E%�9���c9�U�h�*��!A;�_�3�ly��Ϻn]����dY;��y펟�	t'&��f^x�N�ղd��� ��ebES 32������W&+L;&����s� �V~_��	�k��]�H�㶎��H\P���,'�{�%�x�|"��E������@���c�r�;?ʾu���ǿ�u��rb� ���ڗ��?�B���X�g&��,nk� ��0r��~Y6j�]��[��༃w�j���5�h���4�l��o̼����0��C��I��y�'0���	v&�����tR���@)�t׶����U��H;=<��̡C�;��(�	�]^��ǈ�s�0pc�
�8�G��=h{/�ZzW�b�Ih�b�C��)�~�hu8�"�u%���Z8�Wu��d.J$��R��W9%J�i�h������=�:���"!�mSI�M"��?yZхnf/�MDӏ���6�II�).�:�h�܅F_Q�+��41Z�^��x~�:b#�$���ٱm�@
;g'^��L�AI��.5�19*<\D@�9���d�T��|֯MD?Kq:E՝!����ks�"�E�!!,�Ll��!x'8���ԛ3@�թT�����,��u}����'܎�V$�3'9�Ztx�����!�6ow�$�� ������Y��b���P����/���fg�H���}��)��Q`�V�	O�nZ��ǡ��'HC��Pţ��s>V8';unj�F�O�/��ovW�1�X��#�^BBS�*(��'��>��U f@��s����H.��J��<��S u�C��x�Q0e��z��Jc��h�E�u��ͫ~�����+���^�h ��d��Hȫ����+[J�����I]���=�`=_Y�Z�nv��ӯ�������)�V���O;i8CyǞ�<���B�=�q��ɥ�ɭk��$c)<�8����8�b��'Z�89k{�����*��y�Õ�z�[Q5+R%\Q��tG��W�(7�U�<a���Jk�N�
>�d�/�ir���H�Z�>TQ���ؿ�:�C`A�knR�s(���9��&r֏FWB-U��Dy{�n���e;�X�U� ᪴�:-G\e<�¡[�7bY۱�y�%v��� jMpamxdN�At��&����9�Qu5`�%�|+��8�]$���af�4Lb8���R=@��6p��ʟ%��љ�a��� ^$��4f(�!�@Ņ5�M�ߘ���s#Wa�0�h�w �#�������w��z�>��_֫Q�tdW���#��(�8:x��O�,�����r�u���Ev�,�g�K^CA5�����S��ꐿSo0<^d�B�#M�+(bh���A��\?���n#UTb�.i�\\����X��+=��b�Jq��:�ŝ-{���ޕ`~���iؘ���\NI �hV�Zo�Q��6�l��wU���sH��$����k-�A �з���#���o�Y�SY�M7���ܔ�Y���d�C�34J�-w29��L�&�e��#�<V�4���A��Kn�t%X*�߭ˢd���y�"eՠ.�}'�4���
���y%�pM��`��Ih��.ޫn�����{6�t���Ѵ��+��o-�{!�� '���.Q�p'���Q�f�[-�>���c�f������'Y�@IJw��Q �rG�:<P����ŝ�X����#�`3�A1�s�'�t���v'�*�)���oB�����	C*��\���'>��_/���G�A���	��Q�v��a�J-j
�8����lp�<���k�s��X�?���o�j�l��ձuՂ�c�H����O�g�m� 2��>���+�!��~�%��y/�U~���*��u��q�}�D}�ͫS�n�	��e���F'�~��M� P��xO�B�d7c;��������_��L�����ϊ\Cᙲ���d�1y�Tm��%Ԍ��	fP��(x�pcJ�g�_������iqe^8C!��,{���^	�7RK��>�����{�s�ZpFI�˩7���i�c����N�E���;���2�5�Od3���';%V�Ep�M��eu�S���մ;2����b]6[��*��QX� �.&r�{@E�P6��^��!��1�S�fD�d���� ��(U��`D����J��������/��O �y��P7�����ԇƾe�S��D"F(��gkR�΍ga��ꦤ荠<������jfd���l]���0k� �W�m����u���km�A�a̥UA��F_Á�L�G�Fѿ��S���r�,�Ùxr�A�z8�C`X}a=��>az�ތ����Mx�ND�+��T�Ns�$��;����� �B��D���u�-������O�]vPN{�Y�kB!� ��N,o�g���b��'�q�м�'�@�A25y="�e�H �}]�g�6]BP��[Im���ee�$�x٘6j��ߟ�"�ݽ���r���(-=�rZ�ٝ������R�B{�zq�'k�Jr��(l�nؗ�E�ϙt7�+=��n���cY�i֮�R��H����&lH�T�㻎�7CZ=����UJ��Ge�rTׅ-��5�f����Z��ՠ<�ET���,���wKL��nJ�6�O��9}�M��J�T��9�����m��BY
S"�>1v�����ʀ's���e�x&�u=��F|���{�`�V{{��@������;-��x�Q����6ؤ)|�Xe�#�#�ß!V���_��kE��g
����8h6����.[����=��Ĩ�w��Fb�<	~���V`��X2u��W�kY�M�S��W����e�'I�$�� ��L뤆���c�G+�U�MB-M�>�6Vn�(4vi�C�8V]!���8�W�Q� _�K'��}V贫nm����D�[7�i)k4����{HS�ÙB���V���Y���;͂l�X��,�����>L|��,�N���ߥ�dv��r���V7�b�F�|�׍�i���C�9 ���BJI��!���ǹ�jF]�J��7��yۗ�f���Δ��ŌzIm�7t��=� ���t�wY��ʺx�;^�ڮ���#YV��]�?�ՙ�������n�~@���7�qa�;��`,��Us�_i�����֏�J7�JurS�r1B��!�L�ݕ�4��������G���!�}pv1?4��yXh��-�dZ�5�QR��	�1�z`�� �X:���Y���=�̞�У|v�E��<\�����֦�x�	��W9��}׽�ԧe�8,Z>p��Ҳ�o�O�Up������aY����j�ۙ����q/ԩN��z�`���=X�&J�2ۭw$�3*�g�P��#o�z�p- 0���3��!0|�xP�*�jD��gbZ���N�{s_�7��O2�z�/�6�gc�}0�����Iؒl:�t�h2��=!e����[h��o����^q�/�	`��D��W�RZ���̳i�$7����\��a(�)��֖�F��y_>��u��4TCHW?g.<��	9��A��7&������Z�>������5Y(���t:�#�i��N��_�.w�b�����R�O�`JZ���B�����P�(�)"�W�ZPï��?46�N��}ւ)�:�:�p����h �� �\�/���T�#�������U�) ]�X����������L��{�ZcrG�~<���Yr.�B~�y�s#�D�XC�#
��uQ`�/9��V�&B��|UD':�[X��}^��钛�7Se��N�uf�$����ܝY�9��q��*���'��oW���f�{�|�5Bm�&oy��5��l1���%5�����H̱z����`�c��%ntEȅ��5��v�ch"4>W����
3BS�ڦ�eVx�Iv繍�O����L_}e7�_q/W���q�������%W�(���8')9(��J�h�!�=B��H��+\�H�f# Q����0P�h~�J�?�b�aCca�* ���/�@����yX�m���z��]R�P.��]�pȘ*��0���&���r�ˎe�|�f%tW�d�Ϧz�FEb�6a����ѵ��X��2��/z��Sη�s�v�@�q|�����n5��T�6���rN�bߞ-w�������W�ȣ��ǀ;Ԉ03pP;��_t������qS�����y�m�?S�*ܝB�X�1n^���B��"�W2É��c沢��%�C�$�$���Y3�$������n[��Q?ĭ�
��}�$�p?hk�l������H�z�}S��������z�֭i��IK� ��g��.w�83�� 8c�x�w4�uQo�j�vSb�#>% bع���w�۬���)G!�����򗹀�ز��@�H2w6ȩ;A�E[�"��>|X�u;�{�k�ji̋.g?_��_(r�d�~�"�'}��94Q�=&؎���l�0 ۱x�=?�s���?�n���:��H�2��b�B���~m_�����������OFҘ8�◡�g78��}Y/�aa:sIk���09*��d1FRbO�����	kk�������XhR9��F³q����v���(����(�|����2L�߉ǃ�M�v������������M�n0U���B�%ScN���#ҧ�ݮ�&���&%5���aD�a6�=�܁͕@.�u�_[�y�x����ƀ[^�}U��DVڍ�;R�E�cy��>�њ!Q�,�QgiF��zS�)��wl�0���d��.�+�P#�gKz��S�<Iu���̺�n��	ʱ�ܳ{�;^�� �3�M�	_�p'�,׽�:a�3�V��ot�4��sk��G�R�9s�I�b��s�:	.V
�E��ATs���"���1�ٳ�g,"H����;�t���5)�	�ˑ�T)�gXM�lU���k^.�̾���e�L����>A���ّO�0��b[�x~H���!���m��H]Ϣ�WM��Gз��d�I�(iгhhDO؎�� ��Y�^�ߐ@��U�hס�}&�~Ѽ ׬�̐t�$�hynڍs������bZ<Z}��	;;%}����1��bhĂ
xQk�S�5�<�I��q1َ�bx�K�b=���RB�╘{����Uu#E%f��UnK�7������j�����Dzg�?z���L�����mN]:�֕_Z<��:�`M�ؐߗ�������@*G>��B>������ı:�iNQm�h0v֠��[m��Y>?�L1d�[ά�e�}�)�m�hT��ٙ�Zx-�>����Z���/5�-���@k=������O=��d����=��Wt\2����ǧ�ƣ��.Z���Pp�yDP�"1�Z3@=�����~w31˛"� �S��äTDo;�D奍����;����J~���yЅ)|���ԕu�&�UD��2�HR��y��eR4��V������8 <���R���Bq���m`�>��2�燼��GiC�4%��}3೑e����כ������Y3���&���_=6ۋ�)�PK��LcȂxQ|���u�j`T���͏n��1�����x����}��4�vFu�~Bm��>?5z���ΘiFa�A,^���*��1�h�~�z%��%�I5@A��ߒ؁2^b$pQ�Y3���O$Y�XWT��>��}�g;#նK�9��X��/�
��tp��(!D�ܠ��� �����y�+^�_9�<˭T�a&[?��s��w�r��nQ\��C�Pw�!��#E�a@�bض��e�kX���^�W�dL=ȥT�$����Ұs����H?dL	q~�2�(��ߓ7$ܩ�Ve����9�EPv	�l�G3��Mߐ�b^[]4}��&�����W�)z��P��	Z�¡>��a���r��S�Z�~i�a3ڸ&�̅�+ڡt���@�Ε�.r
a~��[ ���_�W��9�VF��W�a?��'큃V�(��w��[�T�?c����EJM�xAV�|l_wOk��B@@��=֗
'��c)1Y����bTR�`���@�8L���?�>P�BvE�>���$��֗cw���2���:��'� �f�7��ŚSm�`���_��oSq�v��[��MP�.�S��2��8����d�:S9J��m"����!q�)���؇���vy�f�)}ƒ�_o�R����Z�"m����y�࿚oQC=&lo�ͤt:���d����|��q���#�Z�6א�4�9܎V����|�nr�4�1���-���IP.�z���N��{��aGҤ�A���:������)�K��n�U5"�A�@����y��q�r�ey��ٚE6wR�3L��BH�m���2�!�C���g*e�F�8�<�p�͊؁=��`�� G^�B�:u�|7�#��ڟ�S��(�a���]�5�j&;��g��4s�w��	6 ��c�V�w t[l����';���!��d*��❩�#�j��k���ĵ�<�Ԛgh�>�f}��j���k�8����a!1�w,�:��!?��yA��'5)�U�f��X��۱?��kE7|0k�-WF�,4�ZT�Xs!m������f�}�Kj�q[�PVP ��È\�}[+DG��0`b��ҧ EF!	�sŪ1��8��J&�O8�E'n��;ʐ洘��sV�S.��=pi���P��$���^��n�4�r@_UE���H#g��j�,65��T�E.9ʏc�Y�j��#85�k��XQ^�t�Bx��JjZ.Otq�畲9[;ns-'6b���GB�B�_�����n�d�_ޘ����x��g/����Cy](>�1oF�/���+k9N��|5i
�G�'n�/'��W�h[ĝ��q�&���x���7#�`m�R�;�C]�`�N1z:f5��A������_K����˄�g�@vV��(�O�?��ơ��\7�i�i�F���H�2��S��0�I����ܯgY��Ee3��r.ɉ�%���L&[���T�Q��w�g��]���UҺ!}:o:kҡ.����#h��E��*�M��]����-!k):�#G���jd�q�j�L��w	��IF�z���*D��z�TI�ޥ9X��;?&���Rϴ��/�@'�	:����q���ջ�i�#�Cα�?ϋ	����� F�w\e:N���r�O�����jt�Y�U=���y�
���E�@��F8Z�ۺ���������6�E�����y�D�!X�M����2�'b����E���-���1�o�{�$�H���}'��-��qa{֐���KQ�y�l�+���G,7	���X�L8e��橂��J�PD&�IB �@�;�)^�v��t�yG����c>���֠�����_r2��׾]��3"Mߌ��r;*=/�������g����T��D�f���!�WctŠ)�S���iW�o9�b�Ե\���vh9��s�JY���1�c�窣��w���VF�^e"�H�x ��r`�d/@�o�4-a2���7zd��w#�,�z��J��o|%S.8���T�l�2�N�8#��3�汔-PR��S{�ISJ���!DHVш�X�eY�4��! DM���Vg\ef�����~]kW�	8���(idj�-���
彚�ps��!��q�ELn�^�ތ{*��Zޙ�f�z����ߵ�:.��$��� ��tX'�C��a�޻cGm��2�T3�������o���N9��	h �ptB]�S�A�3M3Yh�h&��Dm����miE	�P�����zj�8A��q���;�|2��C
���PQ��ھG�[KѺ>GD�+"�9S���4KL.+��A���5cR���R�w� �N nP��	��I���P�4w��>���ٙ���9o'<Q��9?����{�q<_<��@v]�8d��љ�7�g��$����e��`%֩XYլ�[�[����8�,���fH�
L�q���g�&]W�9 #]�IR�����8��xز0��*�
����|L���1ߥ��9�(D��/ax٬\x�<��N^�b�i'����ʔ^����t�p���+�x�{q�j(��R�@p� �
T5]�mE���߇���-֬'ֿL���0���f��C���a��>�vh2\f���8.`4RmG~?}���b�
�#^��
� ���l�cy|^�a3��v���(�U�R��>Q��+�y��t�`����������2�z2�K��C��E,�����
�]��e���P5�Q*�ηD��h`��ՙݯ_���yqGJ{v���q����iEp��wM*%=��S�G����.۳H`_��څl�+ZL���s a��p:�kНg:6������V�T���L�Z�k���I�"X~dqUaM���b��~�;P��BH4G������t��m �؏U�Bf�8]�2���7�sk(�KJn�@�#g1쫂5c]_��'_|b�	U�1�	�y�tK�h{���-LPx�-3��p�S�֞���H(��[�溂�VdRo�����@�0Np'�b�$�6$�2���u��u�_�_Mz�`� :4�٦�,�I�R�T��]hĴt�b�nf�@���[�����}���|���}�7��E| 5$������=�iҀ4wP��Z�s��F�ŮTvh�HGK�߻Ll�&�R(�C^�ڣ�����1xVX��������O�K�]�m�	
>�AT:�%�'��˜�n��z�4��k4`��,���u��)�i��xkO�Th�uiE�Z n�/��lJ^ɂk�e�O����5wڣ��4���I��A���h;g��w�p3)�O��[�jM����,=�SV]�-�x��yJ)6�'E���A�����4����L��|� �	.��0�Eŕ��! �$S�M���]3�5<KΊJ�U�Y��(}_.�?==��ǖO���u�%���T,��G��<H�D��15����f�g���G��Vz�G#t���㶸烐$�}`�i���h���#A��
v~c��ځ7 �4.sz��Ni�Ԩ{�^����L�"�����r�%5(��;5 ��in��Rت2����.Sk� r k���e�-�Qb�X6�/��h��{M��ܕnH��V
=��H%*��xi��}�>F�0I*)�;Mx�P_T��N*@�t��~�|�$J�\f��?ό��)̇p�
�sŊKsp^�'L���֠R�xt������L�����$�)`�\��F�PK���Go�t��&��~ J�(v��h� �P2l��a�����5��y���H�����C:*�2fT�&�ؘm�x���5�0*���u�v W��ćG��H6���_ͥ<��<��;����N�<,"rު�v��.X�췁���3Րm�����+��$��K�@�*w�.3�K���$�ҨrhY����N����|�
���u&�[������z�l!�e�H��(�kA�٪X�*��Us鍑b./㍧�]/�4p�X	[X�Q�}�A��)�`��ѥu�.C:�i:qKFQ���i�<��-UL����=ςPAT$оz��}��W��t�P�~jp��c�MO%��U�1a��@#k������!gN.�}�?	BP1�*��_����п=j-T�<��b)]�3�^`͝/��c�~�ۢ�ܟE#a�-lg�Ե��0��)�iٯ���j��2�31����UH������/�m-�4!�C<�N���2�v�j�<:�DR�7��
_L�#V��IO�,�[�&��
ogq��p�����M�|`��@�'`(�۠�@�0���QZ"�s~�L��(Kva>�[��)W|&\�E~tl��3��Ħ�^|��r�*&��|�������X2��!�����V@���<�'	�J�e�M5;f����,h$�m~�F�.�|y��a��~�4F�?�5(���+��ne[�C�Y
�5��jǡɴ��R��ëw'����
����|8�o��Vc��獦����7��������������XdU�ʧ�� 7�܈���)|�}j{��y��Y��t�a>��=��j�T�=L��N��x��ݙ�,�~�/����q�x��]r����5B�B���h��,�Z�2���6���uԜY��1�J,ơ�r��&>�_�"r'� k퍧�5TneN�{5�H鰡���K�;�u�/�6>�D_jG��J;������h� e��BpަxN�i�'z-?��G)��?�XM���2X�D��چ9x��hF��Sc(yƦ�!��O���9�~n�3���W�+P���c$n���;\vXt�p�"���Z��Z�ݳ�$�梤�t��d �98�2�! ;k�Q]�R�h]L��no�`Q犊f��zÃ��`y9	�#zl�|v�ϸ���SQ���
Zŭ�
zް�a��`�3n2�m��XW_�ݠ��~���]&��m��oaY�Ty�������y�J2R0o��
n�lt��~��<���U���J��ԓ�Ao����+��$�ڵ���>�V�.�"��~n�ܶ\c)�+�=0�]pt�TkF��I�dy���i0��	*:R�����-����s����>(1�m��]�1!�M����e'����L%�EB�����Kƥ32�O��o6n��My�<�$V�e�۫RB,<�%H�:~����wm�o���2V�_��-��d^y�PCղ�+%c?N�orKMBqμ�cQ�k���?�?��~�p�[�X�Dl?B+��K�Jw�������fm��3h$�/���ǭ ��`��:F�kW�+�8�.�p�	�K�pGi�P�Sw���*"A��+]�`��l�ݚ�d�������KJ���
��dж��Š���(�L�N6;���I������=�K��=���3
(r~yn��,��ξ��0L�#���9��jr�0�R[��ٽ���dr
�KGF'R,�&oɧ�fy�Bɹ?��<	� J��C?��Nv֝(���twҘ3ۣj*y���,�S.��Cy�z��#CɘF� ,s3�mΡ�t-
e_�k�9��Q��G�`��O��&��c�287���������MC=u	����s|�f�q� �����������?�����9��J�����'��((��&�|܎L��%��娳�� ��Њ�g�p�X��+n��hJ*�y�/�[M�o��=P�q��$�s��2�	��Q?y0Z�1FRq��(�c�zz�s0F4K�h��%�8Z�]`�`z7����C��΃�#$.�^&����#1.�eT���s�y3����j�mЪa���U�]h�m��լ)��hZr�����~)C�|Q8�>hR5G5O�Z�|i�B$?����Xpge}W,f�-��:^���DG�d�������5���J���imR���'����R��pשQ�̽�;dx��ΐ_\��8��y�Wa���Nz��a��,��@�-��wW�V?����)�^K��ٱ��e|#�j���n*�PW���
tZuU��}+A��F���%�Z9�J׈'ܿ*�J� �ۭ���f����z�,K��_Zl'�X,�[q��L��.��F53��9ɉ�ji�(�{k`�f�7]�[Žc������S��� c�1�&s��"���؟s��O����Ԑx�g,\"��ЛZw�a[�q������F���i�#q5���~�7!Vۺ!��y^����[]�`�4��F �	�R�p���^�c��C1WMU*�궝:���74�TxA�܍!^i�?g�8�P9��ҝ�h<�T�\�ll!�R4�t�a�?W����� �$z�^;ia�^
~�����f)`����Z�)�9�d�㏻v���q������.-�i�[9�s�b)"ҐAI�m�|l�|x��~��X�}8z*����aCALG߯���q��cIGU�m=H�(��N���K��� �X�a��� 5r��64�TwX+7P,�U:<�!YJ*a4� ꭰ����SP��ΨM��-�$���<8uy�d��RV C�Z:��4���_����r�A܊@Y�:�$�d�l ��6��w��'i��A$�Va�:�%|e����ɵ/� C���F��	� n[�1jQ�����|X�M5���]M9
A�c��H�����N䕴b�ƺ�R�uE��D��x!Ed��7v�S� �R�8'�Whx���L�kbP���:�;��}���?{�kEa����_g�	~�1�t�ݥ-_Z`�6),�9�J���o&!��n�zlY��A=�Ŧ�b=ГA�\��j�Ͽ��{�שּ=O�T���4�t&�:�Ӄ�Z��b* j��z����LJ��{z���?�z:>	�ŊkK�٤v�l\�ho��������L(��m�N��Ӹa���H�����A���{�h�{��t�:��O$�C?��IvP�ٻa1���ϖz$��w��%L��#d��3H�}6��EUv���Q�5r� gA�s M�Zpug�'l�L�������x�D]Y��1(K�@s"IƞYsFO�'=��Qw�{!�lmw������395���y���dv0����kSE��Hݾ�lBů�\�'#�N�I%l�9�w9��{ھ��䗾-�������1O��
�Π���.��AB�.�_k!~S��k���&ܼ�Ig���Lk��W�;M�{o34��������i��W>7�@�~�N����Sd�x�w�9��;��A�� ^��˟lnVl=�Y�;�M�umn}�eWL������5V�|:�v,��'����ڒD�w]��]���s�ު�	j����l�-y���X���r� J
ѭ��X�g�J����#.xv�����.���XŮiP��ڶ;&w�A��N,0O�o�S�f]�a*'�X�9 ���]����S}��,:�uJÖ��9�����5j�a/1�ʛ~����W���=�q�� �@���Ҧ��q�x�j����SHJ�[�TN�cz�&7QSg�ý�[�S������΢�H;y���[Z���x�Â�(z1�Ψ��v�,)����Y9K5`�ۣR��ï���Dۢ%T�~%�5�˪[ RY�e�
���N�\O�o��5fH ��4tcJ���g�(�~a�$��M3���Vk�]��-�l��ˢE��B��8?�
Q�i��'B0A�Z��/�ٺy� GSJ��#���_<�(ʨ�/�w��Km��cʟ��|�Pf��UJ�bz(6Lr��v�pd'��S��T�����ə��XCJ!V�Xs�1�����̕�l�C�L�X�{�Z�e�0i_��C=�i����uD}Qfe��N�$蕿:"+�fh䞳v,�����V��P�����eb��e8D�nqZ���;M���@%�/�<��kT��Y�<��u;��s�oE����q�k�,u���oFh���Q���@D�0}rE�����@y��0qc�a��wM�I���RM�S�b�rf�����*�hT����l>k*扫��0�.�;�`_�����0����[�r�NF�*r�w�Y���΢���#�B#Nm�4	SN�H�DDm�+��{p�y��E�y,\*��_WI���Ǥ��9�xO�m��:�=��7��Z��k)ؽ��=l��t���8H�X V"���V�YB= ��K����+����+��|3�j�ޔ�dq���r�5��Ҩff��i��򙧴c����L^��aи�tD��w�}2)�TY��3����(v�5�.F�ɭ�jM�1�T
8sEfZ�b����ef�/�Z~��m�,)�vR�@<�pfV�\�!	�Ra� F��G��4hةD�w��h���/p !�yɀ��^D)����u�Zzи)���c*�ǃ�Ѕ��	��n��-~�];��K��q�F�oN?JB_��8��)�*��W-��}�=�8ԡ�����Q�A�,8{I��6� 5��Vtf���0�cn�K�Uص�����e7'Aք�MCFI!�$����F	�!��js�����x�`ʡ�;6�XB%����LU3Q��=�IJ]Wy;OoF-9Ǚ.�ah�� ��H��_�S]*�K��w��1��Ov]�ϯYJǆ#Qp7���{Śm^������^g5�C�Z�N�z��K?$�M]{���k���@�|��ف�{sx���j����DƆ㡴Z�t:�q,~��*k$�n�"JR�xM,Qy7�C�ʿ|�[��]��j�S1|p�=�u�l�l���oF���?����m��`�vf�+9:�sU��B���5�B��Y��K�,�-��r|S����� ����DY��\�[�ң
�y�(� ��(������_�o�3�h�,8&�4�C��m4�)zԩ���W~'`|4�0�c�8/[
���< �.�dr*�攝7�EB��l�ֻ�r�(9��`)��-�����L��=:���m+���f�G<{��R�=+���b��M��f��P,�i\���
bM�HIƣ�r�W��k���� ���Y������;a�N.#�J��ǟ�z�,�F������ڤ���B��l��6Jz�׽Gl}�uJ�֢p�CJFe�R��4�l`b�ܖ�A�����gAU\��op��gD�&�#֩���˫��FU��ak�o���^���i�D�@b<�ʲ��rޓ]��PH��䩃M�SFJc ���q�}@"�l�Q�ѻjc�<�Z��'mZ:[luE/�Xf��%���DG��H� �6Yy����/�a��#)U%�gF�qj,J���+R[��/{UD�Sw�WȺ+��_I]Xk�P_B<��T[�9�{Vwoe��┸��6�%��(�=�څKt�m���W	�@쩷D)K��<:�$�m��5�T*ĝ�0!�g��ěF���������@�f8���|&�78����(����&��9��%i>���*1���><��8������5�a(bWR���,��X�8ڬ5��h��OB� h�5�'���K̉�і]8�*1����q�m���I�/чʝܰL�N���ז�z�8jܘ�͕���J�eo3��GX�#�����lW7$Q-e��B-�#��LL��1�Qt�H0���aS�9O�̴���c�������"���YuT��f��� �o�/H}M�I���f��;״��n��F�4Ď&�VE�?t��髜b+ž��ۍV�`�i�`�j��sg�S����ļ�V��l>�4��OU_��)�SV:I�vZd�s�a9.|��ijy��uz��<���-&��� �)|o��r�.�/O+w9��[�V�����݌wX�fazֲ��L�2�}�v�d��H���	P� "��FC�x H_���f��$uA~��U][d�#���fN�l�?	��fk�E�䃙;=�o�LrĔ><��R5��ʬ��=V.���ԛj��.�Y�t�n�y^3fO�M�_L6�8�EQ���XZ�<,����7�:��3���T�B0���}�!�,V��U�2���Wn5�[4鴚t���_6�D��f���F��gN&>k��&+Fa�=�ff�)&8�N�?���(,9+�8d���Oz�k�%�^�0����Vﳅ�J_��n�����0�M���&�R�)W�'%�@F陴u����̩B�Sə���5I�e!�J!�=g���0,0��!��e�$h-�{ؘ�]�[vfs�f��Rө�\w��xk���!�s�Gf[�L���R��_g�J��b��G��,p�v`9�=���a3+����1�B��,ؕ��cf- K_���Zg���yY��P/��>"���h22�?p*�(����u��@�,�¶H��G}�¥˾_03���p��iŦLwf6<u�j��X����>�������M;��O3'3Q�Zc��;�Ky���rT��vA��z��o=��H��*�.T�]/�~ɶ��"�?VX��j7V&7P�����>e���$Q�
�%�)��������9�^*Q��/84%p�A�D��(�Z�G�3��c��%��R��n2D�@�4 [���C�Bђ���5�����iu��b�#G��2��)�1��E��nSZMLd���9���4y�
Q�i4����OE/�}7/Hⰼ���l�����7�w��)��I�����:^f�o���tL���Χ���6��vZcL���gA	�%�AΝ�*���0E�����b}����90>�	H+c
�iu���	y<���x�r������{��9�3�o[ c��!��*��F8���\�A]��%V%�*�k�p\�Q���o+�h���z�C-dXw[��J�0ݮ�[�d-�$� �c����]�5��X~���?����J�(}ݰ��#l�����E�,��4*l���{Q2L�����ѱU937gqI���J^zoڭQE��]��d���"$r�#�h�x���*9�n0�=5�X;,w�6��>ƍ���~<�IPe��Ě��=��-u"Є�q�,�K|�6���g����\�R�� hN��Z��h
��7κ��t�s'�e��ȫU$mv"�9��<]F�B��Ha4ղ*;1����O&t�_Ʒ>�e��s�����<����6�c
4��8��C_�q'[������)j�����_��t���w�*`��v����E5(�҃��(���jE�Y���g�0��y&�Q㽓�b<����G6�r���C|���g�+a�ɳ4�d�R��ÿȳ<RX� K�3�+)��b2p��� �?�Z�U�SD��a���16)��fy��f8�E������Ħ�x�mU��31` ����7�0xN���B[<�sM��w��#_��5� |3	����'2���ڌă ��w�3�����|2GeѥَC�N���6�٤�q��Ħ�s�ga,�����������TO��K�<�7
F7���-FV}����B�:ǮG�x����д����,��EGg#��:������&���
����5?���׏\��% �^�����֪/�,�gv�p�z*���t� D�q��F����/ �t�m�[�{�5�OE�Ғي��4���$�Y{����l�����z
�}���@�G2k\��a���&N���?��h��w�j�b�g�C��K¼b��}m��K��o���[�cU(j�ΑO!�_�I�_�NG;�wm��,"��A�d`��t�瑘��^O��R�G��A�+u�t�b(��<+����#���z�L��B�K85�GK��V�Hÿ�o=�f�鴚��}"n��5��L_�KU��m�~�1�9����9�G<ׇ����#�#�5�i��۷.��av��A�Y��c��"#���Eb����cI��}C�n�����|�y�u�s�3�����l`�<%�=
wyv�9ں\4��)�wL���+|AM#��%�9~0ׅr�}��ј73ib�a���*�"+�mb/J�(|q��Ar�~�7�z5/ ���z�>�:1E��Qh=��Ey���s�n0��w�*���-���A�����|����Iy���W5��qj䗭,�<nL�4Fz�E��+�Ѿ� f�~-�����K���E���F-�1y�����Ej��.�Q�M<�碟{CJgI���0*υcPt:ft1-귟�#�)C�����j޹N�x�����Mu��d�\�G\s���<;�?�S�.gTֳX(%g��]6<�<�����Y��T��da�Uz�I���������j�"�;+�(Mf9W]t�-fq�������p�bs�G��^z��S튕c�`��e�x���H��� ;T�P�ڊ�|Y��=��hR�JR��=\�in�.�LG�k�R����t�п�>F�nV��bC����Q[+r���s�Ň�>6�~K�1㊶��t��9.��4��jm����>0���5	��&i�0:g����l%,u��p3����]�����
�[���UmdŜ�it��[���nq�]�U��\����C~��Vk��P4l֍.K}eB��Ɠ�N��7�I]�v�d�xR)��#�����������}������I�󕝣�l���c�Ӥ�ח{GDEp�hhB��Hi�#j����W���ѥ�O�� ���n�ޥ���Ĩ��(�!Kv�� �1����c&GE��,����jb�@�z��D��JϾ��K|�7ũfx�)��\w~�\����E1�B�PQ1��X��$X N�a�K�V%�OM��.kY2=
�0�J��P:�g~���>`�䍺P�ih��V����T2k��{e�|N^���ԩ�j�C]B�ƭ8��5��T��\8��t!�!�Ѝ���T��m�ZTD���v�w>�fH���`���(�RI�L!��b����<(�8�6Z����E�o(��>m&���,Z ���H�͇�f�,��V�@��]�AV4v��A�x�bo�i����(uq���N9�����<���'��y�Q�T4vaT�+����b�(V
�G�V4�ߔ�T�?��J��#EӝYY�A��j���}�!��ͮE�_z�p'�X��?�=��B�M������ژM�g&Τ���+�h~����Įb�!Zh�(�ݣ�n �?�GF#�d�J+9�����{/�
��aZb�p>�s�t��u�y�!RX�}4�t� ��b�'��h��[����h�>�Y)�(�>x{a�_���V'鍧��M�)^�s:(�����*ż�c ��pd�lrwf��cGP)~?�ʋ;�	9h"T�ۯ#������ ؍vz�Н#
K5p��r��F�쑄Qgr-�VU�g�U_%� �Xd���`��)������)�����9�J���:���'��A�[�D�)��}[��C��d? 8Cyٓ��o�f��;�m�{�a��t�խ!Kl��2��O������a����a�QW�A��z��V�0�l�z��������D����$A&
Y���}^��O�z��2	��d�r��l4ȥ!�N�FdK����ʄ��Fq��A���Q�H��Z��c0W���d��~��`���@� 7� �
<��������j�dN�Wk;����8�ϸJ̓�V��B�58�u?L���L%�VU$�ײ�{�I��{��+�f�
2��51>Z)�U
ĺ��e�G��J��$��L����;�-�6��YF�͒�B��-�K�װ��I�z��C �G�Ջu������=&dC]!�rM��yIJ0�*�u��8�!�Gۘ>ώ��W����j��#���[�0�O)jW���K�q�Y��#����е����}>C�.h��D�ꄥ����h.^:�Lgȇ���Es2W���v6S\|"���G��nط�"(O3/�V&ǡg�܉s�I�*��z�{��tҚ�E怋>vG5;1T�P	���$i��$���nЗ���������!�ldk;P|�G��:t1�>i��}˲q�F�'��g��{��1��@xMc��v^�,�kkQ{�<6*Ŵ��2�0(B���������&Ǯv�\⼸.�	�פ����)�55�=9�>�{��1��`��'��A���Ѱ(�ʾݑ�	wW[�d���8�0���I֍	��EqM�3���k��^<[��.p��X��.!��O��B�1��n4�8�>x�
-,��8��I���H>W�,�b>�7 8jOU��&��<P�ѵ0w��V^_� h�ic�m��ECm�[��$�����,;��p*���]H����D^_�Nԏ8<�m|��@�VY֔L[?��%��foP�/���F�>�C��#�Z}ƒVD�, #�^5M����H\��z�'0��3��f�A�ǝ�|N�V���S�9�g0����餹��k8nO/i6�~d�&���;O)X?	��~9�|�<��]���,����B8�5�X��=}�㴺"^[�R�rt|�JW�O>��M;�H������6�쩀c\G`E�S�iq�]�W�0�v#�d�}� ��{KS"��@�Ѱj7�t������Z�c8�}�BH��gT���-�*���|G�b7�n0ܶ����5}�%�^' 	j'@�Fg=�a��j��q4[90������F��,�����ȫ�iST�4����߆�=��J�Rr�1�l͈װ��A
$fӶ�K��?��
u�R�@��򠈈�.��iFX�A���1)4Wޥ}�,̒dߕ�*�>���^�j��H	􌎋���+sZ�^�[�!Q�c_��~T�5��,h�Wo��Iyv�&[Ģ	gd��N}����q�%����N�$��4���B��3��˽,�
�`zp���v�+1�����d�ؖ�)����v�i�M���R�P��rp	�\-v�z� ]p���$�j�V��vf�*H����)�q��oL4�!hȃ���>��jxq��D#�I��|��3�<6���7}e�4Ѹ���S����`i�{�W�ى�+s��T��pd��$�Ogk��\r�Y�oG�6�����L�4qa�����a��-7��*S�^��EMtT�$;5P�s̓v��\T�U��ͫ#���I���d���\}RN��k&<�� s�_�K�s��U!�#)"�N��x�0*�X@^��=�a�%Vf��bNm��Io��;J6"����=Q�(�������Q=�Q9.2�ul)��6V���eɰJ!ugU�)���'�$"Z]7�=iX�aŵ�CA�l���d�k��̿�f£-E������yd�k��D� ު�q%��N�G$�ޮ����y�%��]8z� +��"h����"�� ���ILTb�Sفei��0J�Za8/���K"l�?%�[��5^n�}���9 ��,����P����n-���z-�>䎪�qɎ^ }�(�,��A�1P���-,�a}�Fx��`Q�6�z*�u�Fi�;�OH�wG�9zs�Dfw���A^��}X 	P�Sx���":3���U��ZwY�0<T�)Ī�4)�C�z3�_5Ê�!�n��t�u�!�o3���/��"�ہUX����0����p���i=*�[E��I@S�A
�|���?M<}�i�GX�����=~�j�*:���1��P��QҤc�}�ۀ��.�_7���P&)x���7lx ��a�%pE�ƥ�R��Ӷ�%z��#�r����v+�:�~ΜQ�321lk8)�$�d힙gn��^��H]lǤ��:/�Cz/�J}�����3?��K��r˞�&��F@"e��M� ލD���"��!�T��2 �wؤ��k�k��m$ao�Q�-�>R�} ΤzNK���Sh\Tl+�/�5Ę�%�:y�M��l	1/�����D���b���K��pA� �D�0������)K�EW� h���<��4P$X���Q^�����!��д�����M<6���d�=c�1�Yv����1]nT�����e[�k�H5������3�I9hQ�7R��%�0�û*4��:�?�Ƈm�A*	��A��I>t��T�`��Y��_������nW���H���b�[�((kAN�݈꾧���;VCW����~S0`0�LU�O5��1ya����BNl��=���~�[MP�Y�L�ܾ��pVY�#����]I2�24Q��9 �fD]ܸ��K����b��?p9��)��m�&�Jm3��^��W�2PǱ*��ۅ�+IN���V�wh��W��]Q���`#|�A�J��v/�p��oP�5��5p��^�ʑ"�^Ѷ��(O���-)�����&N���K,)�'}nWm��xi�B�xK)J�*aJF�TzW�J0�� z��=ɪ ����\%�f�UA�G0g�Ox��.\]w~5	�
Ѥ~��	fp�����i��r�]#���h:�iVr�="�_y����ޥ"|v@{���	�wߪb61ͨ���l'���'4�oL9;����q���{	�,\���%��,�nI�߽�)���C�xsf~-��-��'�Z��dUGl��Ǡ�c��~�l�J�
\d�O,��& ���ީC���r4N�H���?���
X�m�q���r"�Mke
��y%��K�3u�9�ć�\���*[���Vl2��̒��C%|��������>���,]��}DM��E
{y$�{����M�G��'�r�x�҉������D$�;bg ��.?Ij��Ѹ�h���e�N�5kޝ�i�e	`:�y=��VLcI>
c�!Qwy�Êr'�2+/����Iz/�1sYr���~�N%�.�ǎa)�%�09Q���x���AQeFdܪ����+)i��#%��#�(aq��e"|n^
�S�E#�{���0$v����/\HI�o��a���O1y�M�#Z�v��=���i�s22�-?[mj�����0�����P^�R��~����̖5bv�Z5�M�jCpDy45��*LIL0� !���P�C��ڗ������a)V�G~�C��Q>�,uf�A���E�8$��s�C�l���Y��S���� �J?���K��ZN'R%�A�9NQ��Pvn������눃.�7=���z��[pJ7��W���IW�3��I)�:n����Tv��$��铖��P�h�-Ib7�ͭ���O֞�l�a�Nw����EE(/�������CɫοDjW��g�H.�Q�H�,�C��Ȟ��:�!��ψ�0ƽ�I�'Nri���I��n0�5��<:%z��tTuJ?�e�,����=�g~@����?��5�D��X~w�.����e���Z�d7�n�Ҥ?6�d-o\_�R�\�()��
���!��W��;�a�<B�?a |=�ݽ%�=mX�pL�N��E���Q���x��h&n�5%���r����P��]Hd��Sv����p�؍�|��P��G���o�Z,pW�"��}�@d\�BZ<����C�� L3`�ioJ���]R��/�9Y��gn#��`�)2�_�E���I�V�%�F��&<|ި��,ƞ�=�&����l�8�]� �0��G����5�
�+p�9�k� �[�U&*�&��/�����Ʀ�э�"�*A���9�q$��4�>�Q�\4����"��Be�ȧl�u����KK��d=�*�M�H|���412����VT��l1���(�9.�x5)!�F��33��f����9<9X�d� �3�<NV�ow��bƵ��m'(�ƅ����G�9�D4��2�H㣝�k��@�x�#G�Cr��������|��_k�p�sCX,M�F�r>��K�{�Ȅ~�ʣ��m����C�q}�R���a�S7F\gV�a�<�@*��Qb	�[D�n�z�U��)�lZ��Do���aݺ=i�X�?�\��r=�����n�O@�~��J@m+d���@�ʠ�q������-%ø1�f�R��a[�vx3�J���O}��i��exp/��C���X�B$5�0(7�Z�[�A�D�E]z�l��<|�+,�ډ�@J������|`�4Q}��H`�=^J���Kb/�1g:+�@|k�Y�b�E�p����]�o��	X7}��^ψ+O�ʾ��7l$���6�U^��t����&S�l)�v]"�1L\����"($�oK�WR��]E)b�ӴV��U����M��%�7��	�O�]�װ�f\Yz���A�]������1�7�i��3Z�(�&*yRmQ�t�PaZ�ۄ���[$�cL��N�>r_�3WU��6<�9\~�t�џ
�Xz;� N� �mH��j0�ȃ��?�'x1���7
QYiua�p�7��&t)ݍ|�]W��P�a�d�5�[b�^�?qR�|��-_
{�KU������}�/��mS��q���kgMM�}�<�~�~ư��q�U?�t>��Z�i�G����:"K���u��'�^��a��.���V�� ��������A}�W>�4��6�����/mP�X��T�zy8Q&�Q�j�
������G=n(`c��j�^���S�>g�>Կ�l��v���!P���)���M�e��Z��v�HpA��40��C1�3#(�
��dHn]��s�ᾁ�(��G��~3��4������	m�8W�����RM���m㫦�1�|���P�5���ef�d��������r�G�;�m�l�O��>XK�2�(M��Ά+A���Eñ�H�N��0�X���@��O�0��i�V���y��������R�R0O�-�G@4�;@����,�7\�2�V�2ai�|m��[�w�@��.k���$(��!�0�V�$T�?2[�s�}���lAB�k�Rt3m�Tg�r��~��T�z)�6Oe�s��bz��ZC��RM���v�(>[��@���UXb���'�e���*,��4�l$X�T9!1&�W����^���5{I��_$��<�1�b�y˂�5<B7`��;�����VS��VF�����2(����P�{K(�Q�G�rl�#�J���v�4�M�yS��`0�p�:'y�NŘ�^���E�ż��Ԣ6/|���-)�:�*k�(С�Ĭؙ�+�^E]O,�=Dˁ��.��>O��pȦ�e��B"��h�-�����ƫ��0��k�g뻈��&l�Qt��>�9�JS�U�W�CõB�]w�����y�K5��qӈ����M~�m�,m=l�[�i��ڽv����s��_~=X�[FE��~*ټ��S��|\jF�ļ���N�4C3���W�@��O��A+�#�ݞ���7S6�����-ɐ�/�u�խ-	��j6�n�z��;��ŵ#���"V!�S���P��v���0�3�H�u�I�����M����q�@�a��8����Z��g���g�����g��@�I�x���
^��4������>���F���Y�P�a��:���=��#��zc�b�Y��Quכ��E�߶�E(�KB~֔�\��g[(�o>� g@0�J߽�f��?=��n������r��}�@�S	�'������GO,�*�8��g�q�k�FvjL�.l��_+���vԝ�?ĮL�v*߉q��ʞ��(�_2�B#C���wI6U ��
�[
�)�.5u�>��JJ�vΫ/#[k,̑��p���P�)��tƊyV��RP�ڛ�8b�P�\���r`mf-a����տ��}�e�_a����)�Xs8���(;�S��}�Q�#����C�O9��ڗ3G�H>���9�X�����`�x��mYO }k>h��xMK��,޸�2ٚad���ں�U��_�)�5|ę�l�S�z��I;K�J���ͤ��k��*�m��Z��i����~�jrra�;�9�@��;�o|��:P����}�b,_�M�vY=��0O��"2d����{�U��i֤"m�;�Ɣ�/�e��j�C� ,䍩��ψ��sޭ't�.������������2��ȹ�ǂ;�}BZ����S(>��(�)s��-�R�t��gZ��؟ZY
y�mU�g���T����DW֐>�Y��׏�T���Z�H�Ӟ�w��dA��;'�Ok���
$�	"�n�*M*O%,g����kl��t�AQ���/��:�|�S�xq�O�O���M�o��c �FHl-�Hy�C��WB�wy��e�)����O�~��x5���)�$������üN�KS<��Ҋ�G�&d���h6L&Q�BhϹE�*�0T=���\��:-����
M�+ON1����9Y��*��,d���R��d���#�������O�T�l;�DlF/� �5��ոM'���\���$~^>W.Dd)���ʟ��WRL�ә�
-���榛���lШ�(LS��*�0�r։И���y��Ôr�������{F݇�/\��AP��������ꂶ�ke��\�U��26�/��t.�ED5�A�s+2�������������|$b�K�ط��$���
����jx��h��C��)	`?��B�0.�DoP�D%��׎�Q���ll��.�E8#3� �L�G��/5'6I"uČ�������X�YLh."�"��cҖl��/~2�`N4#���q�IH��(E��eN�R�OI냮'Tp�3AYI���e!d��[`�mV|3�b�F���z�BarQoy��x��EN������>,6ۆ������-Lݝ��d����=��Ĉ1��u�q�q��kO�%�gCN�ׂ�Vh��3����Apε�Cg���.��!��6��7�1"-dy|�S�@�o���j�C-[����x+�Uz\8Y7-�h��R~o��د.�nqR�k�6ρ����[F-����T����:yD/���fpPSYrxG�=�,!V��K�Ev��抨Ki������ ����5�R��խ�������Q�����pZ�����V���N�s+
k�<�~5��0/�9�:�� ��@n�6.���%���M){-��9���%ғk���@�`��x?�@��<����bw![���f!;���W���:���������IK$O�S�B�!������'�f��,�rh������M����/�n��@�K�ℴ�镮����e[cA��JO��E9P���Ь����r�Ϣ�L�?f��8y`o�@�QD�J�Z��y`�U���NևC�����|�δ�;��dU�ڵ�?�e��M�|t�IT��S�"Y�U2�[�GA�� &��n��
�p�q�e�jP[m��L�MU�ޔ��+M������HM�}�^5�X~��K��n�Z@X
��!�$_P]��a�^���̑��`�H�_Ӗ6W���g���d,bn��G�o\o�����:RDuF�yk��u>��:	��Q^�۩e�J~P$2{��\�Y{�����\�&��PwY���K��dq�0��V�����	9/8�3��i��w�qS�uQ����>�����wb�fa���/��u���UV�/�ޭ/��U+<�x�}<�|�����2��z�0Q������,%7��Uڧ�Y:@b��7a��K�e��YU/e�]��#F|�%P�c:)-�ш�2[i��|�`�R���, ���||�����Ai�X��m�kǿh�{�޾.$�HU��M��Q �b��OSe�?�7��M�����F�2t`����E<|U#�%?���=G�����!j��n�J�9bn	?g����8�_}.>�烓�
.M ���x�@j�ɸ�<�!$V ���ނ��O��sBڈM;�����K�q�"�/����f�>�j����a7+�6���%�����D�^������>�l�{���Qk��b4
K-���_!�������Y��/��%t�ÁV0�l�.����͡	PI�Ps�݁P��+g��*$\�W�A� �q m�8�sr2��;�� ժ\������ny���Ax��wq�6���/�50��ܻ�OI�#ѝ#������I�e�Xd���遪s�w��;��5�-i��1�``|�tm\��!��M�޻�z�\�}@�o��]z��q���e-��_�Tu����e��LE�O�
��8�m���� ~X�"ꮰ.W� Zd����Wgt^����Ӓ�Æ�V|��2VNr���9Փsw} B��&�aM�x�}��������_�U<��b*?���9����$!C�Mb�P�;ڃe�w~� ��!�{�0�/�%�������Y�t�8���F���� M�hi����]͹�S�Md��υ� ^�
�B �E�a�5�Iֻ�&rb9�YW�<d8]�[/�Tѳ	Amt�&i�3��oзcBbv��5`�ɶ)�
1g&/��Kzx�!��hB'J�&X�u]j�贅�O@�z�6����T-5����Z_�ޭ���y���W�t
ۿ^����y=�H����.��$�܂,弍,d��c�:~v�j�l����-XzQ��MFQ �z`��S�2�1p7��s8=W��cq*�D����;��.�.���Ϡ�]���8��8�B(�q؞y���h�Q��I�>BBf�i�J#�A�?�+��7���"����	���h�
��)}86\6�Y�~)�ܙ�Y�EQ#����"��ڙ/�a?���pH+P~�
�/�˾[ǆ?�=�G>��*�cT�X���`�j��d�Wjf��I�W���ڄ�[�Y�Q�'�n��������)�!��l��B¼���h�?��gl�*����H
�
���m�Ԫa���Ƭя�@��R5�zR�2Ꙇ�:��5��W��w�P�N���Fo�TM�*���VȥMǐ�)��y:v�(��r��Ȉ�wg�Xˇ�N�Ho�lC}� *�{�~����֑֟��c�k�g[�r�pX��e�kJ���|��ϴa3D���;��Rh�a��>���O�r�o�oa���"�.��QN�Ҙ����V�M�^�^�#�H�>�`����騊
+<�.v,f��3�M�j��=3c1$|�<[�`�yo_hF�4s��J|{�� �k0U��k |�@��� �H��o�P?R Cf��:di%��1���S���҈�'~��&­35�e�8� �7�ȹ�÷Z�a{��q�oSRS��u�iGo�hJJ���4��)�]�������7��c�V��=����a;j�� ? ?ݫ���9��КN��i_�}Ʀ�
Jև�+`�s�rR@�ff��M�5�E�0�c��V�]z���F׹G���,���Z�4��=l}x��E��Ҹ�.�3��sl�DwpW����TP� H����*8�W��.�{a�j
{� =IS\��3jQ������Q�n�M fW�-���T����:�y��	���"U�ma��-'�/ا��b�Wܥ��%8�l96^޾�3D(�r���	��&��H�yʭ�C
t��Kcm�pz�m.��4Xl^>1M���(�I��ш_X��p5Lk��O`h�nĶ�f��l����9&���л"qv�UIn�i�J�k�V9c=<O.�(i1m�==5�]�.�y;�Ŏ3��V���E����'(�5���|�}��Cj��E�n�$2!P�M	C�iB���`���9�I�?�PH��[��Z���"Y��5�JY�.����Z�w��J���� ʏ*[��_|)ZCVu���m_�J^Y��L���{�}�p`B���%2ă.�ec��RA�}^��)���X��*%����U�b�$�p�:U�<kXY�=_b���C-^����¹�N�@�D��(�>�����=I_��Rz ([�h�a�$z}��� �Κ��L
�4�e�B��b|Q=a8mR�2>Ie��O�y��2f�[j'�c�W`ﵝ�M�ؿ ����AU���8��+2Ž�/�K��>������\S[����N�:7��VE�p�f�T#j��T�̽m��	�۽�c����iX��::s���}�c���ETP��$�,����yq~;�e�2��\9Z\���뿌*!=5��v�1t�C���y���j��[����UeU��:���W��'4��9!>�b#��]t�p�ʟ/�IAՕ���4 �eQ�_:7r>������R"����m#��]��8;�}���@՟{��w�u��*�6��W�rB��I���kVi���VNi$4��zc.H������mܲ_p��S%[� �|� 5�<��)Y�d6�b�ZrȰy�{��ٞ�֭��+��@��&�'h�C�9�F����Ru7�c�;��t�H��'믿�"^��eL��F�N2"<�t-s�c�Ӫϑ��n$����h���A�x�����/�;�@2:n�(%��}�����o�׵������1E��!Y��&�p��0l���d4%�l����f���`�Qz��!�ȁ�6�W������VCÆ;��'�2/�U���Ī�u���`��kD�Un�"6��si*�c_r��TO���EÄ́�5�ʵ���N��5j(>[|g2��2�gq���-��1+tȌ/ �3k��i��^�.��=��Б���q��2`&wedZ5_�OՂ�'Z��q޾��#�S~��⎦*P{���^��9i�o��nj'�GuQ+ЛY�=��u��$�O���z�9y��'�a��F'�m���w[���r�(-�hIH] {f���<:R*���4����C�h�`�D��� �F��6��5�*1.�l�@M���Tq����VG�]dw����W�Z�Zz.Q�Rt2���1*S���e��>�|�}���J�M(�<�*'����j�����_�]Y	��i�GL�@�ff�?�(`��&�@7Q	/^w�.y�(�Fu��ː��Ŋ�>M��+���Z�5�۰Ȳ���.��Y����ݒ�R�X^���#Iϣ�_�D�G-�Q�WI���������9���M���UX�H)�EZ V�[)��1�F�>��ɽ%�t{3��=Ww�A��� �FhH�{#�
�z�B~hb�b5Q��6^;�1v66f���L�*Z�Y%���Sms�������-��a Rxπ��V�.���6{���j�tA��9Zsy�n�����1�<A��������+:�R�#�Ξ!����/b�Cp�����d)u�5fw�?��x���(j���=��,�����3���Ij z�ؒ����q�ߚ��=�=�8ܘZ���E������3+Cѕm��S�W�/�?Ԗ���3ym̡JX���ُx�C1����<�5�P�w�k�^(Lh>[�r{��OO��g��%��N����?p�Bo��WuȄ�����C��x�%5!�s��YX�y�nT`]#�V尫�y�k�����R�k1��[J�0�2:Ĝ���U� ��!�
���E���&�#g����dEhǸ�~t d�;�`��@4�bA�K\��ǅD% e�%�v����|g��%�^$��&�qga阧��x��3����&Pl��SM�&������R}�l�9�.wp��x��!�|�
�4U?w�TCd�w/�<�� �vJ�Ҏx��ق�0R��?\��.%L%�
�F&e�d��Rt�+�ܒz͂�Z����гb���1�X��e�`S%��r!��="�w�/�d7z� ֖|hI��[l�eÁ��;�~/3�|'���+ϭ-pћ.�
�蟴Vi2-��x�8���Oo��ƤJ~��1���j!5����� �O���G-$S����?�AF��y��\(�n���D�˴Q �<C*ݱ�kꖄ0=����W��.�D50�MA`h�6\��O����e"�HcK0�����/�_z��, ;�[�|9�B��=x�/�?��M����``�Z��۱e1�5�R��_0������=C��B�֠i����C�}�~�L^P�z����A@9H��@u�s�@:�k'>��� :���9��]�C[�W�X5�*	|s�,«�!�H�ݔ��s�+�1\�t_����Ui}�Q��	m@�υ�a'�P�f��G`�8]����k�/Rz�v��(I]��-�s��0|�!.���2
�����Y�Eb�iM�OL�5��a���-s�,5Y�(�5�|[k� ��O��$�sH���wj�f�Tf�HcX��O�q�=~;�e���H(�}WĕD���h����<甩���+ͣ7Y�Ǉ�[��%�	�ts��L���	x�i:3J���䑳�^8�&�=^&lA�r��5��f�}�50�З���rx�$��v^�9�ߡz���z
��C�Z:<l�*5�V�ښ�0�����%��H�Ŵ��s9(<
z�y�Toug�����h����.�_i�5&�9��h�7�sl:�o�f�$�|e����H&���'�>^�eV�������0Q2�
��<l�j�Mߨd��ځ�{ӏ�D�	���wk܇:)�|�����o��a���%�!����-CC��(q�d����2-N7�r,d�E�|lxd0K��@Z�����p��`�)Z���ӆ5$������U��~����N��	R 7���[�%��h"�a����lI\>�S��H\��%�\ײ���Ё �y;6Tᡞ�G�X�I�b�Zgl���Р���}����1d|��"�̻*�o�$K/��E�Mvs�i:��,�`Gl4`�	�ߋ�vEa2�YN����7;�Ɏ;��R�l3�ҁr^�	� �̛�r$v83�ܬ�.|�6r�!��=K� F��zS�'X�S���,���>	k\x! L�r������`����{t�5��y���2{o������r!�u�ӗ��3[����r��(�m�l�Y�z_H+�mAld�MTS�Vl0h7�B���aBÐ<��)�!�F(G+��	�r���t����>����]��/�̤����n�Vh�r���euV�G��\!���@e�I�>�O9��O�k)�+�rS@�q�VH'�^;sԹ�w1VdҾ^H�mShOx��g�У[<r0���Բ:�M��%����={�.�D*J��srGs��S+:Z�I+[�G� ,x������1���� s@��Ar���z��=6�us5�>3p(e'��
A��$6��u ��Df=�2k>�$2V2ƂБ�3$s���~��@	��U �s�Ǆ�kЖ��'@]s�VO�(���d�BA�Y��g����S��1�(Y�� ����kŞV]Xs��kP�=��U;��3Z�MP�4c�
���/���o�gzi֜�\U�KN��)u�Ӧ��я]�b=EA��^���B����f��x���������\����xѷ�$�|��B�Q��>^��- 뭍��2lw�EƔp�HIoM�8���ێ�<9e�&	�:6J<�K����7񋑬q��Lśf�~�$��Fsl���!S����J�^�{�neq�w�ۈ�W��82�!��b�j8Ɨ��c����o���,=��Ke6d�o=�O�B�J���������$�3�±�H������;����s߷hu�A�r��25ҕ�n����t�\}\��4�[c�XU��a�_���`���9�L���ܽ�v��ϰv�A��!��
ҠK���9��ba�N �Z��X�w!q���ߺ�(������f6U���J�A�A=��.ܨ��׊m�|l�
��^��$�{1���B\VD Ł��𕋭���S�C2�eQ��W$s
�2���|�I<�9��j��п_�9ۥ$E�u=�"И����:�9w�n�y�Oê�|-�|8X2�����5{f��ST�ym�kr���\��	��$��"�[v7�M��G22��	�����#w�ݦ�y~pJtfms�S�jZⱺD��(�R�k�(�#�~`�;��ԢE�T u
��/k%d��wA�}UiA��v%��il�s���{��x�>�Bǔ��8�]r�aG?�3�_�p��iK:vp��q��)�ͩ]ظ ς*�!��I ��Q�h{��h���=�icma����}�s�+�8,��:1�L�����`��2@�A�=�X�TJF��X\�&-2H�%����t���l-����,@�t�_�BS��-iJ�DzV�C�؝2����O�(xF�n�C��3�D����t�c��qn�%	�(�(��$���;��T���A�P�?m�����5��<唄8�߭�rc�6'ɻ�7I��xyj�LF�g�����ɔ�ob	����-�ԍ[�8��xAS��{U���K]��!�h	�����Uq^!����UjD�̺P"B{(�rq�r�aIy�d	+��Rm/v͞���a3�\֭��=�]�GY�I�<���څ�7�=D���}z(z��ds�GE�e�I�X'��+��d���6���Ulb��D�	�6�=��{9��+���?��K�LT���e�z�4�N$̿y!Ŧv1��"Csͭ���~�����AP*k:6	�I��W����2t[ŉΨ4}�q����� /��,�^Ws��g����Yn�E��߬{qIǠ��b`�jwkld��̚� �Y�,(l�ug�"`L��j�lu4�S�Ux�=X?^å�>aHĝ�r��`��̈́��ַ�2̏lu㦖�n-����F�m�ArL�!J^����9K�m3�2>���l?��DV�� ���o'Sv�,?N�]e�T��N�����C�Ǔ2@?��������a��r����;;g�G��Tc0�&I�@&��@ `|/�\��`�w1�M��[��r3N ͟���n;$�l��Z��&�#�E��.�:���f�7�i�0w�����E ?��NE⪻�{�P�mQm���0�dp� u���׈�b�bF^������/��`WN]j�� 2���\��[�o���*��24:Y5�Y1�o�j�6�0p�#_-S��̫��q��4)��0 Ӂ`9��[�b�a>L8oK�5+�r��SpOD������]��Ú�k��Y����^�Yj��˞�	P_ȳ%����uk��u����;eh���g|f�0vP^��x��L� -�tGDru�w�
��<kf�P�|*�%��$������¶vG.I[;��A�~� �hik�l?�х�$�(VCD\4ƹ�P��i3�|���UW�԰!*�4���"V���4�*��7�`'�?3_��k����T1�6Q�F�qv�CmJr�cv���F#�?y��D�����vؾ;�_Gp�O��K���Ek{eIڍ�&֋u��Tm�<��`��}��+��
������ִx������y]��%��E8)����VI�3Ǐ�Hڀ�.&��ĳ*҄Jr�$@�s�z�B�o7�mg�6�/솹�ob�f�b_tJ�.�3�?N#dt��,�C��{J��ˏ��w7�������R����y���a�[Ig��`�qI��bȕ�N�*��[D�O[�8v���huu�Aqz/Omizp+��q)E�>�k�r�!�L?M��ۯ��h{i�T��3溠��^�r�h�H��t��	��9}�
�|��X����?.���P�UR��派ᨰ�q���d�޳�<�6 >)q�N[��s��R:;u쾭��|�*i�v��i����j�/��~f��"��߆^y�j��'���-���+����}�(t�>HFۣ�I()>>���t�s�G�,���NINY����t�+�W{R����H<8p30�x������x�.r���[�GgEv��6P�?�A��(^��Q��=�1B��<9�Yϭ�I3XN��L�M��oyf�0��� S��2��(���%���V6x��G�Y�׋�ڗ_��h|UsI�d��#2�� �Θ�w��y����rq@�}���g6m��g��4*�Q�S%�=�f��с$|�a�=I@��+���Z-��7�Y�r(���1O�T�&dflg�eF�m`Z/�!�'�}P�i.��*�R���Y+�U(ꋪÖQ��;˅ �I�����f��Y^�)�5��[�⭁k�	qfBeY�Q����:�X�g�Qf��45�]�7������|%mʏ��rQ��qi/��3�����Ǩ,a)�`]ێF�����C�{ݞ�0xE����w4����p��4ڤ��f~�����n�R��*�u@r4#V6|�+�?����R��8TɁ���u$�O	\��� �{S|9�*y�&+�z';1S��
�>/�z��<Te�)+���O2t ��R���{~'�Tt��t(��(?1]	}~��t�m垊P�����v� �����a"Ȩ�K�k�9�|��sz�c���=�X�����A�9���Eh���x��qb�K8��]@�A^������\h��:��<ly����i(��e�s���[*[-�QaQv)�>[E�p�λ��j�$�g��H�m���@���B����w蕊��Ɠ\LU�O�HG�GS��ǥ�$��J�VI���{�A�^�Η����Vb��տ���}z��eĕ�zWFn������@�V��	�s���;��t����伆����B�K�-:y��&X�xr`a�Ǝ�k#|V솃E�Rl���l	��L!��F;&�F��
�F≳װdMY���s��k*��6�O)�~������)��,�^<���w��#[�MK�����c*���N�oW��<.��>�x����[Qf?S�I?�[���k���L��f�_?�J6��d��G�4��11l�r����D�|���P�wµm�C��_����W7���ׄ��P�L�K�5�*$�>�����6���W�>Fjjj�������c���'�$�Za�a�P#�����,V�!7{Ę;)�������@��YW�5G@I\�ތ��þ�b�Ǎ�p�s��R��[���ɶ�X�*��gI�cb����y8s��ۗWBD����O*��k�l��g�A;�@8$ი�ٛ��˛fSӅ���[�9�L�:~�4R/H�:�i��qח[>$�9::�)Ȟ	ෂ�C%W��Z)�$�Ɨ�C�mk�K L��~R�"��������q1[�K�`�)���*���V�R��7����D}B�[�&Jy4�J �YQzL\��'$�@�Klcgc�;�0J&,�K+��ͥ�7:�X����4?"����}@�WFt��N����W���� �Mׂ^@��`�R
�%f��ao?�V�cT$r׏�Ѕ�~��S�	(�߬c�5NrSSiw����Q�ΨǸg*�i
xYR(���i��w���ɿF!��FB]�d%;d���Z"@�|�?]-rj-�7>�����%m^f��h�(a� ���A�������c�����A�Z�������kq� 6i��2��p���.���54���\�U��� �\���q���r��;�Tc&�`�e#h=�a�EQPX�wɓf��X��J�@Ӌ+Cq���K��5	������tlUNQ!���o��e J3WK��p"j���s?֮?�G�\��oы�wU��zӠ�#F�fg�v�O#�/-�㹕���3�0��_˰���@3��:P�u���^Ś�S�,8�ǅ֜3^���k�ܦ�hL�)���k�l#+H���Y~�f���V䩝��+�{1B�}���� ��WT
4�?)`5�3��8�CQ��3v�����L;�q�40�uG�A�:}�"�N9A���F����>���{��3�?p���D�[�6��gPb�	�wm!]ǌ�>9�2{�t�*c]�~���i{�AO�Yc��x&I/l%��턝�hg����LD�Z-Cu������е�k�V���D�P�Oێ����c��F����/�o,�t���N�I0Y!E�Yj�Nx�&�4�r��@C�[�yDd�\oI���{������q,�'H5X�S.^c˺��-����n���!q���v�"p��r����bιEų����򊕂�ڱ���G[6���w{v�]�O�����fKxר>�zm.��ƀ�B��h�y�L�Z����ޗ������K��xA�}�M��Y�w����[�PC���R����ːB̴v�i!yu���M�F�ô^1�~��Z��%���6X��%�_<=���C7�1�Ań�[�˟,���-p�t���3�3��`Bd�5f)������y~�/}��yTh:]���総�+���|J [��6u3R;T��>�t*�v4�)w���Q{)��*���	�}#�����W��&���;��o�nSG�p��Z����Qe�� Ρ���b�mf2,��*#Ա�(i����!���꠿�v\NƄE�!"2�h��Q��s�`$�Q.\�[ͥ����>u�m��I���ckP���-LU���Ӌ���l��M1��⸊V�w�s	#�x<b
�B���4��(�Z(?�-p��R	!�Q�rj�0s� W~���2��r�U�]����=Y/�t������2Qb�_�������_)�~�w�Ef��<�US�E{���c�Ÿ?��ӘN��w޽A�d��(�W��س�^��9ъ��C�M&�on���|�,�f�ķ�2�˪}�����
�Y|5�X�V�9K��bgd+�%�y΂�ܬ�Z�˻����f鬻 zYq�	�����E�EN�D�4�A�n�&iO�Ug?�E�� ���޶��6�ֲ����Ӛ
Ӑ��}^�,��R ��E�N�9vDC
�1i�!�GDզ����qQ��uWyt{u���*�!���/Q��T�3��u������-������2�롱�#KN�Fy����UC Z��a{\~����`ZZ1ks"n>K�.���Z���_����$}���*c#J��1���!�F��Reۯ@S9˧A(���O���O��6ѷ����(�ԹKV�d��H6@�9��N�.��*���F��H�����X�U<�ilx7�. ߱�s�S&�v���W'��.O�pKA����	}��IQ�U�KD'���Y3QT=�G0�~R�4����7ZJ"����Kp�OAo��U�<I�yG��~
JG�hY*i��#VE2�)��xEдX��Kw�k�.�Ѐ�؛�Û��r7J6�,��U�=��0�f�A->a��&��Y1�eAs��w%����{_Wѷ ��e�xx���)�� �6���.qz���1��ՂI�L$sH>����Ez٘R,�x�QAҖ�(,�H`�߽>ģ���n�/�x��Ȏ�R|�h��n�Y�),��-H��aCE7Fl���y��:��V!#��pDQ����rts���eܗb����
�y��^0�	�Z�-���$}Ϋ�m�p���`b>Ƙ[?uv� �7h��S��y��2�~_�Q�,J�轊���8�u
���E����K������{�����M2�l����4K݇X�սh���ՙ���R^�]':⍭�p��:	�k��-Xg�9Z.@���+�Ƶ�k���*kY�dF^� ��I����RT�Ǚ(PE�[Z@���}�c��Rn0��]%�n0E��:��C�� !|�������يZ�S�4$�Ѱ��÷�񇔻��X"��i��CNȚ?9��W!Ӥ�*�86�h����/$h�&pJ��e���#8$'޽�b)UO�Ft�Kk�I���;�pX*���톐�A4Y�prڈ�S���w�XP�S;��Mh�3�'B*.���Aw?Ar"f ��(���p�cfV��l����]*���r��]�3 n+B	�FI��C��d�,��K)�j#���h�D���\N�}Cy� %�_I�l9�ص%�K���1�O��}Fy��9��c<�:^��&�O�4��}M
 ���A2����$Ӫ�����WIGj���`���e}�1��1��]qF��'��s��V�_��=wc�wm���:������8^r�n��\�׷0��X#TB~sHBh�z:im!��e���3��=w����֜&�?%$ֽ���#��c\*��+؞�S[��T)(SC�����}s����_�G'x{����H��L����A8�H��F��>K�^�D����nJ�۴=v��y���d����F��I��Ϯ,�_��g����c�J���f'����J�s> D!r@ @8X���33�J7�+V.,.F:�n���"~6���\(+y�xNT�l�ػWFj�E���R�}=Y�0��3��<|^�og?�!�<ڝ9"{O_�0�VTk���M�
* p�@�]
&S���4�����rgՁ���Cr�@W/hȾ
���N��Ix�x9k�ߍ���Z���D;d+�Jݍ����l������i7��R*�g�c�/���:���*�ӢzĬS5w�9���L�X��?����ԯ�S���v��p	�Lrg�u$Զ�DI}�Y��]՝�B�`����j�[U�)� �ܑ[���B��e�1C�����^�Ó��s�b��O׮S9��-9�h�E���r�T�<�ג��PCB����.��4F7λ��.��l��l����7�!SJ'�_�+���H�a�=r�U*9��y��u�|x%A�`�+�����v1�/�
Ǿ�m����V�M�PBC��.1'`f:{d���L�����y�x��k!M�Q���*�˼�}��y��NZ"���9/+*�DJ��ǲa�\�T����a�04�j�-�*KS�}�V�ߒ��-����B�5H�r��\Vm�*���W�9�A�G��xh�6���*��C6�[|3�h����m35�C3��
����2v�����F�(�(�r�xt�3��j��`QJ��f���������o;����[���M����>��o��/�K��L/j�r+�_ � n�#�b[�ҐR�G�������l�)�|A��x���L�'K��ٷ�p��tGte�&����WM��+�e���k!��(Gz����h�';��6�#1P6,_@R�����b?�cMluP��R�.�1τ�Y��Wf�x=�u��^��=�{�ے���%��wD�x����7�֐��9|�?/�����"�{�E?�̖��Ǯ�g���#�>ky$�NҪ0�ⵅV�!����x^̉��9������sP%�s�J@��F��j���K׸�����Ny�T9d<�"����E���/I
tE	tœ!��%����������4���4+�.RKGk	e����cS��kx]�r�����׋�b�1MG$�6xՊ�k\�^O6���=�ׄA�{9�uu/%��6']F��'��؍HJn*��d%N哚R���"ꭑD�тG-r��p-'�b���O֋:7��n����؛��cZ�����-<�������_d��C[�tu	��=�ߕ7v�h �0Z	b���w�'Y�)V�y���Ko��'&��{�ꃙ1;%��N�W
�\1N=$��zP�F�P�<`q"����g쇩È�n�`���qR��/=V���R�<��8'�K��M>n��C|��m)�׽�B�J�#�Z���}�$�I �{q`����]��q�&�/����-Ó/��)uC�&��w|��i��0���?=��(�N�,�rGl��z�J�
VCv�*N7�,�Yh��a�2C�O�m���K�W�g�������cV��g������XX��h��DET'��:�M�՛��߯�N"�<-����/�J���w9nk}����� 0�QؽVG��8��S��DU��̴�\���b�����8$GBy�R���NW'i=��JCo���Ѹ�%apv��P7�o;-e:�nsQ{�h��5��~�#c�չ�����`6CL�xHU��AV4���=*���˼Rە-~�,T�g�M��m�}�[�����]�y(%���P8XK��ܾ�+��=g��+��L��ٛ/�5�*���%3;Gs��G�.d��u�*��-��������n���6��qq�OҘ;%���d�<��
��>u�N���D,}�m�� ���2��U�	#E6ʹ�+z��v�my-J/~�'H"��m��3ي��z�z��Q���m�d�Ju�����jYU��<�L�T9:G�����}����h2�2ˇ��z�֧���`�%���G��@��r�%�?K�����O�2�9_����L���QA��U�j���|�;�pM�'e��%�����uFKd�1bu� p�7���B�xs�Zro�?c���1�t?Qڲ|����rl@֠U�<��V��I,a*F9��1��߭������Zr:�SԤ��vT��2U� ��#/[��քu��(23��p�J\}`{4��C݂�}���c�VkfSa-���j���T4�ŹJ/"�)b�ْ���>8��s*"6��:*2Θg�K�j�ޜanw��2f�M�v����i���	�l�. m�ԁ�)�9�Λy��'0ǾRh��61yj�&��X�_�'�ɪ��)H��@T����f��#<�3=U���K��7CkIE0���&��D�6Y��#Li�y��<#U�z�	��}	�e6T7�����+��Mǿ�Y���F��`�Q�2�ӹ��R�j��K��"uE�B`�n��,ӫ�M$`|)�h��V�/���޻��ne�g�z�W5��V�"R� �j����u��s����(�/�e���s��|1�&���� �����%s���Z)���g\݅���G�`L�33t��&�AF�^N9��s�������92q�l[�1)UFDU��@)��
_p��E��ӄ���� �D9X�ѥ@�>r:��G�%�8 �M	d^����V�^��ː�Mx���t�V��:�V"�Q2���c�}����{��r���s��^'��k3@v>&��8Wl�<��K�e;�A'#M�Q��d0�D�mh0��Y�����0*�ҽ.�8MN� ��p$������4�H��^�ma�:jm�����4��-7��[�2W�W��"�%��N�G�!i`.��
:y~�B�W!mke�?8�+���J������Y�<^+�2�ǃa���v�PY��M�H�M�e��ٍ�@���N3I�#Ԏt ���$��[l��y������d)As�'6zh�/����6�"f{2Dn��m`�T�s�X0n?�am��T��&��{U3���l��!�㏠s�>G�E�Ys������7��\��h��D��^��
*�spe��"E���)�B�&0m�'��+hb�'e���'�����|�"�5�6��Ft�.�ؠ4,1oB�C�26Uav��s��&�Q' CnV�vQ~V����,OI�H�i�/���?`��,3����s(�s ��W��=�������|��U����0��7����i%���X�������Ko@J�"ed��\�&�!�ďU������@.�1VfQήT:���G�՜�U���GĶJ�L�x��"-���<ԫ�2���.�%��5���ʶ�cӞP���٥2���z�����.����#�E��R�3v�N� 0&�*~��*z��i�S��t��hΞ�y8��u�������!b!��ǉU�}sn��ajJ��V�:� _�yUoXQ�FH;��7:e��L���r1��H�r�� %n�fA�f�S�����9 �ͽ�84�52��?�����!�؉'�ԏ<\��V�>0H@?B]΄��dJ�:�Zј���W�j�tg�Z�wΐ��l���*~�'��/{�F�V��d���J��ݣ�%W�.��b�!}<Y�Oǐ��/���߯D�w�,�+�zi��y� xH�g8�~0�:3.�cIm�)߿�&������i9rc��xL�i_p:�h�q�P�k�+���R�j_�v���d��� �=*�o�,A����R�g�M̅�k8���Ԉb���+��ZBw�$A}� �d!w�����QY�/�,�����EM(�2j���ե`���<&p$_�7�����}����	#�:���R�]FVKR��r(����H����6�P��M�s�t��w�>�D���&�ޗ�e�'�,D\��W�t���c��K[�:�_��r�'sI�GL
��lvM�襴9#��Q|��B�Y���uI�r����0�Q �jew�l=}�m41��5r�r�%��̳y��W�ffa�#����M#=�џ�Y+�#R`R��{)���jZ�J�/��=&�]��N��{��s�
W\��K;R�lfV҄��q�{�a�g�钽�����9x.إf��;�č �����zW��wʉJ������J�Ӭ
���^%;�k�ۻ��y��9g�¼���'� 0�`j�
�L�;�l�]3d���\�?��QH��u�z��d�`�s��a^<����N�����'y��q�1:�:j�*��Eo��<G(6x_����!;�kz:��E'� 0	�W�	G8m>�c�G�6��2����р�Ė�S�a�1{M�~]����eK���xA��n�)�<�A<4$����ծm�3��PѨ�E��`��W�I�\cY��mM��S�����W�=�T����:W` 0���n���О�Y�0	?u�O�,U�k���yn�V@�Z�0ݥ'�8YP!���^�%��7��l��1�35 `�r+�;�xq���p�j�O�zh�J�Y�?)	�Bg�!
�}H��LLSB��g��g�����]�+�XA���"A��k#7�S�4t-M�em�3��Y�;<�2s�f��{9�33���s����F�w�[�wseiy�� ����+��k� �g��.�
��P�1�!q��;�aj09䊋�]�0��v�ŷ���`���V�CH���&��rz�@w�CZ�=��v�F�r���VEJ���)���)�E�R�(3W�]A�O^O�'�Q���d�.(M ���t�3�e���9�� ��V=������)jC�S��������W��Z߂�5_�<$�0��������,â�䠐���De^#l����#-�R2���^Mk9*���@�5��'\R���k�Ѭ�%.��-TŖ�G"%a&F�:�}�zt����]��2�p�w�?\8��C^�G�"+NdG��̣<*�	��Ul۪&��3�U
�/4��`.y R���c�) ��|$��aB�7��mx(���O�����M�MW8�����L�xW�U�
�jo�{�,���|'�v�>1k������2u�∕����I�L����M0���b���f3ܥ�ZDKf&<�g&_C�t��P��@K쇻���Y�ۉ��������|f�f1IiGD��H��i|'�-Ʃ��0`+? �eJ����;N����f/;����w�Z�9e\�V���@�k:f�Y��=����p+&m�r�hQ$���\uﺽs�q4�C\!q�v����9��l�uVc2�bc"����Ig�Dl47^�Y}.����	���]����!=��#9��{E�=�c3��^�ĥЇĪCF��ǋ�^�Bz�y�t��,�	'�j �]��sܤ9'�b`����E}��ތ�,�h��ܚ���n?e��xP޳�@�ul� z���/	����,�7��|���:B\�_�������a>O#I0El��o��)���~V;��	��z��W�7�������'rR��l��Cm�n����X�&ޢS�
*��'T��i�"P�����@���Y!W2�LU��q�������aO_
�YJӠ�&+�C�����'[��ڮ�/<�7�x ��PWU���KS��wVzf�σ�����H%�U}����O�o����xZ吡ס|��=���͐S�C$�a�l��,��"�@��ȅ3�j�㢈�u
ζ�����I�pG��T��٭�����h�b�;l��k {c��I���oɗ��қ`y�	����7�//ў�S��d���
p�#���61��7�	v8+\�SA��zF�!m"I��J��Vo�¢�U�+ÿ�U��,����I�D���P���q����0XY~Q�XU�y���Q@ЪE���oq��'ܚl� C)�q�쓳m���4�/}z�Q|Oȝ5E���a���� �X��ww�p�g�{�?�b�����>����(�7�;U�^��ޭu��5��dPxyN��wF�}�xf�.V�΃06�K��Q�庪.����$}j q�n���;��Tͪ�&�MxT�1_o�Ac�ğ����x�D��K�:������1%\�(a��mDw�>������8��(Y-���G�x6�il�A�D�]��`�:��i�%Z�hx�1��[pܭ�W�D�c��$2�l��Q�k������5#M`��_hX��!�J5��T�~�Q;��d�|���F��/��U9�g�7�� �k֟�@������?�+I�#�`�^k��eV:����(�>|��ȱ��_y&���i�7G�d������!3{�#�K�Q�Z�+�T쭕��#���8^P��%��Z�8/�5�W=��Z�xT�j�������Sȕd��Ų��C��7J���:x�VR@^�t�{��:XH�/�
�9g�L�A��[so(�LX_ܡ���7�p��evC�r��f�.���3���/��?�t�eK�4p:�}����}J�6�<9;�D3R�R��I�nf �������?[O�f���f@ø�CH��59�\���ʕΞůa����,H]�&�v�i���\'.��S�9��z��T=\ ���x5� ��!����qJ�!�ɇ�Lfa��1�'d�T۶���:8"�#�!f��t⾱�*��!q�^٢�{b�N��7���B�HN�Ө��O�J5�)���^S��L�����y�8�[��?�ƕ:�,-�P��5���z�Ď��kAa�#)���xv�1���R�+��t9e��Z���XP<f�/-�BI�����p����"9�����S��қ����xn�:0Fe��,���.9��O)z�P�Z����(+stg!�8ϸ^C�s���#�b>�ш4���w8:���o�)���cG�x=1�,T6�C�J�ϝ�d,W�;7�u&aO5��V��h��2*����U�7��6�ԗ_}Л�S��d�sٝ{����)H���P.V����$p�z�2���8:����n�&yo��v�0��2������]�;Q�<���k[+_�`c���؁ٽ+	�U�^��ۃ\h�]�b��J�bK��d�#-�?�!��\r�������?N:mW~����]~.g]�������`]��=oH�qYx�^hN���	cT,\\�A�T`i��`k��Zkk�β����?ȳy��'%\�����΢0LAG��_n#��� ��4�!�@��5R��ƽH�Bǖ�9�L(��c&�� ����;�9�+�":0>��$O��+cl���~�a��+���i2���aK�J�:c�?����,o獚����鉋<�:.����x�T��=�oH���"��ߩ���x����P$Mǝ�����[t%���Q)5�x����T@�Ki�VG���������*Ī
�{�����i�[�	7!��l
����݃C��5�]�De�����Q�ũ�s|�<��j�]��B��_�O��w���0o�z��X��PN���1��j��= sz�0�w{�z܎Q��/J���׬��ߪ~�fv��276�)�K����!I�8|x88J����H󑫭HC����B�>VC�a�{N�,�Z�tSsx'���d��BaI3sUf�16�e~A��ˢ�t:�I�2e/�(<YeFC��.�|���pVDü|��oK��E�t�
 �
��8-m9@7�ӱ���,1���ܹ�����L}GC:�AG�f��9�##}p�>p	і��@;�b悆|���w�00������y���]��o2ݎ�v��]ӻ7��&����^���5bYBp�Ȓ�	WE�$U��t&봠u,���SOS��zE)�ݲ�ԡy�q�<��wr�������i�I$��<9�=�	#���� : ��6:�j9(��d��w�
�7&��Y=D�y��Z@�d'J�|f���
B�t�O��#o���O?��z�u��a�X�(vbߖ��~9}���B�w�vVys*ϵ�H�Y"�`P�&��h?�2����&�t��G��%��#%U)�n�&L���Nˣ�����O��f̄P+�C��t��/��2�&B�<FAFCCf&)]u�癎	K$�L����x^�
"�� c��=h.6�f;��I�M� �y,���@�lu�h�ė��-!��1%��<⏤褭2�dŵH��=
��U�IsC p^�n"C�hȠ�#,+�_�X���^j_�%�^7�M��=��9��N$�r��\��;7�G	���V�%,�)�9�?����㸟Ȁ�ypd�*�k��L����*e.������
cjs<_be�?w
r�Ō����vg3�_���� ����Yo�y�Y_\��0M��5�фW*�8η�8��V$C"�E���[>����م�*Xe>/�v5��|�~2��7�0e�jBi߹z�kn��'1ǎ�,e��2\��6�'}�P���w0eX���.�=�z�i׾�q��e�� Ա��*�2�Iyb�k	B{u4�on��jn�ô��y��$���)5S��B �13������t)TD�O�*��Y BVB{�YL�{�7 ��	�p|����[�UT��I,�&��<�s���c|TVm��Q8zH��D�Q�V%����Wm��i��3����t��0ف�!	]�<�P/���[2��g�G�<QV(�jx�4ڤ��9)Il�6�/XT���l�6�*��r�q|U�pz�ŝ�	�o�}��|�� ��Ւ�c3�i���X-�w��$bP)���?�����w�L��̚G���jrW�yRP�	B����X�F��_����9�㾷��ҵ��������d��`��g.��ی�'������ }/����-}���3�ʼ�
W�-в�ی�ݤ�`�g��1(Iu��=3�?�6���k��_'~0��%�-�cf?�3}I�����v��B����Kո'n]�(A�0��2��Ԓ)�z;k	2�w�A+�8����[�U�Z�1uupm�	�ه�����3�-��+>Ǎ�smq�_�I����Hi��3�^e&뤠量O�y�Uk(uS�ĳ��r�{��u��*b
�r5�/ެ�2�S�[��>C�M��~����º|Q����.���}㮳Dޏ1�*7\qk�ڠ���)x��|�\&#"EX�Ke�<~�ӾZzE[o+;Z���X\3�˦Q�02�R��hr�Fs)�������	���T2���n
x����IJ���xMi��%�`A8��f�ȩO9�/�,1=IpڌN��U��LC�
f��t���H��hp�}�������M����B�O���DKoG�F��*0���R��ĝ[}��<̼�y��4�Ƥ��o?�Z�^;�8W~&H
j�\q�M�ۇgs�s"��JM}��'�3��?^+��D<�����LK;U�R�/��5����P�Čk�2�ح%�2�3��'��&�=��*M#p䁍/��[��k�ӏ�� �u��q9�չ�L���ģ�D�+1�`r1��������'�o�e$hoN�+KB�G���	� ���:BTsI�7o��xo�;��!���e�4��n��*xq�3�5N����e��q��J��6�:������ ��_a�o���؍��_c�O?q�������2��bʦ3;�d�z���h�-�euiuޞ���/�+��¢gh9�r��S,�e��Q�%�s<�����۞Y���ֿ��Κ���]�L����vV���ԿN��:�)���`F��K�Gj,"	��1�"1(��XOE��[4'��q��@�I�,��ÚU9�j�(C|�� ���Vkb�@�#l��wG�fe��V���'A�9&���7N�T�J���Զq5�N�W@9��1gP[]��,�#vGc��')nnt�Y5������e��EC�.E�������s�x;�Si���~q�g����&Xjݯ��O<ƫ(t�gz��*R�F�1��$}�L0��52s)mO��۷�#M(-�O5�8����7L>�C��a3��G�8�f�8Asԍ����`�`��ϙ����F�[�W]�x)�p�D{��7/�	�e:��,�~
����	�~�{���2	�q�^BD-���F�2���	���e���?�f.�.�e�ⲯn?��O�P�0��ت*��
HZ>X���y�S�����Z��B����]x��pŕ������"Jm�i���$j�J�Ou�|��U�pI����zPsRւ)��7�o���\O����8޿�`�(��'�R.CW�.qo�u��B_���ňܣC�]��0Y�n8U���d��Y{a�����4�:�.m�p��k�{�e5��%��!Ї�}�������=F���~F��;�k>�[�r0��ƤX�4��̒0�p�OHQ�~J�v�o��X+y��E�pt��|#Ǆ!$Q�`D��u��XʻI��f~�<��@Zk���jt/@�8��Z~-zB�	h^�rN7�M�(Q}�c�������n�?�S 4�/��؛��r�>��lr�)Zd�V&���:wmfڭ"|��g��C����F޼�bZ=ۉ"7�$�ʺ��:��,��i�/o	3�R(���	�8��W�@��0X!�=!Z�g �>2���~���N����fm�r{�*Q����Dvӏp�%��9�)n�='�q�.�k���d8�g��^~8�����ܙ�U�E�r����c��KT,ohK���jUZ�~��@/��dە�`��
���s�Ǝ�!.	����pОM���1��`&p��[��%N����˔ݡ�Fe�� X���T��	- _4qU��R�ua�^�E�s�l��l	����m�=����t=M8Z@d9G��O���K��O��������?1$�S�/��Nbج4˂h+8U���b��d;�Z���@�D��н��H�����}�ޤbxeWxNi�^:�>�}�G�q�=C�Y���W��QN}��n8��[~�YSoɠ�c�;����O��8dxm��ty]�d��ʗ0`|�7,�A���d�O�����-y}�!� r����RoҲ�v����Q�8ɝR��8�l3qDў�T4{;���[I�ҳ�C��z�}�m[���a�7Ν�%�J��%��X1x��(�	�͠�%��H��zB�"�q�=��	����u���(����x�k���U�sb�'ߥ�����/gRrJ�[�X�`�'S�[�5J�:)!~��z�ÿ ��ȩ}I1�b>�G�E2�w5���_�b���j�{�����	�P�z�$`�%����B N�K8��������ΐ��7���4��.�2��x�*V�7 �D�dwI�k�~so	g��VN�0~����B��S���S ��QN�*VZ����1��b��[���H�b*�R�s5f��e�.���H?��j�"���J��#N���a|[*�c�zR&�J��٨�<k�1��抌�:��!̘Ln��`��4��i^���<�]:8}P<ڄtb�a�4^BrZ��gb������������EY����b�>ԏ��E�p�`��!�5)Su켰'x�a������{��L��'{n�/�'�s2��W�؇�e�
SY�.R�;���4h�Y�����a|#GU�&���;����F��xpi�H��2"��$'�hS�/������oD����z�6��vU0)f�~
>DX�C��?�]j�^NB�at�{�xŶd��05_�`�Jͅ\�JPү�P� kC�]���6�5�7%�����(��?�E3��L��~��4YST���/> 9i�[��vb�Z��%�� �d�[4���@����#�G� ̑�
ÃN�7&=F����ܓ���3�!�\S�N);������ ��w��`-}~pǫB��L8�7��ض�����(j����v�����5�eV,EI���A-�`Q�|�Q.�7_�I��Џ7��%�x/3�P����46�̗�L@M�b�~�vv�l�-M���d�ZcB� �"R��\���$j4/J~@왇m'eV�D�e��S��aag�]���I��G�ҡU�����=Q%r^��n�GV�������| b���B�&�"��mT���w$�q��`�.v`�+�PhoI&��1]k���IX����g<L���u��1S��1����O��{<��j��:�����oy2��ͱJ���011m.,�\0o��v�aA�?�~��MP&~H�-�H
����7tK��6�9j_HiHe�R�*=��ngo�5�=�{By�n|\D4�1�|�1W�f�k.�	�P4�\��}p���NoѮ���>Np'(n?�^	հ�����B�4O[��^�n9�c�,t:��q�L�h{	�@��)2U�����/�Ƞ��xy�C_�$�<F�߳����kI�BTM�K���AK;�d�S�Wp�a�A���w����aRG�t�&������
v��J��E���s���=z�.�2����#�L��r����غ���.��T��CuE̙#A�g{��͝K���0��[^�g��햒��]��b����S�-�.B@�@�V��	k�/1�j�z�����Aɞ�!(����"�/ �P~y�r[ȚR^���dҁ��AV��hS�����;�h5?g�A�ŝ����wUϚs��� |�F�[����:Oِ�P���� ��:O·��O�x�#��!{M 
x�H��vSm�2�F49���i�C�G�w�SҌb���n���np�b{��'��P�5w�P;J��珖�����Rt�rh(ѱz�*��S�a%���ED�m !TN&PX�B����e����}s������Ȗ��~V�	$R���p&�K�5cUT6T]�kAW��~�4��2�p07��h/�?��s+�U�#~���z�rP���N����J+�� Z!�M3��~��2>�P먴H�A���Ѫ���2�k���Q�G��	�Q�Tn�E,�*vzY��L�w��!ֻ�m�=s�XX�1�A�\�[��[V.||���&��a�eW���P�P3�s�0icߥn���(��c?��D�k
U`1�簧�-�̽�Z/'��0sW��k#ar`�����CS3fjL��ap̺�^/KĶ��޿�ycg��rE;l��Ps���3<K+�0�:5M�Z�iG�ȵ�g�^���;h�b�������b��\�&U����R�!>�eT�RnJ����X��VO9�H��pUWs�eL��q��D��=YU�l�Y<�-��opު~E�OD7�1(��\6l���L��.�[c�8.'����k -��Q��ÖE��so��$�����7+��|�\T�������ց�"�+����]%�'��`ւ�r�lryKנ���^��'����^>�JA�H����˥e5s�����'�ٴ��l5�e&���\�e0���B�Zr���"����~I�����1K_q������������.u�0�i�鉉3�� ��EW݉j�{j��i�m5��}!mG6[.-Z3��
�{+��/sH{�f^))iq.~S�B��[^�n��I��䮜x52�H�0�ue��o��Db���J���Z;�:�a��ݤ0aa���ف*�G�U�h�/��*�/׋�@Q*%B)z%��6�#��P���9Vi{��Rd`��R�����C�C:9���-���>�r�:z޵9��L*4�Կ�R�h��p2��T�]M�C�e�1<���FVY�o����t��E��qf�!
�k�0 BL�ЋW������+���y�M������g��F�G�_n(���w1����P��L��'�yr��R�yf�(���sYHcV9�Ca��U&`�]B��_! ;9VLg3�e���k���1 eO���.`~'�)�
�-�d-����a�8�OH�}	_C�i��J�GPz!.4���<&�J��/���rpF�F�L0�9���t�gqK���1�s�kכ}Eo�\g�v�t���&� l���d� V��4N����$����PgP���;N~.b�D׈4cۀH�v$E�����.a(�1���<���6�~r
����U��Z
�� ����s5�����#��ݞ�n�y1*M��~�#�&�q�u�pO�Ǐ/�eGi���O��F��1��K&�X�~��fa窱���٫+b9�aD�%j�TUX<����Q���*�A�����՟<#�9�
�C��{Ԏ�W2V(^aN�W�B��qsz���W�@�U0|��R��F�I�LnP�2AIh�	�l�j�ȷ���!��k�F�paA�b@�	��(�O�Ca$bQ����U0��B����}z��0�Լ�����KB���w��X����Tr�u���ˆ�|�Q(�?1�KYU1D���@��1�}��}��䙳��ª�DI��;�m�o��5������_��^�g�Eݱմ��KyD�#$�]��_��?a4�l��3��p��y����>֗�E��v~�(Gg3�-<�{���]C�>�Yn9���
)�j��1��'RdV	B�V30-���[�!�1�<���`�
̃y(��������$7��\���A	⇸M~�D�D~y5�b�� �*#D�re�o�P��kR�ǜ��G�����66_�Y�O�S��X5��wA������y#��w�Q؞�\�Lal�0;VYs%�n{mMbrqPn���h��5�.Z�x�F�$>ޡ�̦\f5���g:���Q6�+�s��`^3�A�-K���f�*��4ӣ�"(GR�B�+���}4I�	�z~�&�Kz���>����Y�b���r9�GI|�a��]ށ����v�l&~�&b9�//���e 0�����Y`��^�ƃ���L�p+҈9p��,jr�|�J�U����i(e�L5N05����|��J��·kQQȝl38��ud	�ʂ��s�LX���VO'��Q����� ��r�gKP�M8�s-׊�Qn�X���&�o�Y�d��~0�9�sG��G�yf޸�����sk]=��F�@�]��j�1�����f��C.��CO��ܝt��T)M��?9�����k�L��{gE��F�A�I�q8%n������	:�Av�-K�Q'�32�VZ����V��!,ͬF�!��O�B\ ��_s�O��D�a{*��Z�<���H9����,�Z���*R�|�M�(:�����R3�N�x� x�{ 5�1�J{Fʺ^�SWI}���R�t����Y;#��\��k3�x���"�:�,�u�D��s^��n�Q�&�P�(��ϳ����B�F��b`=|>�r��2�(��Zi9ew������g
s�.� 6�@I������-	[���`T�ۚ�a��p���̴Pm��%č�#�[I�_�d�}�'������koD!�l
�]rB�[�����Q� �P<#�\�r��U(,�[6Ć�`r'���gR]�4�,zJ��Ɍ���c(�O�����V�ػ�u��c�c��E<o�<�#�ӥ�	W�$�&%b�b���&=V��EO;��ߚMG�7����8IW����!!]�A�]�8ja�������4}b�i��NR�4
��p5IiB�#��F�%���jk�Y%�A��V\�T_�2S���5)��i�&��J�=���''Դ�[� 4���Z�t
�^Fêdr�X�Hn������Sb�7.�E��~�01��o��������!}�?͍�ZK`�]5�>�9kէa�o��i�WjZF�A�/XD�-���]���$�+�f���'����Ƭ���0y�4�6���4`�q���Ad�R~e��Q*=�&��Pe�?�.���W���*�o���nQ�.r�
hC���3��81�q9�Cr��;��L,�㕂�"h3C_%�c!O���KF����e�8�6��ܻ���_}1�߅��y�,h̯D�N� �)���4d!���-��*��ʹ�#F��Ӱ�񫔠(���2깮ϣ�#����$����8���+rI �0��c��n�,�-��w0��"���I�J���o��:&)F�D�E��jO�H9�:�?�n�]#�,���d�9��T1�d#��g<K�2x�NU�C7i��.�ϲ�a���l��P��T�K%o��W���ߞ�*�\0��Q�]g4a[M�	ؓe��/C����+�순:�yƓ� �L���&���Z�&�$�>n�H�i�P��K����n�r�B�I�}�����Ǜ�5�JWȏZ�MĮ_f�ԓ���7D��8��:�~9�,�|Ic=�Ó�?�r�Rޯ&�w�0��|�WZn�6��jȉ��#��Z-1dժb��5]�&o��?�w.�	b��D����tPz"���w�u>B�Lp� "mI�{f'�ZD�0�!/f�$1�Q�Y��Ʊ��1V�����q�zz��{�+.@$�aw#��,��ͮ���(W^�^��{�%���ج�e����ƙa�)9+�y����	4Cw�y�Y�![�d��`R�K��c�>���FC�@l��
-���2��xz��`l;f���j�t�2�Ak��{������  �nY��Ȝf��#6D(��xRڭvۿ%��
���4N�؊ad� �i�
}�˖_��F��<���`� �k#��G��0[9���2��,���n�s{z� �W�c�H�U��«�߽
�y�Y%����?�R�"��N6U#��d+���@�B��#>�a)1�̤�J3�V���ObB/_a��N�}��6%����,��\Ė�Y���`©+B#O�M5;G��ϼ.D�)��1d�<��Gj:[W,��Y��	�q���T���Y~Į�~�`���mn�$��֛S(��a�r=&I����0ҩP1U`
G`���w�[�;ab[H#	�3��iC^�)w���E*V.�_p��{E�r�<B�f�C|,=P̃#'�=M�Y$Jm����}���"���
{C�	Ht�~�I�z�H��Y:��u�ig,_;>�3�����7��pĵ��n=�*��?�l:c�	�9�1'�Ș�޽z˛��V�&����R��H�W$,�]������y��Sq44ct���D���к��u4X@fw���$4�o���� �C*3
�=ڊ� ;�)!���0�!�4_@I�ՅV�G�!��^Mr��AWSB�l˰],���0����cA�V��p�t�?l ��p��iY Q:=7O2��4.�����/Q�y{EPi�����nɆR�<*��a�LkaMGR��֞��H���"<]7���}���]/��X���H<����Ҕ��!j�J�:�l��Y����^c�J�u���zbM�|�%���������e�b7۱����������ێT*�Vx	�c��~���w�-dXN=�b��E�����Di��݊^��r���_O	Ԯ*Av�j,٧���{Lwp�y����%n�E�j�S�I+��2o��Ƃ���L ��6�1��B:�J��Tr~���N�J���b�W�֦��`˧��dm�"�8�����Y�7�X���"'s��j�a�R�mSI�Z=�65��0�P���j�LH��4�`!�3��ӅƱâYq"� 軅���;s^���X�(�^Ԕq�p�x<�Z(|�(8o�S����G��Dl1H�2�*��Z��Bl�lf� L���3`�)�y��^�Ӿn���xe������aLJdg���˚�-Ke����Ҧ�=�P|9q��8���[���YQ�PpM,<p�J��Q�k�_�Q����x���b�c@��A⋉H�JfGxd��-ܻ|���)ޑ[P�_1��g%�0"�����I�ɺ�H��C�$��G6KV��A����'�@ ��0f�R5�RPo[�ee^�m�4@)OI�V�.ĞIO-��;f���[�?�����{��֬��C��^
��~�"~�00�+����8�{-i�=�DNt�I���!�cqT�Gq��� ��Ԉ����-ߚ^��n��T��ޠ�;8ə, 0�����F��ct��u����ʸeq�_ʔ�*�U�i`A�!?�v�(49���� �S�"�c?O
W��1��]4Qd��d�P�ÒW�q��(���𠪐����Q��bT4X�_�W���7Z�˔���rS/�ѕ|%�-�e�q�����+X�M��x�y�a���Q�]3��m�ىj����k��XO�gJQ��f?�dχ���UG&��D[������QZ}� �'��?έ&OX9��.Fc>1�Yp�۷H|+�<'?C%�Q�w4�N�-��B�YT899��6S���_ҵ�j�Sľ��� zw�Zn+�L�.T��k�4y�%�9��ߏ���=����ώ�Ur~'��7K���á8��qSH��p�_� �����$]�?��?�hi���F�XT�E�~^�	\v�0�G�yݐ�6$�+# ��6"�@��]+�Y?̑RԖ	�U��wx�=?|����cy]��Ϳ£y�)�B��J�~�S�s2��Vٚ��F�cpx���*�6�zy�����M��8) �Q�hw��5�y���Pt=��B�b�(WJ����I�N�LC=�y(��)'�M�u��	=L��C�y�$/x�=�V�	r�=V6ճ�(	�DJ7�Qߖׯ|𝼉RzT��D�ܰ��y?�m1�N]}*��f�=��J�T��d��{ɴ��F�p�'�����mqy~H�X���
��5��o+Dm�}��Hi(!��A��xx�:*�'�������r�@*\�pd��/`�8��v�?bg)���
�8u~\x@-��U9X�L��H��"����ms��
��x+��P �7���t�(K��\�����
�KL�1c�Rٌ�;짭A���!�F�A�u���^b�34uw� ���A��cW�ajv�6/Ƅ[�Gp<ɶ*�w�ؤ���_�R����9��һ�|܁�s���(�#㢺m!B�l���G��`�J�vC�y����x����Z�L�om�_^�|^�Ǧ�4SC@����f��X6�X�L�~g�Dg��! ���8�v�7�Š��%"?$��_'C12��KP#���~Θ�_1B�`�+��yL��m{V{��Ȼ0���_I�W޾�P�֪�U���Ǽ���4��}NL��5v����.�r`�d<�D��Z���ʢ3��R�T�+�5�E��P��F�����V��j�(RG�<�4JQ��z��W����2���^�S�xvAs����{��7G䳮�����q��2��p�o�(9Ŕ^����T�+�����ފљ�Χ@�-��Hn���`�$�������3H���� Y:0�sk���4]0"�}��q,�*u�-�-X�:�P�
=�<�C��y��,_�|����̥F�0�[���~�b�� =%%���Y8_Yݐ3*��O��O�G��O5ek`u.6q�9�b�*=�o���$�OU��z!OjW'oW/��d��>�Ք��KxkگY��)�:��Ț� �zʛ�ȉ���EC�G� �!_6��0ݨ���w)�m �|��E�4�Y��=6�@BL�4My���u��L������3����08�3ݩG�xmzϋ�;��e�7�=�E���t~�E�{�%-�+�-�B2D�d~U� z���4�Lf��$�_�Y#�<Cco�Tycő!�p������d���h̉��앐 t�p�f�鑦N��z+jȦ4/��[E�T4w /�mq�^#C����qGiJ�
�����B�'����-S�{�4�̾�Ce��Up�ڙ �7bN�Ǳp�^���Ny��C�@�~�BpFD�[ɇx�s����l����o����VM^�*�R4�7o2'����f�~�zXB��d.��~ �C���j���Z�(�DB�3���ͥK�D���)-<��}ˇ��b&ôq�����}p	�R��x��N2KE(���G�F��j�y�H�g�0 �I����a�I�'�	Yea�?�$^t����5�d��$�r���k�S�ʆ��2葂~I>b�;f��
0��v>^4ըlB�<&�FJ���}BВ�x�m�1:�ѧ�6��Wk=^�X&��-+��?3�nR�7��6c��搜[ޢjZ;��R.!��ށdvρ����rԌҍ�:�8���6�������=_u`/I������u��3t���A�/>ִ�>��qaf�3���ʮ¬Z�F�Kڝ��ć���B	��J�i>�y�
��&�l �'��@f���q�(*�X �$;�"��¥���*�F��t���{�F�Ze *���������g���R�vFȘsH�&W�K���q��h%�f�՝���ez>|6}Id6عCy߁���-m����Iϲ�dx�Ǐ9�Q�̂Oy䠕(!��˴k,zT־�"g7��S��Wý����I�;O�Jo�p� ��@�[���#�5Ji�����_���[��������^8~��>���"s�S�!♪����7�2|K�|_�Q�QJp�����yeR/�`����s ���8@�sz�|b��uH"6�gl�b���z.��ǭ���������_R2����w����-��!S�>�q�~�y?4I�^�#|�1��|��K��Z���s�@��|KhBM���5��?2�^��Iq��� D�쫼�����{����F�Vȵ��V��a ]��� }�m6����I�$�M'�����Ű<P�!b[IV��B{�d�(]f]������Z:�t���Jn�_NBWC.�L�'b,X���b��������ʅc\m@�֢��pȺH ?h���J����Cn	p�>*��a���ɺE��ǂr�Bo���E��򔟪��Z]Z��Ĺ����W[աT�yS �@��-��n�H��ӿG� ���P��^����cR�;4|�7܈���:#�J�9-���(~;��1P�1����>)%�!�^}����hPY�i���e��H�ϛ;8P��x&���W��JY��i����<��{7O�/��b?f��E;S��]{��bo����^<��.7&u�gߒ�
w"�Aw.H��(��<A��ݿ%��-1��M����
����U��b�w���4�a��Q��iP 4tH�`ˊ��Z�*kD��i�~i��V޿ `7+D<�,�tC�V|�z1�)�C�m���� ��~ݛ�������/R�i�����^6�2�|���/��fZ�;�#<,3Ɖ�М�Ѩ�=1Ii@kW��k	?X���as�^ozL���y2���$y������dJ\30\W��	�ć/_;mA�*�P�Vz
g�q+����t��e��q�#'
Vb9�z^�r<�s�K�`y,oA�(ژ�hV���&-�h �a�e/D��ʱ丟��mxi#	�t�q�b
�����)].)��0�@ �G���U5���5>7_S�f��λ8��7���c#G��Ű&�u	B��6�;T�D��>��K��8�:]90#�IX9y��T���Qk�q �S�ڙ��(8���+m��}'�@Y�UF�I����o��x�vD�0�Ld��z���-�� <eGzg)�0! P���6�2ˤ��Ǧʬ���O\�fh��	
n!@�U+Gi�޽����o'�,H?�£�~?���-,�=�o~dy袤݊��ЂžfR���PK�PJ��ӢH!`Ћ���IAn5�*|����9́�R�Ȓe&�����]�OS��u��D���T
^�~�[?i���Ո�(�_ �^l�Z�w��L+Xna�� f������h݀E�!�l^��s�����H#¤F�!x��W����,�-��21��}�k�w�ʹb
tF0{Ҵ�Z��Q�a$�󀖪v��l6��J/ �pxnF��tW�;o�{2팏�j?
������L�;�Q ������aڄ�VȠ��sW���fL|۲��7�E�
���H�Q���a��'�����GG(	 ���vbH�S�%2]���(Q��O���r	���U��f�9���d� ��������|�����;x8hRA�p���c[��G�8;h��`�Bz<��a�$��ʂl�l]�����.��8�6W������Ja��R7�!fn_ب���k{��>�Av��(�}Q��u���J�e9�D���v����`�&G?"b�CW$�]��Z�[���3�:OX��"��~�Ll���Mm��!V.G�����~��s���t�H��B?����T�81p���킕���W�t��-#��.�إ�1��AJ'P5^ű�}Xi;���'.w��^���3$|��?��x���۠����
�?M�ۭ"�y������� +p  ��k�q
��shḲ�M�/r��lR3.7��H�5�E���G]��B?4-��f:��֪�9��|�C���L	�ݙ���rkF�H��X�<�w�n�Y��gR���9YW��M���RjW�^�=f�����C������D��up��C_+���F9)U��(�)���7�g(��P�q����U��!�V�հ�R`7O9��T�,���i�6��`ͪ��X���<�/��x��@zВ�~�۝��_�3�/��]�>��G������֙}$���w!��c��<�J�۹WE�g"�Tx�N݈��,�5֗��u�<A�j���p{�.8w����F*2����:.�� v�������S�LZ�y��\�����	9�M.�=l��7��&ni��ܐx�L	S��Tl�}mkv�z�m�s��,�nlx})�R.�l0N�HV�tm�?��e����疙��O织�8k>������+@� P�(d��6�g��?]`�Z�%��C�����F�5s�䆙�d8�"��Ȉ�� 1�ձ�	'�{\����"�%E^n�   %�F5͌���J̔"� ��GQ�F�Ji�o��e�欫���4���~ㅬۼax �������@�;!� ^�6���U��6J}@�$�I��x�%FW]��@�9]��_Ĕԛj+�8�ё:u�u#q�1>@B�1�R; �����v^MS`;�����on�HFw��#��gA��}a;��9��c|�m����τ�������N�3��`��f�@��W��k���?,�vk>6��re&��V(��Y�^8�G�^�R�%�I'��)�� Ԟ<�i��@���M'��b)�Wz�0f�h�׫������o&ѫ9��X��Ou�GpR����
��b��q�SV��T� Q�'�P=-�	�ˌ@P��zF�<b�LQ^S��BPu�����TQm������,�������/��g!Y����]�t�M0�?w��!�tI�(L�_��/]��t������~Ab<`��.>��a�do7O�����|��	���׺��ՠl�G���o�CfV��e�T���	>M��#���K���狤��#t�C�1$P�ގ*����ǗOBxf���i�����Rf�KQэ��;4�7[jW���O�k�
9Z�0Sv�쐸����<t+��j�)�	��J���Y����	�W0�����O����5�+�!o���i�&\D��h
1�PQ�g�l�9��/u6W���|9V��{�^fZC� �*�����5��﹬@oW�GE�z��
�����3خo5q�9䲔�NBs'�Bxik�_����)���sn�����Q�jW���_ޭn"� ���}d �x*p��i�V����P"L����2�o�L��|w��E�%p��B�xE���r���<��'�3�2;��]�m�+�O16��ŀ`����q��%Ĭ 0��}����)y�LBӢ�{��ؚ���ni��	x��d$X���g7]���!3��u�_G�7�7��.[�b�;�KB��9����"��	 H�M[͑NY�y��y~�Ư��&?��G;6Qp7H�����7R (�-���}�T]��A���9%p���s-�L��黮�'3`���H�����110k�_|�x�Mߖm�%�[w�k�ΒQ7z����m��0��rř�Eˋ`������L��~U��w��Ʉ�A����$Q�Y�"���R�[с��VV�^}�q�DZ�(�06��V<�=r��S2��qn�|k�F�-$���3��b��F?D�)�6��Ylx�D�e�'NzAx�مʺ*z5��%�����	B���M0�L���]�Iy L�<�x�T������l�'w&e�
li���-7�m.�f�T��)�;�%�L㢟��W~�m��,
֒�S�R�ɓ�;�m#A���]�����&�:=6���C
�:�{��>L�қq��!�%:�h$��>����ᶇ	{�ƴH�z��ZT,\L �7�i�� ���ǯ@%Y����vx�C\`W�_��M����.&�y�����C*��W΄v���3�׭��$�'3Iw<	Ję=E:3�jA
��.����#6>���@N��#y'��ܐ����Dn(ul�7'*Q�C]����`Bĸ"=�=�*�.I;5iK4[M`����0��|`��#�\\E<Q���j���7q����	��s��ba�@7��G뒭�}�g��g�{���(�b��Έل~�^�1�`&��w��MF��dF�Z�|�oG�8�1����Y]-^���a��d3���;�	����%ru� ���.��9l����ŕO�	�j����V
�hw��W�y=�<�C�Zn+ܗm$b#�O���8Ê���%�"%��%�Ա�?A|`��F؁�����ƤX�O�V!ߢĳU��u�ꕮ�:xh�CPGBl(�:��l�.�U@%�FbZF(���5:fB��/}#��>�i�L,��#��b���ic�5,5J�9���wc��K�e�H�O[���g}:�� ��`:BK���&�q��m�!F{��2�`� �&�1x���!L�k��>���9���(���X��b��׷����l��x#���O�*�ƞ8�tcLq�!�}����/��et5Q���)8�|�V���?5SV4�d�r)�l���t����X����o�����P4$����8��q6�~.���6M�r�em�)	j�(��K�w�K�dX��,��!3
���߹����'��{�k�q�M�Ӈx��P�Xfֺ���C����T����Xw��}��K��m���з�&˺��2O��"�4)��w]���^jj��w��N��,��n ����^�Ϭ}	�,�Y���ز��2��W��/�M�,֩�;��{K��\>�K.~�-ׄ8T�L�V�	J�Q	�Bn��W^^��ݹ$Aԯ��tb��D�ŵ>\��ᢚM��T�Zq˔�{:���s�4Ŗ�-�¶����l��bѣ�3��������׆��X�v�ڌ0�V^)���K�[�P^+�������B��ۇgĮh��N���֠z& �����u*cJ#��PX�d;�م�;�d��H}�v��oa���bT}}�%���݌���1._*b�uy/�^�l7_�[ODĕ�y`�����>��eٮ���&���'1��/��aY��b#sM4	��Bqv���~8it�?��?�BZ2i���Hd��I����*���`ox��������K�A�d�ΰ��*��,�P��X�՝[:��O��Ui�hd'�0s&�@m�y��,�,�\)��7�ґ�dx$G��H�>�8��E��}�x����*��
�K���E���cB�
K-l�,%,�UK%��sx��.LU{���O���wѩ:FЄ�fa�����C����l_%�0�I$�6pҨ~#a`y%�s�4���Z�ٖw~v@%����!�(ܓ���҄����ج�񆴭�5n#5���!��f�o��L}������v��U/�倐�yX�2�6"��n��}�k�*k!���jq��C��h�/[�n����x�C���Q�/�W��2�&�:�av��s�`���@�8|��"��i��l�e�M�L������
���T���KF̋�M�ua��d/����B�f8�����ɏ��u�ގ�ɰ�AE���m������������"����Ȕ��jٱ�$�O	�j1�,EA?O@sO�:�����N����#h ��-����*=M{k���<����Dϧg2��} I,��6��.��Ws��<2�'nTY�`anr3@����ktdd$y}��.Fm�!Q�4�����5)=Be"6Ȟ�,�sX��'b=B�������9J�.�N '��Vf~��K��4��r�EXڸiOW�D�(�g�!���w�y#�9RYC������@so[��V. ?���T��Ϊ"�p���1Ath�������vU=��h�6�Ի��n����*�Dnj]�ځC�=�x���7�`�UR>�m����DM�,�\5=�K��jQa�p���d�?�ː�絔L�vIK���#YȽ��&5V�(bP�}�Q��}�g'�xn��a�X;��-���
ID�����ʆ��X
�?���"�Cr���a����uh@	M����_����������|p�3�/��RI(~��j�N8�"l�w�2߈�����R�Gb]��dBL+V�]�7�EAFrP�$��\*��<*Vh|�������Ϟ���2m�2F�fG�Ц�q6K%�õ���4O�@I7�V����hg�<M��s�2?�%��� ��e*���a��V�I�1�Z��q1̙�9�2kD��BY����i�<�n�����8:q	����u�j���lig�����t(�Tu�Rb��:�ry{�>oq��)7oO%і.��+Z�B��}����O���B��D��k�<.�eOP�N~��_�lc��Y�xIG\/���$ǔ��h��V�?kQJn*�|�%;�5z��Jl&�P��x���O�`o5,��(��ڈ)�Ep�,����|��A+���R�b��,A�w��S$ة|��������7�l�����g�]�-7����c�F�<�y|�d!�;�:}��bQ�7�aO L��,|ũv��A��������N��ϝ�쿄?��mB�*S�`3Ǔ��~�U�gH��0��Er�U��@?�a6l+�K"����x�yٟ(�z"� �Ҹ&,��y�Ϲ'�,N��:|�_똫�~�-��[���[4p��r��ˈ~H�E��e�M5�7�PK�ϔ��6�R�uu��}���Y,޸���Ki �6��Y��U+i��s��WV�:,fB�@�M�>���1��^��4����pu��_�	�d�X��:C/���ԔF�˸� �����_3e�0D����ͬ!hu�v�wA�3A�Sӭ�5r"���+w���чś���s�	L%M�{����x���X� 	�P��6@6��:���l���)*�~�)'�V~+A��򏁥�Fc�|n�+�_�/���I����d �¦�|I���W�+z����fU� �i�C�Ya0��ש���f�2�F|��)z̢��m��j��wy�h��]d��$`�<��9��k�K���ڣpy�'���U J-U����n����m�fӛE�Q��L��g��{C�������-<�{���`~%��11�][�(�YLc��ձq(]���Ȧ�x.f��U��Ī[d�$���ٸ���/�gFg���(�$A�,����`����嫀�����b��ƌ��B^�\n��V�4��A�=��:�q�d���G���Y�1��UU�1��5Y�9?7�w���� ��|�9$�s���h)� C}'�����ſ�eF�[=:��#�,b�?�ggo���)`���ľ���D�6�{'l� ���Vp�������p<ȳ�'#ȱ��L��`w�����(�
؂����w.71��~S%������[
ψR2��t%m��S��}p>I�T���3Q]+#��
B� �̟\�	Mz��k3�r�l]�ԇ��@$9���/�lu���l�l�˗#RAcO_l�ZMmY��h��9ؔ 9��v3XU�u*��*�+�e���>�5)���i�}5q�r�A=�������IH������x%�Ρ�i'��ac��ê.ߓ�]S�H��p� �/ҿ�qy6;�8�ЉM�W��:�CK˷g�8��L<q"&�:�}���.�<zqh"s}[:�����^O'�Z	������|&��#i�� Q4@���J�͡��Ӻ.�!I}q��Q�1�e����$��C��ُ�\v�Հ�B������' ^j���!�����l/��fxR��?k��V)�K�ث��K�˗?��.w����/|)5J@:i�21���<�� ����$���5wMȉ��x:Ů'-y7�zY��M:��4���b\�I(4iL�ox��9�&�֪8�́����F��\�s�y	��E���Nb�+w��Vx�
��Z����
�(�$��@��!%��?��P���(ࢄ��l}/��x��Pc��aL���(Cޏ�z?����l1D�4���D����e�c�Q�C]��H�\�������HL��]#ϖ�G�+*��_� �]>J`���*ށ1W㨊�Wi	��_��s@�<(-���KNhp�u}+퐓(��{�3<�ʹQ*(��=V4Lҽ�]qo�+'
�lHH8��,c(��q�� Q
o��+9E���A���a��C3�ٸ;��j��	'�^`��XE��t� �{�����a#?��x�\����}Pye-�ɮ�L�����)��A�N�F�*47A��.�g�״Ε� F#�[�ӡ`7���]\�ɕ9��y[��I+�/)l��,�%�a8����Q�����T_e/=!Qк[�#
��ɛ�aa�uz�X^<��� �����cm�l�(��@��3�`A�=����e�1��A��[o=L�m�6K�f��f-���J��nr�ej1]�ᓿ}b���d|n��*��A��&�n4A��+$#�L��55���}jy|�Aj[Ć�mj�H��(�V�^G.}�L��3l�Ņ_�sv��Bn���w)I'>��)�YY�����XGL kV�b�c�mH�Ѷ"lI�;��m���w�&��+𽵁��Z�ˍo����9�����+d���PU���z�cB� :�\N��IR(&�]����3��3�PN�7�%E�e���6�S�6Bxx��>��K�^��
�b�1c�#�]�*i�&��>-\�*o1ɋ@�j�"e�x�=������ÌΌ�{����a��x�{����|�0���P#]+�A�=V�B d�{久��hn��8�>~Mi�ǅJ��}	� �q�A-ns���>MoTݲ�)�W����a.ae1U�=>���9Cq�m��o�@�<��x�o}��m׿y� A0;�2K�
���ϔ�w��N��(�8����`�#1?�����7N�|���(�mfG9yy$�Eh|T���V�omt֫ ��>�B�������r\6��L�[�W�It����
��)r,1���7�Hj6k�r/D�k�Ѡ+UA�����������u��n|D|�������R=��O-�:R�3����a"�L�(`Rғ�~���ا]&�B,�Ԃ#�4z/���\�$�	� }A���,���B�f��+N�>�A�@Hds ��M;��d��|"Je����`�+�w�=�FEp{��'O8A���t�?T�"P��*s�Ă=�<��d8Ǽ�;c��t�K���?m��T�K.�8�S��3�asdLI:���( �[�ke�k�0nc�7�;���M�)9����+�U9�"�*f�Z'�i�Z��f�'�T�.�(Uk~'��,b)�e�R���ò)���ז9f�ؽ��e���'ri���e�>y��V^d#���/����;�!�Q��,�97[��;q������$����u��g�9{}Y�nZCD�_��襎{��&���mX:{��+�W܌d���h�3 -0��A^ a=��rh�3�� W^yTA����p��f�?�J�T��z�y�������ž�씔P�G�+L7��[{����8���n��.�ɨ�n,���r���u���tN�:1�;s�$����f�Z��x=�%j���%�͍R�
����.0:����Lс��%��mi��߆�J[p.>�8a��#oQo�t\IQ���x-�k�׽7l���ä5L�+�sD|����҉0� f�.3*5T&�?/^���p�����J&�v0ti�ȸ�~~�&g�PmTg�`j��!�H�5���3Y"�͡��'Dּ�;@�����5RdK��(�{�ᰃ0�c��ʭfV!�>fpi��媟҈��S�}��F4o��f�8<�mb �O��6fl�| �\g� �m�o�:cE���v�3�Yj��Z��rd}]�OA�{7"�r���Az>y�<���rC�$�.I�l|���g�ln?������"�������}LF�H/�EZj���(�ǈ�v'M���{6�;4��߈�٪��"ѱ�+�๒cE���3m��m�/���Z��:ֶ��MX:��x{{��-Fw��X���O]5}�S��,��h]=���iw����k�����:�ѷ��e0/3���f?F��)�^���8������L%���*b"�˒+�7S���z(�	�W�|����ȷL3��W��:�/�ǂ2������Ʊp�/r0��1�I�8Oћ���٢]L��3�%������ԍ�bw}�@�l���{H���p��n򏴄�K��=��OI�w�dFП�_=�t���i�X�k�]��Uу6nk~�\&;�!d��cj����d�@(��/�Gɵ��)����wT7j�(�A=�U��sfo
��N�Y��G��4���ei@Ļr�zs���R��0��\�.�N����j��~%�r�H/?6��P7��C$����5�y�y�h[�BmPھ�����C�Dw�@��C�D2�Ik��d�2�s���d �ŹO{�"˨}?F,|S�� r�=���4j-�i��8{J ba?@����F[w(�k����%_�H�A�X5�1�e����A�5���D`� �I��oV�t��c\x�:|5��m�>�	�[5�q���Δ���J�)���URV4o���n��/�ޜ��u����|�=��A�(�'�xؽ�y�±��'m
��a��4�c��h�g�^v�����:똙�ʳ�at�C��M���������$��7@���HG	_�
v&���ׅ��i��+q�N�'zOs���?k���A��G��A9F<��` 3�'D���B݁�[�)Pߪ���a
е��z^]��|�7��됲cfb�B�u��(�&rkN�Ckg�P��H�?E.�=%V��e�Ǯ���C�l7��6`j�v�ĸUP�&V�Q���5�۷����Q��TJȭ�3��H�����GU��	Y7�qꯔQK�Y�����T:
M	�A����C����w�ߏ�ڪ�؞�&�92�f���8^{�}��[���L�3?��ۊr�IQmx'���"���W�<�Ή�{�!]P�t�a���.�%=J���)�PѴ���҃�!u8��y���-� "8KHi�H�c�!U-�5d,��Z��I��=<������Y]��i�R��۷a�b�nG̀���x�%���=�WO�~��7�tЦ.<��� 6��kg���.�U�(l��k�,Y�����Ƕ̅�A��R�_C�Y!`�N�e ^o����F����ל}Ъa`���nē)A
�X[R�B�R�/P	�bM��s@��[Lt�y���U���n���
���e{���6�7�Sޗ�Mt�ʟ��if��n�K�H��u��2�w�w��}�*�&�b?�p�F �y�p���)�,���Bz�e���&Xr+~4���e��o�?��nV���-LX��4�7Ӡ���h7漉���i�_�LR��b��г�dA�ߎ�q�W�_�`+�X-;�]��kf��4����;|�'�N^S��h���u�wn2�!1�v��G�+�q�}ˤ�E�� ��_l<�8m}n6�ں&�����������55�3�fORr���G�-��/�y������~5��z �w��yI޾A�������3��%��	�\R��\�ſ�j�4l��xCD$����r�z�ێrV�����QKx�S�O���2Ց���tys<��؏�H�T���R`��UV���nwv� �h�������GPؙ���M�O$h���������2vX�\BND47~��z#��ծ�f�5�x-�us����曤5�ǆ�7��|�E҅83�R��2��5x,	��0��kam�2PlMa�z-)����9�f��:qAόJ%-4���d��Fͪɲ�t����l�F�C~��=��E��&���5%����r�e��މ��u8>���g�ic��Ò8�Kp��Vpܶe�(n��ův��g��4n���uK;������o������ʵ�7�}��빈��'�O�J�ivT2��V�9د)��"]��pN�Jj3JI\�R�T����Faā�+���$C�U�X��L�K�yI�]�� �+�;m�d�G��+��q>�/z�7C���b��l*����0]�[^P��
�p��-�K�Z�q��j��b��덝�rdZ�޿�`&��{E�b� f���=2�<ZM�<�?�����~��s�z{�O0�R	�ma�v_Z_ma⾪��@��!X�1J�l,�n9�+�L�lb��q��>ʆ�|���x�y������z	g�yurK����rr�i�	�َ�����pm%�թ�������L�;���0�0>��,�1�F�zA2�=L�)Ku�����A1d����3���G�d�#������a���Z��o�̶��J	ԇ>��Wq�.�V�31�e^ �9��s��H�������,��> ᡌ??r�*���E��`���S�����-@�ƮD��vg��]�<~4�'�Q�v��e��?_"�^�@����
��3(!f���^���l�ܵa�m�ث����hJ`���G�H<k��X���?�TR�d�M���ݺ��ˏ+ع*D��,�,�7R�ELP L) =����	JU�-�|�(�;�)X&��=j�7[��ۑ�v]�N����V6�@��T��lA���E���nG���N��9ؓ����,��{Ѽ�$�#DY�SS��H���6���Nn ]��գ�>��a��o�e���g��)����o�LH[��T1�R�`˸(�Of,A��vG1k�7(��/nYKݹ�	�gJ:�i�����3������H��|���Lk�,RR��y�<��c�n�q�7)�3��	��w�q�~zz��D�o6M��:��Q�/�L|,��B�x'�w�RӋ��q��Hl��f�c�p}����1��0��r\{�Vw�&v �6��.�sA�v�9�jҵ᫜
UTX�b�7��̮1R���l���T�U7X�P�kOT
�mT_El�v[�̮}3�¤���)e����#�#l�2���b�bL�nH���V�����Ȳ�}2�1~~�Xcm#�kjC�������VeO�CrM׮����k���\��c���sKJA&o�M�.�Oc�ƪm�$u*惮�Qpb�՘\�3�].ѿ�~�葿l���-��9�x�"��+�Q3}\�~p{kG��ܱQ��oeS�|)�A$$�&�vp2�&')2��SX�B?��bؚ枎{ǎ����u�]A���jge���4
 9��]����y��7�ݷ�9\z60�;�~�Vk&V�E�&��Ec@O�u��zY��B�S�1���̱�QfD֜��m��PzI��2����C�w�M�N��BV��������,�A�pÒ�Z Er��)�G+{������e�(Q+T��u�1"��P���I
u�at$�SgY�kxu�-��,2* ����ҳ���tt�%��R��O��]�%X]��ٚ���)�5;�T���I�� P#y��Oa�By�	Zi���~�K��V-�t�VX��kxP�]�ܙB�����r���xo�qL<�{y]ZHǑ��SI��K24ji�"Ɍ�p���_76S@g���]� (�* l����#�5���+�����"�b
���!�� �WY�.�j����On� ��8ݡ��k����T��6˘�ĹN��>���]�9��b& �����HfWp�qMZ.�N`	���b2��P'�=iR���kH����,��'�#p刹�Ed�^7ۇ�5t���}xĉ�<X~���J�:�3�Ud�j�m�>�M����9=힁}C�9va��������X�)4��T���5A�!<��3ܦ @n{�\����l$@��f8��J�umiD���#�������)yK�t�܁ m~pQn�Qw��=tA��珜����pP�z�%�k�~#���d��"$!�� �yS�B���=��y6�t	�la�DDQ��ն��]�
t"��Ϛ֫7�M�2Q+�b�=^�Rw���R%bqk7J�ܞ�����>v"�y�#+w����a�H2Nn�,2�_+�����G�C�߂n�cd����O� �=W�1�b���PE��C���.�8���M�|�K��m����p�S�I@N�H�bC��i�]c�
t��lơ���p���!��)x���[b1�����>�j��nzB,�|DaE)�;(3ET�!��GS���+@Q,貮nF����q�6Y'*0�{� ���A+|Rw�z���l7$���eJI�ON��L�W��t�#��-e��Q��d�9��}�Q����C��&{w/tbU���Ǣ)c�ۗ�Tx��	����S�����iڈ��$�cdv���q/y�cx`K�u;���C�U�ś����H��=!?�%�+g��Z�����soʬ	���6hd�9�#8��C�Ǩ*�pX���(�M���\�w���+C����X<�X>J�g�L!����9@����$�E_��,.���7!~<�����]��;\�~�et[��ۻ�|�˿x��x��aPA�U�W3��C����'Io@g�WE�F��bf�f��}��_<��B��$� 6%C�fM�T[���<��xĔ��J�HB������qwA<�=��q5�|���J�
r�P�$Bk�����ؖ��{q࿵�V�*�в9t'��F5��� YX*+����żQ��9uݖW�RC4�ڈ$���R��gr�c�.+����}P@k��:���U�7�4��&��HE��w��̬�>�c;���aJ�+���u���4��QAbQ�on��*���X}�5�+gy�|BCr�6��J4�cS����j�)���iUhإ|\��idfY�����K%f����ǿ� Q�Q�jI�K����Pq�-/����PE�b�'D��qZ$hO�ʢ���#�ܔ��^]B-S�������O�Z��c2	kd�<��E��zނ(��x��������8d���,��	61��^
2�`nuf+-Z�/-����!���YYJ���E2՗�4�`�	Pd<����Z�p%��#��izG�����t};?0���Sw6���b8=���ԃ�lD���L�/�)�< ��@�Q�zA�@�ͺ[L����M���G�-1�Xj	�{q��"��0��= ���'j����R�KkS%*/30Ų���Fj���ai`�}����@��ơ'�3%�T� �$�js�ӳ�.r�w�����0b�5�:�O �LN��@�.�{�|^mr>�h6g|��T�,Qa�_��\<�,���X5�A��0�jM���-�����ǻ�A(��J�p�I�ڶS$��
~N���!L̿p�Ǟ.��Kf*��7��"��]��˰tC�!�ʯ�%��0�<���ә��2H��)�j�Ծ�L~��D<��V�C�&�z�|�3��~����l����3�g���8y�Nx���O<�C9{~�U�C(�=���S���x����Y�������X��6��,��>�`�m��'}���yd���G#(g�R��i�r��j�n��al��q������P��c+�#��(�P0��oh��pB(>p(Ց?��˯�Vj<���sCΉ^�!*[�&B���J��|3 �yj1�S�4��8ěݻם��DC��ae%B�A"�Lљ��0��Gl_�w7���B,�9�5�%�IoN3�$s�	5S�~r�+����ӟc�F�2@[5O��i���C`��y�=��_Zցxr>2s��Ys��fm/yP=ީPj���>� �D��	�������n���I�k}.�9x곺��8^R��D�?N{E�gw�Z{v�?��D����%��I����	�
��F�e&q�N֐?�>W����̗y����e��v4�t~̪��Zg�=���Bv���]$��6t�5qTک/�Wn�� �������q��|3U ��cS]V�����ՠj��!PY�Dq��°0z
���hN���F�`�'�\("~���V�4����w�$���ؘ�#+�����x����Z��q_^�h���F5F:$����ȸ}]!�����q�}w<�98�_�}������Ɣ%·'<���8Ys����FoК�\���a��M�7�%�e�b��Ae�{���E�X�C�,a���d�4�*W�͹-�jr�L*)y/& �c�� �t$�(t�4�Y��q\������g���S,I�H���s��්����ڳ<�����h��/��K��I0�M���ُ�	��,�ą�<TVE7B�u"�%�i��4���o<_�����>�l����M��ȴ�h�j��e(�;L�������eu��������	��J9���6h�%��=_Z@4B��L~��	���Ù�`M@��q�&w<��������M�	�&�-������ܩ8�� A["`�s����J����II�s�Rg�0S9����C�,I������L`s��S/� ,uE����Mku%��u��nfALy���cl��'5
�����	�u;�V9��@ΰjxY�d�H9m�"i_�Y+�HFяn~��T|K�Ca\��?�0v	+7`�ک�#S��KQfo)f}�5������	��@0(F���/<F�	U��`)Q�(�@N��Z(���ן�Pa���e	���V���ǡ��p܀�9��ف�)�4Z����3���68�sz�H���I�>�΀D�M�n�("�Xdo��Ԝ��}@߱����d�{���
��?���_d.�2�Zu7�8%�;���`7&������R*n��ܧ�҅�����G~�b�3���� vm�?�=���Y�Ǿ�{����\N������s+H�L����Q�|�0�O���M���Dn�i8Lɡ%+�[�1�a9/��Q�Cz娨<�5���ب��jhS��;���P�ic�C2�`���
����4&~��W;ᵀ����
��m��
��V�y��
ȂF��fѲS	3��)r|W���g���Jn޵�e7X��$W� &�����.�_`������'V��0��� �v˧�b��O(��+���"<U��I#'J�����͉���I��*���@Xe!����6m�J(W�����zڝ����&'��YJ�y$gB�T,�������VS'Ju���M��|war���O��.������/��\��>�U��ÿ��P�%���,b��uu�ו�C8��MֳS����a`��#nw�{/e���'h�%5�@�\aW1��/�+����L�=������ܧ�:���c���å�����.��p�/j
m��i�^q�������=��@QT� O��\ݩ����(��V��4�l�w�d���h���:��ɸ��{d�R֪^�R�3�̑��f؎	L�"C�iW"eG8�-��ڨ���ᢛPSE%dD����W�0�Wl�LWX�G-�L-�	����I,r
^K�秗�P�@*�$����m�,` �4Q冪Y�u�ea+�w/�'��#x��h�3��� ������6kg,!����>� Hkw�&޶�Q��X����~	=^kB��ܟYc@��� >l�����}��46?1�W+���T>�$���<��~H�����Q�L{_����q�8���6��>���m0�&Ա퓑8��,)ߒR�ė"�Ey�k]���K]���^L����r�+~E�ec�c�*＝��\��[)��u+���𮷡��̌�/�Gg�d<7�[��w=�J��e�(�tqK/9�SP1�v���uj/��H�=��O\p�:@���tI��s�o��$�`x9�|��z� ��.�-Y���bx���Ӷx�o7���OH�����D�W2�
H���9�66�>��./пiL���@���QL���ҠY��(��%�� R���÷2l�]1Rp�AѽΪ�����I��&B`�v�#j��|��u3��f���ɬ�c8�������m�o��;*�=� �& �>���l(��/)hJ���=J��J�v�y(�NZ嵭�~M��Vk��@�C��pu��#�Ь��c2��=��}��I'�!�-��uy�~���6���'!J����D���y�:�v����-^�% �q[��
n��O	QV&k�~��8�/�K��貭҂=N���ϔ��0 �#rh����dЕ(R\b �G���0�3�;�د��Sc��Ŷ�����f][X�7L�L,b�̥d���?ԏ��!�W�l�"�qf��|��\���Ύ2��y�}۞|�\�nn��Dh4���3F�]�֬@j��q����e�R.J�Y�@�h���Y���7w�.'�lɅ�s&l)I��bi	��Xg��3�"ʻT�e9]q*�ɪ
63��?8S�4n�}F�ܽ��@�����>
^e�i�<e����?���EwqDxI��߷	����I���n�j���C�3Xu�����:6��'�;��"sܷ;!�+!���Ɣ�C4F=lkJ��fD�go�������3�����\&�������7�4���Q�DD�ςՀ�D��?I�EgJzB.���.�㉎ۓ	k��v�f�h�h��a�P3��E�����@ߙɿ����/l�*�F�"�<~AP'�Q{�bI��h��S���t��'QY����3��G�aL�=L<��@(g���ŏ�FXfH���L��52O��w��E�0�y��07.����}�&� g#f���h�c��9�{�����Q]��̰E��!�h�����y��\�� mgOpo��Q]W�1�����J9;	�^آ?�nj���J�Z��c��Ne����������.�h���9����d�KԁSVh(��p�Pm]�-f�5��U�D�,�b��I
<eE"�;{��bL:QW�[�]�M%���˹����f5�
���n�o���'O�4�T��w(�ҫt��c�_Nu���<!���&�x#�w��pZ&nq�,���7��,XIcm��T��?G�eTl���O#�f�]��$�𒘠l���H
���b�+{4�/{?vf0h��5�����D.�a�� a��go�#'@��J0r.&[�o�����5p0X�#n�Z~E/vD-;bY^5�ݎ���;���M8��CB������xn���O~1[rk��=�I�s3���`1�zn�bh��1�S�ǡ�Mb�R!_c��~�����ϰ�CLx��hԩ�ϴc?�ވx�r��}��"x˧S��M��H}!u������=Bw��F����N��f1D�ْU�E���ly~�=0豌�5&W��)��$�H� ��\�_�v�jV���r�6�"�kv�����6b���()����z��������k}�H�&�`oI�wV
�鮨�<�����`�h ��s�͕�9�]��ۃ��U�:��a�?~�+�OI?�&���<$O��#/���Hv��]�S1���y�ś����޶�:��B�A��=�����^�*[Ȩ&݄���N6�$��(�:����o���e��{�C5=�j�~a��i鰲=�ah�c����_ɴ�V�M8��������r���~�,b���H��:���M�	�xޗU��	�Wr|U5
Wp�߼F�-ʃ?.o�1&�.�q�Un!de��w|�C(��Lx7VI�K� ��ص�O#Pᐫ�)��
�g �l?6�cY/���y��>J�Q�j��n7ڙk3����M%���;�	�[p�S���m��1uҶcg39�U=�$T8�����a����)k�gaHI��M����D��k"'�*8��_�ɘ�y��li���ɵ��1�����x���ơ ��(G�H�9G'{B�PoMc�S��2_����c��� "P�y��6�5�Y�S�&����V�`V3?,�����E�`A�q{t����B��o�S����d���],U�/��mS~�=zJD
�ũ�e�cxk-�^%��O�2�²=��%�gX:��/�̐#�H����#5���2�����A�hQn*�i�lge��̭Ҥx��R����(`?TI� `��W�:xf�h��O�)3�M���6���3U�8Z"�`��'�[���@/��ϋ%7��]�tՇ+?�O_~L��3�Ic:����~rr/@�N<"9_1�p�x�/�#��Q�.!7G��C|�?��H�!���G�Zv_+Ry�W��ի���/[M<���Z��Au@�f�> C� r0�'
�˟I�����}��>b��@	�Y�<T6��6���(�Ds���)im�n�V4' ;P��򣙆?�:f��D��M�8�5dĲ
\I	l��&����԰j���	M^�YχLV�9�^m�s�__Xجn(����S�� Ϯ���7=k�w��%`_h�"����=\DH��wrE0$��v_�bx��d0�zQ ,�^�����'|G�@�^�+����z���R
b����@+  q�!��.&�߼Y�FN
�5c:�f����Qn�����6}7���{�}=�j~���X�|L�֌��[|SP]�R
�UK��{�L?���-fW���#��:�}�ǜ��K�:�����������k4j��楟�u3ê���r��A+�*��b{Z&L_�����Wϛ���_�M'#����������[7�q��}���l�.����2=VE�E�~���];��=5}�ڒ�Z�F�S�Vx��1��Y�����W[�`y1'<�,) �b#;�Ql��2�_*�\����x�BﰥZ� g�qT������ݙe�ƹ�,�$���yVx�hم�ŭ�1k}}��,��@Ci���팰���Y�S�=Q2[%��o?�����N��W��iB;�X9 m�����$)�R$Ý �Vc��;v*��G�7���bhQ�ݷzc�W-S�4��P�����!�{ ]�i�r\)h��
��M_m�͌QgB9%�80��0h�$��Q��mUw���iY�d��tt����羲i��3��CC�����[���K�p�X#��I�w��C���f@�
�d��³^�&�������Z5&�a��g�nj�p3T�������~��d;}T�43����z�g
���}#� �8��9����D��(�����ǖxS��g�U��5du}x���q�>��}�k4z�[�P:�K���s��c��Ji(᷾njnV��swT��I���Aƕ��*�_���Q�Er8))��Qk:�~J�z�T0�4~���#�����ߞu���	;k�ϕ|�E�g���X����%C�*��^�zP�"�.N�!N��M��2�g��]�?�]z��p1Gf�.���{�,�J��˅�W�|^�`�ם]�8#�G>���'�����i�`�&��>D�^H�?#{��R�ąi@-ɹ� ���U`����D<�;�Hv����*��?��^��z�����?��-*"�7�eIՔmjES5w7X�c�]n�nV%^P�N����yc�S	/��ns��b�x{[���6�pYn��Q�������6})/�>�E��mM)eU����vM����������Ӌ_�`�'?�  "b�-J��`;�U�:T�C�4i|�I�G\�����O����6�%Ɗ������΂��IP��u�}��}�\C�S1��?O0e���}�����z��jm��(�P��[BR�-T�ze��~WP6�khr�&0�$�^r�Sj��|�ߡ}l��W�	In�+4��>�����˔��磲r��} l��Qe���ǫ%P�ڝG��?�J��[1�y#���u��>u���,GrX� �K���g4�Z��.�>�5f�dH�C��yo l�0�}��R��57�C�l�r�6?���b=�I04�r���bJ%~�[�"��Ç��E�w�\L�OIs���8�3���N�8�s~g��-�����,�0\dI\+ȉ0��B�&��4DAᓳz��&�Bt�FB���3�Ǔ�{Z�e�q�u?� L$�ya�;+��X�=
��Q	ĳ���L	���Qo����f��+�T�A��G���\�ڑ����e+��$�L��6BҲea}�r�����`�{gxq�6j�?H�C-��1�2�L[G�Щ)kHM��N�R���l��_ɼ�(�Y&Z�q��{��*I,iX�Ă�J��j���M����.�?N�[@x±�|��]�>����:�+�j|���&�_�K�21u�Ws[L��7U������N��xISfCWĢ��{k��~@�vm���6�Psg����ޖL`V�WM/.% ��縟��VK	���N��G�Pk'o��,��=0���J�f�0���F�T��%,^q�����Ze.k)؟5)���8�{���s=KJ>Nӆ��b�U�����sݱS;~`��º���>��@�e͕<W�C��aΉ�g�&�*�����g)�t�i?&��z	ğ�k��@(g�SdP9��AJ�#r�7��5|.Ih2�F�!2�m\|��a�c�-4o��zSY����(��{{W��]�b]��x-�w��h��rn�C��$K_���k��������$է�3��4�ȾAH��l��T)՝��Yխ7A�8c�U?{����ʰC4���mj8lˠ+z�-�����>�2����1=pӯ5�|l�p�asb�|��D(L�����"��(y�u%���۝=��OG�8�C����䔆����$60�+a�S��
�)S�_�u�[K�g��,?xv8��G4�7����D�sԸl��`-�=���c1J]	���j�<`;���a���gC#�`6�g(�,�����KG��fL���Y܁�40+��DW�w?e��P��B!������'��D��@�����pxp�i��*s���/(���f7/��*�͒�����9W�rֽ��:,����e�=�c'��B�B�]�R�o�21՝�1QN���k-Z�AaDw7)V�O�X�l6��t�m �������J�{������X^Q��L!�_+8`刡�>Sr�\�a�$ ��cZ�U��b��|K�ס�XCω<���VQ:�_9ig��@bC���Q I�*���GNq�0O�0dD9��>ƞ���H�	ynTR���a�2���@ꊩl(��"Jn�&�#Fb��S>�u�WcOqV�D`s��Ԏ�E|�"0Ұ'�u2�f7Ң�,�*7�+/�����)�L-�)��H���E����ҫ{PK����F��%�rP:�5TZ��b ���y���v��)��=M���[~���vCAx��*[�x*/�a�DWQ��w���8Ӻr�s�m.��^�0X&�;�+{6�27��1f��d�/�c��7��
%� �U�B��|���j�����_eL�cw4-���:+$c����L�1��dpZg4ե'Xv��'���PP���`�J[>�>�3'I�%�Ѭ�v<�� +�+آ���~�gm�*7���D݃��r��ꭁ�
�h��ᦦF#�n+8����*K����� �Zk���
6`��b�'ӈ�ܓWs���A��ZNݯ�N����gW��[̋�ğ��d���u	���cc��/���n�����}^��ܥ5�.X�f�ȶw'�5&�!7߆��a���*}5s�B�7�;��hc��y՝_�M*R����&Y���˫/ߚ�iw�z+�^��H*����V1`����y䫠�(���d���آ�� ������ia�tPL�/��|lL���᪁U(��g	�I4SDh{������(�\I��B��B(U���3�f`�V��!�A>-��#�����Q`��R���YA��d+2���D�<���/0�7�+zn��5PO!�vnm_�o@��g:�דG�B���L��B�Cy��X��ؽ�~m�)���;��&�
��
`�b[���^Yi�� �X��Xb`�m����W�w_��!�Q@���g+s �B������?1˃EŐ����Mc9��U*�>��A�t����LP�a!���f�$ ��_F���\�X���n��.�J��9Tu椬�9`ˋ�w�O#��$8X��������I�*�m�h$�*���Q?����{�Q��#8EX{������ٶr�l:��1RV�?��K�w�X��T�\.*FX�s<nX�164s:/ w��D�l~��b>�+Q��h\7���Pv�')��_�.-|Z��#�������/�,��+����k�0{�I|%ڄ��x��oc6�@��)4+� �&�����c�D^�p�u�h8d{���
387�|��c3��(�����Dg�Fů�O��Q�
�֥jv����;�L���)D*�J��|<�*�;�r���b�ֈ�	#^΁O��L0m?���$�GMJ��4�WN�<g{mځ��0d�5L�P��6`�SG_1A�Ѳ���N}�lMY�X�LJ`o�%`���� tiV,x�	]��uǱ>�FC�(���L/�U�m_<�7��T�u�4�7�c7����5�>F�o(���X*_�~���`u�V�w����V~�9��W;�2��~V��8�\���$��n^���|�vbC#s�&���5Ұ� ���~4H)��F��GO�aI���IZ�vsv�oL�agM�S��◝�<�v����n~�Qr�6O��qm���W��%
y��q��bfW��"VH��'�\���LN��>�8����z���i�Jh>��Ӊ��~����l�x�<Yś'PU�ִ�5�d��ipHQ�ӱ����R�4�F�\;4G��/E
7}�P/֯������GRT�O�Hѧ�c���$��!����y4Y
/H�<ޭ��9�f���l��Ŕ0�?��i�l��U��BJ�IuKRx��.��	![��8&��>{�@��ZH���9\�0�|��Z�����c|6�ys=F�M��8��e��K<d#�{�����ڪ��1�J�@��`�3샭���9��7�a�R��1�V��wс'��ɹ!�k����!�y�n5�>�z&��Ģ�Y@צY�w���_�"8]���o�����E�:�޼��b�S Rzz�h����2� �����h��}�z���tD���J���[��#O!���XN���5���T"��'9<|[�H�&F��'�����(K=�^kƁ-���6�|H4<�Y��~ֽu�6 �D�K	O�(�D}f�'��>�J�o��W�e��H�������5@����y�RY�s�9Ksh�����r��F��K��XՐ=�=+#�+�4k��8jRc�[֨�6����
⤜hE1j��k����=��L�sw�݇V�j p՘�Z 2�,ql�V�u2@v .��q�S'����R�b����;������2Q}�n���0��%�6W��b�ї@�rD���l���pC���I8;���̠�S`�f��n��!0�]QH�+o[Y'�)��dl��_�?ɗ4��`Nu���n#ԅ�K�	%����7<}=�]`�z�����.	�Ib�f���M�=E���SE���w��q!�C���6�[8�]�M8ڦ�I��͍�Q�(	�Awe�s%V�0\�cy�)���$ 3`F���Iҝz"D&��L�fZf���nlz��+̑g�&�,iw���GO��,P���A+��0���T��ۻ�P��@��PP-����bס��hJ����w���x���sZ6���0����R��@!2@�rdU O����)�N�|�~�֘�W�:�?�1�*�Pߧ��@~ʳ)��DL����Æ�tݖN�tʿ,��c߸�S�=t3����YY�$�~���x�_Ru�,9di�5�Vu0d�e�x	����d�,�x�0�ч�U�4P���a}��)D��ǰj�8��)y�EU@��_N2%Q�6������Z������R�=��Ցڜ� �I���M�@�J�?�h��0��7�)�\~�$��G]����V�:^���ɤĈ�Ot�¥���J����L��������׻�JO�F��}m�K�p�ƹ?L��zʚ�N}Ӵ{��K����ڑ��҉'��v���@�_X�ʹ�{vϭ���c�1u���O�^�~>�Ӫa�J\�U��}����8<��`B'_P�����n���xW�!�Y9V@,�2K�h�5��	(O~�Y�?��v'[N�"cf%|��sl`E�->|��q����;Xz٤��ܼ�����f|j?���?��&��+ �wȫ�.(N���8:�0(v�B�۪d�$���0��������+��S��Q�t��~�>���hV�-���;`W�b��fcD!�����2�k�\qw�@�R)�l�Z�*�����ַi=J��,����ױ��9h1*�iªC#�φ�ޠ5��^��Y��5]_�o�I�-�����c<DP�ȭF(!k�ET۠OQ�v�Ifȸ슰AK�%�I|*��e���M6h<��o��"�	��:��CO!�L%EKHШ͚��rg����xj���n.q}�]fj��L�2߆>��=ʘ1��ǰ@�v-s5��g��%�����>	
?�Qٲi�9���G���1!�5�J���L;�(��¤k��q�-��,��cY�H�4��J��UT��{F҉~t����Kp�E�*��kN���k��#���vj�i��(jV�'���lc�^�o��59f�3�վ�.s@�y�����P0�\��-mu����ҘB��=s����p�U;e�f>B���)5�R�-����d4̭�Ex'5�~��?���:P����u�Sb�CG�K�&0���a�7��/]�g��7W���<4םq��Ȗ���YS#,{*���,FH*�mѼ�a��O�t�=]G��+s�j_����ww��z����1�Yj�fNJ+e�1����(�]�I�P���'��=~�WG� /A�����~�/�&c�߷^#o�DԆ�����X�e�v�&��}u�`�|�s� �O�@��-dt�3�bXʈ��^gD���-l5�tZ��Ҥ�ͱ���4Z��UF��w����$����$$�x��:�d��a�9��|`�AT��Ig�x��"Ak^ȡS���[��j	N�D��c�A	hʋ٦?�V��1��I���ϊ��ۄ�N3fYL	���}��
�af��hY=��I�}+[���tU��|��3�f�M��zcLA_�֛I"�TX8�>����h�9D���n@[���(����\\�d�����@��� ��ԭF�����P�����~�hP�Dt�'SAA_c�趰���2�&ͷ�c?���g
��w�6c�%����\k��!@1d������G���_�g�sb��	ȸ4�L�^ZTV��#�=�����z�N� .��_҉Z�'�!�
Cl���1:�1ʉ��z�I��� �4��ʘ�/���*j��+�3P�M�*
e QT��Kż�"�0��JR0;��?ڻ�7�
��S#Q"�73@%�&`�~c�91�.e,r��X�x�B�	��V�Z����F���ﮐp!-.�HS��B�(h��{q$������8+&1s',�5$a|C=��Z�q5�fގ*��{�vz��:�I#��۳D�R�J=�MFCN��s ޅ�fA[:D`�����z?�<�^�o?P��fkm�G4.������>N>���=$P9$J �?�X:Qa,��;*S��Ӌ�,��}Ci3�1D�3�2^���)�qݰ�����J�M7J�RZ����
���`�Q f���{[���0�3>�b�>�҈��Z a�u��>�1��+sK���O�i&�j�v'��?��DxC�$�R9�G�c������)��Sܸ�A�s�3�f��x�]b #g�׫3!�tob��fw?$�w�*�
���|l�8Jr�f��^�j��6����\J<0.`?{r� ��tK#+�g �n��̵d�*8����Q<�<<��WnFS~��*�,�j��ߵ�`NU��?P1�ҹ���D{�7w��Ik�m�����y����?"�s�j�x_S������X����#���ݡ^���۸���1��3��DD݊|3�[���iHۨ���T�,W�Ұ ��nۿD�Gv+�R.�]D�M/�g7D��F)�?�BZ�m���	����|��/���H����&�t�Q�� %��ȯ� �(�Ix�Yzm�0�@T8���	eM�p�mV�eNG׋i̿��r6" /]�T�k��Şy�P�?e���2�k�sr���7t�:����y*������5����y����>ե�M���`�I�s�	����8�{ 5�!��2p����e����)7��c�/Zlg9h�^,^��`��n�8����L�o���z����h𝘮����lwy��l���|s��T�r�zݛ���?��3l�o���m9�����XG�o���*"�]��-٥��, �+�a��g�)~Ԣp?,�,��9Xj#w��6!%^��+�+�i��N�U��>s�nV����dL&P���Ե#��D����� ���g�hpe�eg�w�^�;��;V��`�ȓ=�N�����.?7��$�7�x��"-d�(.�&�O����v�NX|)]�����A�W\=���S�F%�WPf;g}Č��QS�u&!1Fdt_bs��RH_��#k��kg�m¿
�X"�ԘI^0i,�ً��{6ݎ���R��,>�~�+�o��cr��O��rC`��6�/�jְp���U�,�%�ij/��N7������ۨ�t�,`?B�#�Wqp:��]pR�y�
�ȶ� -R� ���?RT̂3��Z�L��-'�[����}��	�^��\��.?.`0 5]/�?�����byΘ�0�G�v�`�O�Q$�G:�8D:�t�Z��}&�6��0��w}!᯸c������>I�֪��uW��hZ |^�l��6E<ˉeF?�	�V.z���v S����H�L�|Ҋ}Z�p\��E��9�؀�j��L"���ֲ�7�Es]�k$_���CT3.��.Q��l��a����$�f1K�G�����c�6��ΰ�@���A�=]c��ku�ҕc���W�E���k�'��������A-��{-{�^�U}��������cg,>�N��]�'h1#X9�/V��;�3wv���t얻g���J��Vk|��Q&�M�¶{�0R���`e}"Z�y��E4[;���k�q����ا�IH�PC�LW�Ԇ�0X��-q�JT��!�n�ƭ+��P⼽(�QO�ٝƅ�J!C�~71�0�$FvC싰_IO�,�ny(�j�dX��}�'�^q�K7�.V�} �[9��b�}U��X��H�z��R��,W��_������:@?#B���:D~��-�>v�>MGV�|��#/7f%n�}<�����DFBs��q�5��8��7=\[ƍ�&���L���ދ��h�t|&�Z�y��h�6�&�WM���X�� .��Q���^3αI���i�&�;@ye-u�R1�h�B�����@K)2Eڶ�Ve����kr�4H��96̷A�3oI��
�7Y�� 9�l�$�v��(G��1���G�飴�T~T	�󋭂vJ�Z�=5$Ҕn�#HZ�mq�8�������gڴh�Edi��R�?&QսA*�绽���Y&d}��<�F�^�_�T,��*8;�
}�H�k ����,Q�&׻�cAD>Le�Oٱ�,i�M��z�?9T3�Q�zeN	xpR���n���x?v�v-'U�&^ӑ1���sO:U=Yo�7���Tc�CcE�F{dLI)4�(~;��`K&�y���/�=.�C ��������p. յP4L^ρ�u�{n;�r�Q_���2�9���Z
�?5o�O���f/�7$WQ�`�{�d�~2-z���+��K�S��h"m�P���}�;��-��/
ט�Xs�m㖸�$nvc=����k�K�#���l��>�?K�4fO���x�|m��[z�V8Z,6�U�e�2��C�xJ��N���爐�q��%�����DL�ǧ�u�<vd��dG4�m>��+;�<�H�8��Y'���,�B�S:��y��n?O�'"���s��PPW�ʃ����U_�_د+p%A���e f����΋������h��~��������j[5�莗���2��4��~�w5�x>�����OŅ�h�[kQ��F
��u���5���7�{�����L���n�8������.�9�KM�����C]���kY�Z������>��㉅��[0"��C�v	_����5�=�H���i��u����q^��1��O�;��%
9\����i{šzȄ��%Q]�B��Qp|,_� z�R@�3;�+�����Rڧ��(=�<���k��FY^I�T��t�4Z "4�r.�(�Vi a��W��4����ڃ���B�����@���!���E
4����]�h��*�p�����g(�݇A6�͔��lђD��wz8�7�q��
J�k|w�2��`A����2�"��N��-_�Ma���Õ���ET�� ����̙���)���B�������jQ鹃d$<�,�eB�8W��@�%����H�P��~�@+Q�V�Woaӫj�?���Y̡j�z��Z7�R@�����ҕp�Op`�#�G;6�D@Ym����Ȭ�,�Yu�*n�N�(*���O�����u[�Yc�U����b��HW!��M���x�������'�}~H�AI(	X�;eXEF��jv�s:Uen�-���M�Z�U���˹�סsU���l�´1xŚz[��j[�6�i�זN�,����U>,�;�'�{>s&3y"+�&~�,'ͲMU�b�E�SVy�ᱼ�s��Z���4b񖿴�1��S�D�!�	`�`
N�E��F���ȅ����i������ޟa�~��v8��*2� ��_�."� �����~iw����g�tu6k8Ųv����o3Ig�$��grn���y���.MNl�J�m��[�Y����ؕ�uպ���U�;��P{Pgtn�+�m�kܭr�,�D�t
����~�/�����Zi�/�l3����m�2��]�q=`��M��cl�y��*�|e5*�v��CU�"� j>�LF,�k� 3�){��J�I$#������_����>I��3�Ԓ��id���E����,,�g��e�ֻ&���)&t=�w����6f<��ϙ�&F����O,�&QL	&�V�a_���Ȫ�_]�m�mG�ﯦ��?��2������)����^<z����mKo� �z���<^|�r�;^�2|���Cf��հ��'�I��D��i	��M�G*�H���zu���[��e�4�t��,��(�1�Â�e�я0-9�2]��F���,���K�p�PyI���,�n��y�8b҉ͭ���'p�c�z0���{�Ŝ�|�RK�4�,FhQ�Mj�U]B!���A�a�Ҫ�IY̅���{����J/��a3�C�v�������@�S6*ھ��ѩ����+�I�^9���w�O�ۛ5HG=;ʽK���[׽�rz2>e�BԔ]Q�C	_��r�a�]��7B���=��d��#�~x�^q{�b�6r�[�9ɺ��W�ȁ�k��M�s�|��e��[1��a���=���r�u6��W���-<^G��"_�ёt��ŀ�q	�䉆���/t���<�A��j��29ذ�s��j�e�V�6)�6��
�fBy���w��+#��ة`R� ��P��=���J*��{*�J���}0&�����rY�ax	/���
%�PN��oL��_�)]C�`$����֠��
��n�c��Y����6|dk���zFW\Pt���}	�׍<�C �)�֒Y�FfrAG�A��ޖ���ȱ_o�eI;� d:��)��36]��%�h���P�҂q����{���l#'�\%a2�w��&H�� ���t�p><{�V��I�,	�\�CJ\1#��*>:�̊������j�%5��u�B�t�+�D�����;�k����.��23z!����|66)R�Fb�7w?���W~L��������Mj�ܬk{���L�5e���ZS�9*�.����5�ʢJb'+�zI] �kL�b����H�؏;�CCI6F��/��R��	���K��Kĳ`�VPIċͰ$D��]+1%3�g�l�n�y�O��֬O��5�Q�&��#���[_Ɨ+QB��qG�~��@���7*�Vt@�T1�簈	ݥx�?����%v�nR_[��4���IV�1Da�/���p�}2Lgn,���0�,���52�y�Yp @�2�G�C�	�C����`��˚��ƸC��	t�>m+��]B�a�X*G�w����t\$k�*�Cx��V���M�y	>�vsU��+���%����}⑤� {�U�s앇|!#,�	�0Y�-����O�;��6�;5�g�TX�`9h�A%l����ࠊ"fո���غ�^ew���P��źD{Hv�=�#2�p�C��l�Ii�BC���p��7�k�N�^X�V�Z�5qU���)�]���:w��6���p\)�q���:W�-��"�9e�k��-w���_,2�&�d�8~��j�2��8
�|�X2�Lm�W��ٺ�湹�'�?��V�[��Z8��'�2�Y7�ҳ���0�p=B�����/��U+��Q(?M���/b#��8�ܞiX�*��B^�Ҿ�ے70P��i|�@�Z8�m|lR>kZ�E��w�zԶp9��X?���s�S^�$���eb҂Q�,�١��H����F����yV�@�����L*f��BG5��s�N4t5��:ѹ|f��&��E{����fk����L�����ڠ4u����w�>Z��&Hk�j��3�XN�$�~�d�yZ�<Y�؏H� �g^F��Fso�h����i�A�U@�.�=��� Fh���öq�߽ٛ�R����;z��%����~њ�����|c�~:C����L�ȸ�6��rlV��h��=���?��A�"P����=�ao'�U(�/�m��=4��O`Z���o���_}��?�� �t'�CJ�z����>h�|<�yF�K8�ez(l�m�d��Q9�9E,eH��tK�Qk�y<�Ox2B�T��D��բ<LJ�T���n�Vc�h��q	��_�
��J�w?ǭ�҂h���gQ���PCC��5'�}��&�;GiP|�pΊr�����0q(O��_����>�_��i���/�
8u���g��N}��2�q���V�iF k�GS�	_*PBM@�_0�c����>�!���4c��+�c%��	$��l���;+��D�VJ�58��GD��̶�GA۳Ď�А�PLk|��l6�ƿ�X݈��`����U�%ʟ�?�q\���5�,����:�]h�.�D]��`fn�o�R��( �R1�O�����[pZT�BZX�"Sؿ�Ci�[��N�_p�7�i(փ���ܮݺ �UH�pe�B��wT���H?1�&\�/|�p�'lp /�X�lky0�m�<��3:#8�/\�&�h�V��ɠr�W(��X�~�|��y�_�B5(e��E'�IPӅ�<�.�1X��͉-0�S`����M���˯����0��h�(wSI��H�БZ�����Pf��)��Q��\�иԸ��k���F�(ߵ ��vRx�k�7;�p: w�Eՠ��@�k��B�����[ɐ�]�7�р��tk���}��HɎt�s)���\�ڕ��N�9G�� ��y:���d�tE;ü��\�7�,s7����m�w,vϡ⡭֪C�9�]���f|;�lr�+��-�|"h�\B���N�	��>�n��kp �Y��4���_�r���F�$�o\Ăt����i�]�$�?�\���L�j�	G^��v: 	���(S�}�h3�>����
 E&��j�2u<��'8��Hb�Yڜg��bU@!=�d�!��D�)�[6:a((��R�~��=�M.��{��cT�'��ʣ��n �OH|��'�Ǜy�Qr�L"�Gu��Z#�:��Ш�����!���H&kԈT"g�ay-�fc`�]
��[�.L����z�;�U��(��E�F�Ws�+�������I[�Ȝ�q�����1�v@�0F��l�FL)���<����0�ydqР%�Ex�Y�,�5���|�N�~�:�[f�-�#*����, G�0�m��R����j��+p�h�rTt�cZ�7v�
�ǈ�땫
M��),��!���M$��-e�z*m��s��|�H���� ���TU�T~��f�G	��|��#4X+GzT��n�P>�	?����	��e����J�)̬��~��D�����T¡tNͨX��RX��3����oAZMh��#h�Z��\,}�UG$Jv�9���cIj�a*����ա�� "^���+��a��9���� �:��·O�8I2^MF�P��Ҍ�f�g6���z[I ����*k�W$�X�5����B,�Ep�o7����B�^����2��,���`zU�Q(��B�Y��PI��4������
̸��>�'�ipZ�nC+�T��7,���rM�����[��?�������91:]�b#Xso��ֺ�^�yrR���F��O�36�F��H����W��G�Ύ�`-��S�x��nx�������AF������|�Fw���n]�٬��w������(�	|Ya��M�����s"ar����p_ڮz}��%0Cq���T~	|��d�"�~��J�q�(�zn��'sPӝG������Z�	'N�35�!�b4n���h�j�Oۃ�قN��D�M��bp�D��:~����u���'�v�2(��X�ߠ�4�-Ʌ�B9�r�F����	#�J~��x;���_gƯ��
�ӳS��@^�NF�q�l����~�����Bu�#4a��*�
�l[��npͲ �H��Ř�	��f�mˏb��KFc�xL����D��+-i'�@}����A�_���<���h��q�3���J�;+��y3b�U�ޤ�n#�I�uv�<J��3�*"l�v�p�h�V�0	srE��\XeI�(>?D���_�OV�ߪ^��d�4���gr�V㯲� ���ah��.�˟��T��L���C�W$��VC��iA~2^�� ����ǻr�d�д:'�x�M��C��q+�lo���ŕ�R0�"��|�$! ܒ�YQ�	8��U廾7����~ �{�YK��{��`��woN�q�|V���Ɣ8g	r T�)�C�(�*�pȮoc^�%�_W����*��C	���O^l�ƅ�u0���^�����|���R�+���G	�O@��1n�Б��Y��ՙ�	��!��X�2���̷�
]F,���}����^�kŒ��`���i����V���Y��6��KasG%'Q�ǐ���h�Z�F��[�t8����V8���W��_q�)Xz��ԑ�܉�]��y~�����'"�S��r�����A����O�X��g,��]��5�����W�k�D5I���,>2R]������=�P��a�1�XU�*̈��{�`���=�������x�G'����.ڻ)7@7 R��յ�C�y���Mi�&|6G��8x1� �/�]��e���k�>��o)��hϔzٽO��V�!V����T���kp
\��WH��'јhJ��ܢа.q��F.�	#�<f.TʫDt�t5�.׆�n����v2�����Ξ��}Iu
~$�>�R�T���m?T=O2��T�L���		V�!ޠ:?�Ǌa��5�91Po�P�0R'b�(<��t�=��,��_���P����fn��V���k�s��#ݢC;�YqTPǵ޷�������) ��ԧ�,��W����[�;��T�%i�)�BS�&_������3��|�&\hV(���z���au=��ʑ����^���N\Cp���D����O[h-l�bJ�׌�n�ْV�~s�B�̿��Qc��[R�^���+ھ2��V����C`a��,���bP���B:����(>�����I8.�A�2�9���҅/��Xw`��H�M������n� �'��=fJcC�I�r((�x�j�X����h��è�,Z�T��dc�W���7/b�����s�O�I���c@j*1������ޡ�J��g$� �䏾�=��w�H��~y���t��)x�Ә�v�`�79�.�P�6���w�����f����9I��b�⦅�84�w�]ݍni��ʛ;*��Q�������f����P[��o�^�m;u�w��Оz�eˠ!�� �&�o�xh��)�п|!bY�0B��1�IV�j��Yl`FO�@�Ti�Gͥ�Y�맀_��#a�&A �?|p�\Q��Q�Rc8Rހ���(R�|cm0�i8>c�����][��7���C����e�Gk�'s���	��Ǩ��`)k�+lrRieJ-���>�WN�#��9'�6`�JE �F�{���S�gX���H�Mf���]�d|�-�y��iB4+�`�X�Q���(���Z��z̈́Ro�����U��&��V��I�daF0f��~�hW�iȳTjℓ%(I*�7̟c��Z����f���y�Q�[G����F��JӾ���W+��g&P�G�Uޒy����S��8�xv�TN��#^�}�d�ucg�Ӝ��<ME���M
<Y$�^j��E�j'���wN4�F�us��>�xI2\��5��{Ho�o�\���d�z1(���\6=�!�C`N7�I� ���юlĂ�2�͕�'���6�����A� �}fA��2����s���B�33�c���A�������`�6����@\#�kd��o�L�s���/��}�B��F����6or�HK�{�Ƶ+��*����\="���l�D>�!GH��$4	� ����2\�x��3�'�z����\g0w�T��ȭc{�8roΙwOt�>��|cH#΢��I��-ݦh��k�B�,�4p'�3�A��f��lZ�����l�����l�8��zs��g�fǕ%����c*v%��M������������K�����RѰ\�C��l��@�sT� 9]���ۓ�K�)gPNd���G�.zs1��4`5ٱb��/�ԟ%�X1"�v�dHB�1��(e'��X�I|�O��ہ��3��H<�Ȕ�����\"0�y!�>��;|~�ZP�f�\�7[�Ë�x�O?p�PUJ�i�`[�ܦkc2��G�ƌ�~���~ӋA�ap=1fs��e�$���:�Z��"�<��Q93��ryF?g������o��W�ˠe�0(�����G�U����r+J׷)A]Ʃ�k?V.A���pG�-º�*0}�2W;I��K�Jk!Ӄ����g�y�2��da<Ē�Q�.;BtVamٸ@6�^Qm-Q�#@±��H�:E���G��ݝ���^��:��+(`�Jy?%�;J���`9��9��8)f$۸j���B�(�d@�>���,_'u�!\�H�:���`=�b�5*j�o�#	Ǡ�#v#Cb��9��ߑӾ�^��{\F�}��V��S�BZD�'���p%7'/��i9�0J߉�(-w�� ������*����+�q3�`��W��Ю������oɟ@�؋�\kN�A1רc�-����겗�?|��O����/g��
��LU`��Ʒz_L {+<���U��g=��̸�Ʋxl�l%�\�����)7KIv
l��!i���V��c�]�%�!G�����`��5��^�J�	�g
o���=!�K����3��),����1p���؎#+,sFz8L�!�3H��@.վ~�c��
�*fFsLW�jp<�z����5� �1Z��r�aa)�!2nT �ȯ$�l
z�o�,c�2i8���KU��*����;���+�z"J�����+��nC�#URq,\�#tn��!��h���|l�:��_���h�_.� 0f���#��p	c<��k۸�hx�Ia7Q�s�rO�FZ�3��%�Ab���rC�ez��ꑵ.ʗ���var�|��G�T����p��~"�L�f�~����Ue�B��iK�-�R�8& 2:��T�g�L���A� Y���u��B��/���[�����p�l�z�_sLܡ֣�,Mǋ�@ʺ6+�A��i�8��Ⱥ�둬Mp�.�4[��V7۞$���Po��S��9G-oy�%��Q��G��[�L*t ���C¼�P�W��� F&l�"N*=V��,��"ִ҄C�R�A����?��O�}�E��W.��V��GaX����O�Ϻβ��a�&�oUEx���K�M����N���O�΅�֥5����V�
\���������I1�@s;jk=�;��U���r*xA\sRdW�;s݀	_�r�<l���.*+糐�&z�_�ۂ��"0xgkm���G	�'��bW�P��'�Һy�"͟Q�c��6����j�j��D=��3o�]���D�������ܶz�� KF�@��$��WI���
v��>æ<~������Y>�H���>����j�;d*�R����~��m�T�x�(O�Y��W-�0�������,h|055���<�e��S:B1L�rbH����}�ʤ8���W ���S�%�ݐ�ʃH�t�ظ��
�>��Ҋ�ǡ7���(�mڑ%t2�(�[�4��������V��O�f�]���Eo�6��$����*SΌ���v�~�ff��G�����{.�T�����W��'�6b{��I�lE��uz~2�B1�����s(Q�#�I�G�I�� ��s'�� 
�u*(����D���ο~�ed��AD~�(b����8�
qCiC��u)��������� ��kݳ|a����=r}:�
��e�
(r0��2�#��C/�[/�t��]��k�"Bf�ƽ���b��o<�`Ͼ��A�3Ū�P��@���$�7���*�v�%�><k���R�&�^��9��g�5}*�f����C��H��᤻`C�����Y�����b����Q����:�%q̓�щI��_���oU�c�.e��eɧ&�P�(���X�@�g͈��CVW�"�#��$�C�2�B�׹З��YD�r��C��[�@j'���J��T��Z��W�S�`�S4��Ň[�mʛ?�B� �/��d�lr\���Q=|��#�Tx\��j��En�YVp�E��$��нD���2�gb^芎Ԛ��=g�� ��W�\?��q#y� o��Nx�,�1�؛�H��u'��!\k��nvxu$j?��w~���������3��F��N%N����%n�����Bێ��C�u��DF�NyCU,��#Y�,�rw�ő�*1E�M-qM໤4E;�	H	fu���6������$se��
WBkH~��9t>�b�����e�a�}&_�N�Nd�.���n:�_kSB���N��`+=H���E�V���F�H9&&��ό����[_��i�/"���&|L���!�!��0�<��"&jbu��ĢH(���^�p�a�w�nr�܂�g]����>������;��[y��~��at���AG�L;�=1��tڊب�wFj=���XŨ�b,x������.��b�G�(��F����yA�ׄZnȷ�ʞj^H�#� �n�EpXzi���u�3�s�o|���"�O�� �����?��!8vS��?�	�+���5	?f�7��_��J1J�+ʻߝ����V ���&*��$����f�#|y5[$������R�~��Q�-
� �[�|�V�3�)h�����S�S��Z <
�¿���[CV)���r��%m7��rY�[#U-y+�Kmj�Iü�A�Qe�� �l��x����������!�y� �p�(�2(O�F�0����.F��pt۠����tv�>�� ��C��H+NO�n[�4�HfT60�^�`5§o�*+6<����)$�1�\m�2�.iij���/�-i	��H�"Y�+e1;���Ӝ�4�<����4�x�s����u`�}F=�j���I�J�7�2��i0K��yg፿H�C'��*���rmXV�f���l�dT�lT���~\ӛ�!	�*�+�}GO�_��T"ޭ��8�̐#.�
�捭	y
 ��h��[�R�j!�--W��Au@D�3��<<��b�ƈ�V��ҦhnYT���x�����nV��u|�
,�`te-5�ι�O��ed_>+W�ë/��b��a���{�O �Mҥm�/ӫ�;�q��e�I�.�\�f=kΫ�����^�~~p�Vʘ��"��O��>�<e�Y���3��,Z�L�Q�0V��t�	����L�9��Ġ��.8%
;��0E���|�f�Ϡ���́�=n<t<(���.�
���'�?<����cHK��Q#;k]�ݸ���\X�>)�3�b�����KI�/����tlﳅh��o�O���L��Z	U��ؓK:�Ì�X����i>
��N��>q��J~�)��Zr���Ε����8$]ԕ���в�I�L���H���Q����E�3�"p�b)ӇZ�:
�n���R�ŹL��`@z�"M7��x#�?�h�r���a/�G) #��� K�5�zSmUp?�R��o�O�)��Z=hX�t���i<7�9�Z��D����f\��I�3��+M�����w	�f�O��'D~�o��#��\pr�$��2���Fʡ��e|X�gyt�e���+�l['�оt�'ɧ��?�"v��j���BQЛ:���sE;1�Z���{=�T�4v��OCK)v*�$�����uDۆj�J�՞v�+�u9k�xj>�oe3�>^��Ghj��.��LRQmdѕ8���K=R,.@�H��7�w�	�QNW ��J�(��z�v �7�Ḵ�fK�j���<Ԁ�*D�7��9�wmi����$��}~��H 
"$+'�@��)A{]��8��8d<V���M�1Eo� �����B�_��VE�c�Q�5�SY�o�Q((�j'�o'�#���P�ے���kPDV�R3[�h��+���,R-�b�0߇�7�F|r�n�}��;0$Ѝ�=g�:��j9�d&�2>}�/�\��F_Z������Qi6K�%��y^yn�gO�²��r��1Ĵ:�6I��U���ya��ҝ��:? ��2_�t��&KE�w�~;t'�N�c��$'��'	�h�u�p�����n�\k.����@��3lYr�~R�������e��{�t[cF��5���m:F�� `>!��c�
D��9�b�������~��.G���Y?�-0�*9�xB<��(ap������Kt��ņ�/�Ʊ�Pn��Āq�1cJ`�P�0ˣ���䁇^H󀨇NԊ�J����g�{܄{C���Y-��X�7��*6A}+N �s.4[��Φ����.%$ٱƷ��L/Z
�C>ѝ���ա/�u�qS��Y�j�v����@}�rb7�ht��|�� �/�^��%E�F0fR��@R�<+7�חÑ�B�O>�KG�v�oN��7���B�H�Ej���7���-���M��~�`}6嫠�p��0E�g��J����6��u�:�?�}�#Q?W�.t��	+!��<��^�r	&R�y �*�jS3����������+J�������m� g��BW�n�Q`�T�11bK-����Zh�;&�e�ϮczF���B��
.�]�'�.�M.��|����q��'��M�K��qcx�� .�0Rw��ox�\kՃۂb�Ԙ��L�!r4�3(��7��2��rd�:��CӒ�5�v�.�2�Ozv��Z�*�z�M���j�-o'�v��sͩ]�
�oK㗔�,Ah_�!�(��)��f޲H���VPT�����w�]��k�uZ7��r8�1���J�����آ�4ɩ˄T���5��f}O8���?��֛��'
�Y[�k2/�-h�#'����~�{�A���ve�$ C���Z���85��5E�n������ᥧޤ��M�� V�]��;o�� �8eNv_��_�()J��*����K��-���t�n5?�zV.Zb �s����*|ն,4�ʝ�t�=�#�S�r�.v6ĥA�	R���C�}B.�5���N�n,-�ѻ���Pƣ'fȟ��ByxfR�dм���ŴB$��_���N���J^�9�r��X,.����Φl?U�a���IƑ������̱'�;�x���n����Ϩ)xv0�Ly9�4�ڇ2�w����n��O��&7V �ں���W���+	���c�wQ��*hvLn�����ZM���jq�@�9�D�a����SA-�4��Sgp�!=�
��)�;N˟}��b�9��e�Eq/!s,T��|&���sl[�ppjԕ�i�^�B�ީRV��
���5U@d3�%:zq�=�0��}ډ1��6W��oјU NV�O+�2�/� �����PR����=�D��j�V ��b�0�~������r؝��SE�u�2�J��H{4t�8&${o�f�bG���ʽ����k��U�i3�|rE�����Xq���3��9j��zH.��:�u�ۮߺO"0�-��M�ꨔSI���3���A/O@@�C �JEw��� 4dLw+�W��[��I�5g:8v��TP�/>���G��zc3V�(�ܜU݋5��9!�_]�"���ޟ�M��dNb[�3X�>sua�vs�~��⒤'T��C��f�Fa�a�q��XU�.�����?DB����� (��W�����hz�_zt�����{ɢ֎�пww��l�Ճ�^:h� l��'�����i�n7��s�60Q-��u+�}]�.��_��|�y��W���Lj�v��VQ�V(]�4~�;0��x��m�WM��:�y � �zz,|�,�� ��C��;F�H�9ZB�5T�B&�i���DG���}��!�/��	צ�<|_ߪ�p���2Y����Kj�X���#s�j�8�J!	�P �����M��s���w�fF�^]�H�W�c)�5�Ԍ�Ѿg+���r�|�B�v�5թ��À6�E�^�3L̞��D�*^`�a�)k�ɔ�,���>�񄸎����w]!.?~��=��J��UԤk-�����N�FlO!��!s�L͝�] ���8$P@�?I�7O��P�de�E���NE@��(I�Ji[@^�BU�������jMp3���u���%/�c�L����P~���d�z�0����:�.5���p[��k�K�G����4F*I�W�}��CWp,�/5��LE
�iw��m�#��9ù�� ��7���x�c�0V����r;&��/,W��z�l�؃��,9�$��y@�n3٭HPn�A4N����|嫨Q��:��k�ς�y�1_����Ī��ƕf����e�p���l���QG�\�
�p���{I7�8�N n�,�D���<�22V֪��� 5^�]dWI]��r���>���=40�2g��X�JtR��b�Ý �@D��Z�wH5��W�!� �4��Kxs��㦤h�R
4���� �aŻ
s�41�F\W�قSS�m��7�@�&���f��^�8��Y������EG~����X���:eT[ ���-c��LK^��7<Ql����6�a6a��~���F��Q����w�prBӓ�����<7O�f����@d�c�#%ZNr�$���ұדuG,��g���߂���M�+AF
L(�ĊD��p�1	��ޠ�B�� ��Y�7�.E�Ĥ/���+�ۼ������w��KQ
�����e���X3�>�Hi�u�� �e�˫��xS��	T�]�H�o4N�O�[ �+�4�a����˟���/��*���pV>{OO΋(�h'� V[��%��`�e����b������:o���0)�'�Et��7�%;�JVG�Q�I�1Q
1����yü� �=�o���<��4��J��˪y�X�*���BL�V;���9W�L�yIO�8�ы�$�i�[���^ߪ����/B����D�0���â�ʯN�),k��Tg�c���ʗ�-��\�%mCv ������$�x�b��	%�?�ybF2��[�3��k.#ga%V��hLj��>�8���#��b�y ���_I�h�?D�B���J��gY�ڞk;>��u6�-	��;R�#ZP��l|�P=,eQ(�O�������&Ku~��:�_Q�nE�S��Ł�cdHW�Or�$��܎��bM����/H�'���mU ٹ���	�������g �^^+��f.���e�˵5�4��dE�gb�yP�-��}�5���e���+c}{L)�r}fBuAT#�&�ݒ��@��J�-Q��o_�-���\W��� d
>N�r=u��72�t�\������q ��*����#�@&}��1�o�)�g�.�	�����=�O �>��/��4�c��q����L�<pڙ��[���t������a�9��6u#������o����	>!C���zR�z�j�e�8���~��\���`�_�@�o�P+����Wu�S�4�Jwoc�q���e��'�e�ǲ� J~�h��Y�� qQ�|�ԝ) ���E�8���2����� ͨ��?�NK{eV<��O$+3)�;�eg��p��&E�ʋ�3��z{�|	��q��(�����\$��sf��j��|*�,�ʦ�1�r���&w�R#*&��$m���
=��/bo\��![�����3U�2!�!�#��r8�Ҳ��~vv:R�����j�Z�&�p�")*�֣��^Gv6ʧ-�'1��N� y��|��p���%a
.��_����m]��2�H����EX�����ǲ.��}���[�R������f��j��%��q�V��:e��VۂN��}�d�΅��-$���|{h������P߰C:��;0�u��;�RC(��{K�Z1�"I���e�)d�w��_�]���������+�,���#��eyU��o=��&5��,��/:[NH�)�������&�*B����ꘊ��/n�h���!̬~p��OF�!I�M�/ ��4�g7;1�(�hr���֜
�\��`�|I	M�5O��y��8[��a�Zc����<!˚�\��gl!�࠺T�=��2���!W_^�U��r��
�4#���C��#chL�B�/�(��u�̄ uȁ0��ueVgc��&v���H!�h�c�Gɹ�_�-�n�uA��>�q�P/�]J�n�'QY�c~�Ba�l�@?�
$��{��^�l�o�UV*���an���8�p�vVx���l��]L.	��6��Y���r�X)e~�Y,tc��	��#ĕr6�	��O9p��᫱W��T��N3|uW�"?��y3.����|(��K�� �^�ݲ9J�E�ѥ�+صg��^���o��7��p�z�/��c3h����'���K��1��2)�N��o��~��������;]�Ya��/��:�E��6�p��Q����7L��|�6��ncum����D^���ՠ2x���E�3*hCve�2���)վ;� ��Nr��]F����F�^�SxB/���V ,��Y��u@�>qSA{�m��pmp���_���n"�ۊU�M�1���������՗@Sam�E'��{��f	�v���?��_@�F0�WWΐ�I�qp��+�!����v����N
��1�t�J��#�4�(�����tX�9P����ۀ%U.�\݌�LZy�ӿ�&`>�*ɇT��D�G��{���@@0"ۖ(I/��w�%�)�8����������9f�}'��PY��(T�� zn��XU�\�{.��ÉȻ/����{�f�\ü{�R�>���0���a撰����THm`1�-�������v�*�n��3KC��x��^�$Y��x���>��x~%ջ�r@f+�ٟ5cY!�ad���;���T��"~ۥY�D_4XYwa���?�(��dS[�!=��!��)CZ��=a2��z��Ah���!�����*�d��'˧~%�1�h�Яr,qH����9����<���k��u31�xH(F�c�O��P�3�o��d$$�uih�Pvm�~m'�m�����1���{��k~���,Lm�6I�hr�k��UzF����?0���¨���h�T�i[!�5D�����E���K�V����<��{C#�6Dv�_�>�C'#�"�O��r3�|���y�Y���x�8�Ǵps��K����ߑ���r=�ו��b��}�ח��F��W)b�[��a@���,(Yg�T���a���P��Z&��s���_������+���:L9_ �$t��Z����3?gj�
��}��8$��Q�ڄթp
2�,K#i�cW���@�p���n�ި��<sh�=��+.�����WP�
���?��f��CA���m\9��+��Nn�t��87m��=%O��Z��n��Û�K|��P	�p	�O��æZ߯�`�w��2����K��$��(33y�?[�Kr�V-1�Xn[P.bOk��<����Gާof��:n�@���s9��^��e�ʂ�Fo(3�ݙ��*~�V�݌�� ��� ~u0�a�+�Yޥo�˞`�vEv����U�M��sG��oC!2���Κ��B�*.u�&�b�)�J�8JL��I}����]�>4H^h07×�U��r��n�#.�D~���>����=J ;��Lw���$_��h��\�2ٌ=�I(���~��w"�ۊ�vS����%�n�OpW��B��В<V')��A_���5|%z�,Nn
�s�[�A�ͨ}�8%�l"2+���a°��� 6˺���.����"Yq�ߦ��N�!6u�L����Ρi#�J���A1�p���8��#l�2��d��GQH	>7�ϛ����Ǆ����\��H��Gz�R_�{U�=����0j����� �V������|b��l��m�eO-��J���ݿ��}���'2^��w�[���f>B�։4�ɭ����唖}�A_a���F�K3Z��P*��[~��9�{��&ąO�g8��w1��^�"��M��cV����e���� �)��#|P��m���?"���T���_a�o����My�uCe����y ��-F�L�;��_����bStg�j�9 �b=/�8o��M�+i��P߿~�����X��v/��7�Ldǖ_(:�J���T�W��0�=���ak� 'D,��	��G�W�Z�Ԛ�y�O-/�� ?jSqoK�o:Wd�1�����E��P܋#-�2���(yI�NCu%��Ppq	~_fk�9ΈqR�h�)�V�c~�7��~��3i6�C���BS�@�A�v��9cG`��]�O�D#��;�e�/���/�q��~�E���Z G�vO��<�o�&#�ژ��Na�0�,cC��Ur.�>��bV3�J�R*x�Ʌ�P�]�n`u�y-_Wv�bk��$MaHBb�c&w��!���%���[�ɫ\^� L��=���:�a(��@�h핪J��#�����4:��ߩ\�%��S��/��>e�rnM�	�%+ڔ����~�oA\���e?9_����z�Y�������*�6q߱s'4��f`�}�ɚw���u�@GJ�]���e��o~�Q�1B�&f�:^=�S�3�%�OV��:�H(�D٥��'�3�RO�����	F�wr�q�bٯ$��|�Y�R!�
돿b
e��Ch��e��+]�R|ӘYp�^!������lp��bH+_�v�|]��/�8�yi�h���gw��l&iA��i.��v2D���#�p5ʤd�� ^Nt����[�6��>�a9��A����%l�OFRmڱ� ���o����>�	� y�8pߦ$�V
�kH��%Lpv]U �s�=w�[вd�[ņ{�atE�"����gl	�]��R�� R�;A	�����M���\pW�3j��o�	�%�������c�fV���-M�����4��P�Q�cZ�Z�s����y��b�q��W���#���^�>���;�X�ri.z2�Q<��]%�EN6�Xj-=�~vk��|�]�6�����:��fxR�z�ا�l�225�0�  �o�܏I�X��vhf5��^&Kp��Z�bx�Y�P�'�8��������̸[��g��H� �h��b*���d�O�i��/]����J~��>X�2�HO�L8��u�A`�5�L��a�8��{H��,-�	<����m�Ÿ3�
��c�۶V.�;ވ���<��U����,��7�f+�dʱ������0�0����h��;����n�bi�p�w�~��ƴ��|(\���]2(�t�����#�/�?&�E�]Hϧ��=�9�:o�p>��,�����;�ߡ���D�b��[]�I��=���ڰ�z���i��P�:���l��ջ1�@K�稑P��C1 2-�3"��ׄ�ioB�f����n;�т#�4l���D�;��<����MO���ȡ�ԗ�� �*���C	�W'�QSX1c�Ƭ|�֌����	c_�IZFn\��tz1�P�D�V�$� ��Xi��>I�7��ϓ2��R;����Xa�O�^������v�u�di ���1J�n D59�{ ��l�;M4��_lzy��w�@�,(��o�ev��`B�I�@D�7D&d�h���הUg�w�7�3�P;ܟO-�D�Ye�Λ��Th��~����D��aA�@}2	�bb�j-y|
��6�W�q�4��v[�#j]�H����sf`�/�N�/��#+A�|�;hu��1p&���W��"}�C`�\I���f	���&C�B�}.I�B���}w���!����g.���G����fL�Ł���FPom�éRu���C�x{��3n<Ƨ(
y��;���&fi头�^��]A��QR+�,�����J�
�un��H����D�8�Jb��V���yu�A(��ò�9�Ι�h��-_�ڔ����P���֦ym�&���ՙL��"�8�S���6��ς� �P�A��<��	"Y�8M�Ba��EȰy�_=��
ϡ���xh���a�M~{*,y�(�<b�>��~����]ñ��"X�
{"���y� i
%��Q�$��k���I�20�3\�n ���u<xI�]�q�m���Vb�O���p��ނbkq݁P�ꠓ^q{��cWg�s��9�#V� � <��sǎ��8S,���9\TTk�S��(�h{�O���p:e�#�j=�����" ��|˦�U��]����EJ=Ҙ8���YͰ�U�ʶz���=���9"=�7���*�/��qK*�u���3'��ט��=��|z�(+J��������aH�]�0�0��]�Q��$.�T�h�o�z������6����e&�gy4�W���=�'����"�]����5����^���x�*�i�n�;�?�d��b�	��R2�ܨ��L��4�4�[Z��z��\�QF r�u��i2*��P��p��|^ �On����x��u����M�}nr�x�)dXx+��Cw���i�!L[��H��g��mtؚ�%��_�j4�%gi�a�4��S�N�x��us����:��Ѹ9�-��e�>���b>����5�*�r�fb�y�U[q4�n�,�K;:��� y�X``�gHZUGޢ���kF]ָ�g}5B��xd��U6M�J/�şȒ��I��$3\B����GT�$�]����_��n� +�"�k2R�2s�L.'-%�A"͛�����ꜭ��׋B˟�#����E��jʙ��)��F|r�{��?Q)�.K*��M�I]_W�� �n���-�4�_^�e�Dg^+����5T��QJ��}=i7�Z?�%P�X�fw4��q�+�]R>��kq���<�5v�SM�G�;N����Ii�8��f�^o@��:��<��D�(Ԅ�f�V�=��N�xS܊}澐�H�27��7*2�`;WnB?ʜ�I�)�T��kO]>�%tets��
L�݋�T���;�~�J8�h�z�:��p9'��ƌv�	�1��"���qJ��G�,���9�2����	���P��a�0o�G�K����eJ�Zv����yj	-c�7��80�s�u'KC�7�N��H�ㄅ_��J�㢊6T L԰!ẗ́��)�-X&珿����`�'Jty_L�7���j�!J�ؖ���M��!��[���wA������Q[A�+����aJ��c�o&J��sY�
��J�eZ�_��U|q�����s�k"��׃��5[k{��[/p$<(c 0��9�
�C� �I5EK�L��u��T5�F���,�u���@ i��=�HXM�3�n��V�Щ�꫘x[�k���,�x��MXJ�	˫������R���J���&�%�P+����t�e��k�I!)�@w:�{�P�e�Q������ͽ}�D�2��b�:#�T:H�\RfE���\i�p���/֡�[_���7.��q0c<r�@<�<g��H�'�bnpv^���\rp�����#�Ux�ԭbEai%����(%l��ڴ�=��;J�}粎�'��9!y-�?�����g���ޒ�f����^�@׀�'��{g�NAO)B���j��L[9�s9v�SG&�1�ͣ�&)��j6�����A%�l�`�9C�,�����f��@L���-��K{�I���,��d��_�]"d<�#��sQ�T-���'ζ23��.����6��C����?`�8�
�>-`�Ա۳�;b	c��$� y=I1t�Z"���0�E�9�N�ep�Yu�*I�P����l(s�C�_��
45�jH�<������ZuL[o�u�׭V�'v�U<;�lZҺ`L�H�n�f����\��E�'f��x ��1,����Q;�D#�p��HWHuS+k��Бf�=�=@|�)�L�;
�<H��V�������}$���l�/�NEdJ�p�v�q
���-�H�1�O�����?dg)�N�VYt��Z��)n�]nڇ�����s�;<�+� ݇,I
��N�V�,�"��8Y��+.��:������ΞI�b�O��A��`�>�<�����̟�+�6�%f�r�����L� @�$���"jg�;6GU���<yȝc��d�C�8���8ї(��H+z�_�]0�G��!yЃ�T���N�͎�ΪR�7����Ŗ�!��m"myE��a,<�� �q���1�����ȓ�K���J�L�*�Ac3`l�VDb�������
BcH��R��������x�F٣	/P<S (u�Zzs��t�j\�TCe1,���~��]��&��㝳;�����I�(�8�8i�@��q0@�2;0����&���
��M���Z��ףt����?�f���r.��L@��.t��`�͚c%Ƿvp86R�hy�`J������W'�"����al�_�u���Ƚ}����5z�3��|p{('h�跘���\�tk�U �c�V����|�J�"� J0��Z̡�E�G�>���i�=`��`۬�ϣU
ܫN��di��eܲ^�r%5}�Z�����#<��}o�����,B/^?�<�;+q�&H����g|1X��9yJA���"��b�@/�����������V���U�Ȣy��c��V�6�7B�묮<7�D��ý-�LO��=�ʾ6T��l�|��$@r,q!�Ft�
��G`����a@�	����@�bh�3�S,���o��ZK�i+�6����$g��W���hS���'W"6$a�-�b~ ��*v�}L���m�z%C�vY%_ ~o��2F��}�MσYd�2uq�d],�4.d�cj������q�;��HF�~�zU�����f�����"\C�^)� `m����(�""��W_ ��Zr���r���:z�3nT�l��Z�7����-�󋡅�G�_1*�/�)�`��s�ø�y�N��ڐ���9Q+���0�0��(��-��i5��:0�����ʱ�n�?�  �$���L	@��⣶�,�l/���S
*^���r�n���6�}'f�4;毦}�)�̏�����1"�AK勷D���d���?cH�x`��c�X���%׾�}K���W[C���(x��$+|3N��LZᱳ5�Cz��!�B�yk�$YL#Nszn�9ԃ<`e%j5���W��JG�R��T�'�/�u�![ւ s;M&��'�w������AG�iVJ����,�/Dn#]\���᯹}7����O8'��0C{���G�S�8u�a~&E@��I��8�bft
R}����)���/)Q��N���N���"vøp��6���8� ~��.˘���'�#}s����o0S��W�>a/�Q���K�:A�3����9���,����(�FB�M�@(	��b�N+n�B9,SWNz��0�P���m<����j�u)R��OC�T��&3�!��Q1j!�%&�
�ru($�#Q�=��2����v��c��'_R���ݭ\��ky����|���v�	���'ll�%Q�+ܣP�Н4!����-�tH$���?C����_�!�!�EC�4$��2Q�[�Mr��h9{�h�{6�J$S�^쾧�]^��V����d�j��Dò[o��2xY�0�np?��N�"�.?P����pT���
Q�؛�� ���l>{(�ߖ���x|FV̸�k�6h���/I.��iг����T����P%X?"��%z�wq�;��x̹�
�l*�)B��	A�'�8���%o��4��RV߂�w�i<g3��	<P=Zp�A���܀cg�)r�pl�9Foes�{�E7�X�#�>�ǽ��P.5c�I��5�{�N�Ȓd��;��x2�#��K��m""Ra��_��~&����l�z�o������VoW���������#'>�e�H� ��?�Bޑz�x�������B�ꀘ��Ж��7���m��F��Biw�O����"#W���i�o�)$N�Ŗ�������-��H]�����"�l�w���K��sR�߭�0!�]pݠ���`�W�H.=k:D��l$�͎`���tiA�b�ݭ��Q�I�KWi�,��Rb��.�Ψ>_���� �I�}�����mZ"V�wh��19�f��	Ӧt%]|�Dl.@���K>+��֯��A�A��z%��"�<x�۳���`M�u.A^L"Oe\��{��'8�AY@�7}~�����ǌ�?5m�Si2�Or�e��xbz���2~k�y����6S��T�>b�ob�Q�b0.���c�ZL�=d���f��k?��g��y��t�F��@�5��-�_��͂g��U�,��[��E��l�H(�ӡq�����,�ו $^֤�B�P�wK�"a]�Y/�-�-g3�f�[�d���	�x��?��z^�=��rd�qD����rDQ��0���*̭�{{U{�:��4�v��d�8]Tf�����Q�o����po��`�ؿ8��,�2����I�I�@��!������q�rg7g(qC��8H���I?��8��ۓն��b��d�(8��<��vi�EＢ�:���l����#�B��t�@<{��H-��~�
�.w��h^�oO�P�	sA�-E/em�%o�jh��6x��;� r�� �OZz�s�s�C�V��7�Ūr3�#����
���q1��t9�+Rw��%�R�xɛ,{ZV��wM�#���?��u��c��Vk:ԜOc$F��i�-8VS5�*�Z����!�q�.���c&�.�m<I�%j"Ue�Z)�1Vv���0�Q0�8���1�v.�@k���7pJi�A���y��ݭ�*�s�_�6-_�X�*$�V�}9h��qH��e�J
f��+-�S��8(){M��b���J�@��7c�*��U�f�h�D��ծ8�xw` O�y�Z���E�L�)(ag�])��Y	�'��E���U�R�6��ބ���$�47��������XA�1�j�|�q�#�m{y��i�!��%�WT�)b��#���+>�z��ҩ_�I<���L缾��NܩA�����&�ֻt$�ҿ3-�&��Z$��V^�ڱ�\�[c��r�1K��L��V�&���.U��kg�yiG��ShL��C��9�&�;p�1D(ʢ�R���x>S�ѯ��7KQ
��(���U��ľE�l�K����u�� `c9m��7���`��P�.�nUlpS=1�O�ꍯ v����3���N\
�H:!�}<m���R��i�Kz�J��"�o��G%�b-آi�n�T �*�#9�Ǌ��8����Y�6k;}�����/�Vt}~���cњy���4i"(nV	�F,~_�"�c{�$?B��'	`+_�W�U��Ώe�`�y'�]Q�a񎒟n+5�[X�37�v0 ��ܱ%�G�e�^-0����g�X��%�
�,$�N�<`��t6�{���7����(-7ui���F�>xY�T��a�3����*M�G�9	�aHͦ�fډ�VJ��'Bh���䐼=�-�*�Gr����>ݘ3v��w�ՉD7����a�� �����.�\�h�|L Yk�?=���U'�IY�}L�u,`����� ��6��t�_2�)W��8�<��#HJm�&�|��}�{!B��L-���	�՗-�X��:�[<_D�o�N��8�+u��4A�F����	�#�y}#щ���BmD�)�^۔���="�z,�U�a�	�:I*ye�u��"*��s�[<6�P�B�+%%�R��6C�58 b��u��=0���n�xR���=�S8ʝ�oS~�����y�����3�z�����/�0o�(�̋E�#��<�v=�������e����ƙ���囻`��{p�23~Kvx��I:U ("�üѱW3㤸��BHD[����|+
���,*�U��S�lY��5 �$D)4c�&Yj��ݾY8�
��`���'!��e_m8�-{*�%�=��$1�SQ�=�䦨G��b� ��\:!t��t����Y*���*�W����o��m%��'Hə�v�@3��!�jh�$�&Lx��[�{���6ñ�;C}��ޜ��m�-�~��yi�T�Q���C`FH\�-~����_=��7Kh��,��� t-�ə;^M;]ڳײ�^E�Y��)�+���Q��Pm��Q$�R�G�ۆd!�҉�5�\Q/���M��๸�J� @uʔc�|l=���[~�����W�Qә��� �{�Xj�X�'k��$y��ǑO�����n�4O頢2�֮���b.z�������O�lҲ�<���w�9�+�%��R�ִ��\����1�Pǎ=zrRޮ��)�yե;��.��������K�D�+<k;sG�icIP"gU[�:OD��'���������݉�a}�mr��yc}i5S�|�:8)$!��`��%%�8m��Xb3#��J>�$�5ܟ	����b\����"4h�vŪ��P~XU�(�N=�|�5���=r����	��3��yW�8馌�#[K ^f�÷@ �ig*y�U�T]|w�V��pErt
u��N��/ת�:{���Qb��9VBL�	�֪}8^3��������cK�c�~�Uj2m�������u�|iI�L�s�q���og�JU�G7j��T�h��Ǜ!��`0Ȼξܵ�;{�M�<��h�7+e�� �!�Q�#�
a�|1Z�ˣ��3��Bfŵ�6@�q-�0W����ʺ>Հx�U͈��}N�^ɖ":{�k ��9��BPA���s`_�~f0�P�b�lϔ��ߌ'�PM��L�T5�𰣍�kf����e��AO����v�8<�3�~��ȿ/��.�������E�C�$3��5��@�olF�؅�.��S�Cb�2���m=R��/�� �H]m�3FD d89�	���~;������	�"�{@s}�1�YF�<�b�on[u"w�7�j���.��sI7"p�>�r�� �fX��k��$��,ײ"h$�J?�}e�򣑠A]�U����~�w)�4�ۤ�8ǚ�񥈫�6�R/�^f�c�����U��vG>A7yZ��3jS ��p��Y��X��v��X�询>\�_�⸩S��~^��ngS@��G>�/@7 _a0|�v�4��A_�ޚV`y��u�~2i�{���#�=�F��{�h����?z��S֯^(.��h��:y*��U8ٻpH+o�
}蒷-!j��s���#�T�������Mxt��m�YK��U[%*�֋fu�;SP�	}�k']��� �H�0	�x��v��0� �x�dE*v#�@g�O�&��<m�iF�=[�֨���0�A�U!D��@,>�S�m߅�$r��֯/F��;~dpΆ���n�DY������`�b��V=�QL����h�>t�)Z*۽p`}/f��؈t�ǃ Z���F�K\]`�����v;Zs
�k5��l_zI�&s<�_̙�q�K���	�� �А��>uc��b���?=Kf���z����-"��6rz.�:u��\��.�3\�{��\yf�� �Å!c�5U����ɝ��{T;��uVR�3.a��E�C�h�� M�%	a��W]��u{�V���D�ǲ˟!���\�0�%��q�=�vۛ��	ڴ�+��j��R�t�#,��%�Ҁ���`�Y\��(�/K������=Kh1����C�	Y�1B���*٦�f|�]��m'$m�G���*��yJ�6H{á�;P;H��K.W������n-րqf�\2i������ٹ<�1aϻ5F��K���ԓj��f?;�ܵ�XZ�P�����+�3��q�ga�MoP1ƾ�y�u��F��0���a�b\_P.�:����X�"ǯ��b��^X����Ġ�G­b���gL�ֶ�ϒ�#�#�N����'�13��e�o�Th����NA��@�6����Hh���l���,�?\uz�JV�4��^YI��A=#1�Ix}go#��j���v���WK�uz�g\�H�Iۓ�S ~���kT�5�, L�N���B�k$$��v*���H�nѨ5���q�T,�r�'�Ia�(�1]N������䡭�f�0�!����)���H7�����!"C�ɩ_P��w��W@V2���Ely�[�Bi."�����pJ����d2UĖӚ&\��b�b�a��I<�L�M�4�2} lO���c?e+�12�J�k��F�Ƒ��]A�,u�=E񾮡hÑ��bǲ��jrb����QC�0�����_�,�V�H������Q/D�R�A�G���meا��lM0�!�Ŭ���T���~c?�����*P<�ζ�Ht�7���(h����s*���F���h�}�4�w�-⚋L}���ȍ���z)e�P���Pu�n8���5C?ͬ[wجJ�jMSZ���Ȭ���KK��}Y��FJsi��'H�T<�
�M~Ɉ�(W��q�ٓ�>*�?�ϖ�.:������Ju��灵Hj�a?��E��4��5�)�J��j�TbRK�y���k�$.������ܣ��{U���&�=����Cem�~��l#ǂ�'G�����Rbg@Ӎ�Y+�Nk�BHy�z���.��VFq�;gՠ�'��I�H��̉�߇ŋ�6�	���p)6!X#znu�l��o-��_zt��6�)(��GE���lg^�ڝ�����K����s�����0�4��Խg��A}P2lF%���a�.���#�,�
�&[��K��g�$&EQޖYf��#*�|2����@�T����2�������s��ً�g6���zka��\�IW�Jr4���&@#�ó��arǖr.�&�B�)��td|�;���N>��!s�L�9jUB�7E�-���5ar�y_��B��bW�^U{5d��|Y�w ir)�R����3������������5Z
Fn�'ڦ|������?�#��]@WV闩���^��2qhE�����bA������AU��4�Dö���2���+�"��YX��C��2ը��Hmu��XY���N�P??2�tS�@t�6�[/�� �w�(#b�~��9�A�<��ry:i��:X6f�T3d��>��5u�J��H���-"��"x��x�d��P�'R�f�`<�W����K�� F�i�\���{oQ �2U��t�ܪ�י�����{NG�p�ܕ8��{%�<O�BWpbr ������YXX{a����ג��C�;�PAe�u����8+��x�p�3"��xF�O#���q���ͱ�fkc|�%QgKb��I�h�|P^���i#5Yl�+p_�F�!؎�fxn{.j���e{��Tt�h��KF}I�k�@Q�y������5`e���2�9̋VV��j�Mٞ�}�U�C�.~d5x~� ��e����,B!���}�y�1T	�ݹ�+:�3�[�SX=�dzQc�$���*��P[��o�4�n����:`,�g�u0f3�Yj���k��'��Y���k;C8�&�!HnC�*�5�u�V�kET���
�����A�\f� 0��2X�"&�L/�l :��B�[,��rɼTLv����7��`�k��O���f����S�������yQ�^��o�p_u|)�K����n�h�]��kl��
�"�e��d����.O&}��LZ��"du~������i-�Mꐔ+�����`Tl���Op�6�zc-��l��x�Z���#U�� \AH��>I�t*I�T�E% �h+��|�9\^������7�O@	�Գ��[�̫#dL�o�@ԛ���ՠh�&$�[���?�.0���<��r���+@t������:^-E����98A�����\8����D�@�M�� 今�C2#1=J��mrRN�GSɗW@�/�v��9n�ES��r�*��->���%���e���$,+\���cI��|-�&��5��\!�t�c���	PD����NC��	�h�U`}�Z�7�9�Gh�������{[/L���!����½�u�S]���_��wR��
2Q ���U�T��6e��Qyi�3?et�S\�σR��sK2к@^= ��e~3)=Ў�X^s�L:�~E�wh|];�^��8�[,
u{f�s_����D�m���R�]�e���̫��~J�EC��OQ�G��q�@1V�� ���s��)��Ԭ���r�6�����Bcm���4qC�9M��5�1M��x�q<ko�������Nui�Wт`�g��]���4-*�+�Q�Q/�z�q�u��`��ΙA	?����G��"Y�z�����=��������<�B;�4i>��p�/A����"o��z���W�R;2�@�x���8
x�ּ�i��bx��G\���t�	l9O��Uϙ+�%r$շ�x�>3��N�I�be�o��Y���D� ��.��T�,�R�kЯ���߶���@�������|�MZ�L�!��@��7M�;d�t�:������%���(��}y�{*)��8��d�� �)H��?��ۉ{~$
]�e��s�dyc��G���v�#�Ct��Z��cZ���[) L_����*W]�ކ&wQ�0���&ፃ�a|�������(�m��<��0��9�6��~��5[<�~pX��Dȟx����1e����Q�u7	��OC���v6��z�2�b,C��U�P��Y�j{��r�A ���ai�sR�Xts��[��>�L��$¤��~�T��������53�8f�>g��N��"�C��?��x�؉�c�O��p���"Iȶ/N�5�ld���2�!휶���b1�05s��=.u���Y�9�w�:�j����������}����&q2�&5O�v��������P.X9ԁ	��t2�J�#H'� f�M�!V4��%P�sB��p�ch������؞�評o̿ڒ?��YY�p��G~w���Z/L��)<Q�eD���	����E�.���͵W��F� ��B}Qu�����ɴ�F�%��Ih很�Ӆ�Z�L�S�U���ŞՕ��gSBo�k2j�(��n�C�n����S�ַm��v7�{B�.&�?�k�\T*2�t�'R3>j��*�(K$f��\��09�6�?#>��&�o� ���� ���_o�U�Wm��좽i�'�N:őel;/�>|�ek~��Ƣ���8҆Us��E���w ��O8�|\���2(K1�|�e�y"_&��������L�cLQR<���Oj�D���M�1���Ɲ�~��*�tj��=?�"C���?{߰��#%����i
��Aj���7��XȥQ_Ro�`R��ε�� :�]8������Ӣb+�iy<�xBs��FsJ�T�z�\�ڴ%�0�~�4e�Q_ݳ�@@��A��z��ou��r�k}rR�ɘ�dN5���Yz��5�mD�*��9���� ���_˻E�Lw�P�H�[|�r+Y: M��)9�w[)�i���͏�UN�s,��O!����$%e����p���U����qޣ4��M��"m��9%���N\k�R�� sn;8�3��1H։N^�@��i��N�o銴D�3���)��(�	�b��(f�$8�#���ZK�H�ղ=����U���aKt�qXj-��|<�S�����4ނK�Sl5ʦ�V�=A��XvaPwNFW9����s}�&�0��ں� �Aj���c�U�F�693�z�I����q�BS���D}B���}� �U^���]�&�ݮd,��g��
�T�`}F���6���r��C��?ኯ�&?�I]���bO���H��ۇ�¹i�3QV�Q�xA�9	]�c\ +� (&
�i)�/�^3���=�o�Wu_�RV~y ]L��0���G � o���]8b�O���hM�:�"X�F$l���5����v�r�ayt�������l��3�b��r��~(c�zc\S��l��@T��/�\{\��M����OM�/J�7޸EU�P50.��hf����|�CF�x�l�mղ��Rb��ax
��:�����T0t8K��Q.�Y(�>{2E�Ab��/����TUmE��T�����@�2�S�U)��n+s#�;Ͼ��J2�����1Q���M����!��A��"����p ����Pvd��������{�M딽7�����r��RO���됚�*.��fs,&e��v\���;������qX	_��l�J����8'!����lP�s$�F3(ɘ���1 Q�"TBχ�G�-j�Z*�K�X���[J�`��D����u��!��jOB��M���s�Oj�k*�MAjlv��?az�e��״����5{�[�c:(�m��[|���s��d��)>��2~�`�S���rae���	V޽a�~s5��ĦQ���=@��t�0���'zh���̶�C�֥7�@����$L5�!"�@B/P��R��w���;� �5g���p�=�HٸJ�Z��̡��oU�S`0vl�5�<���qp��1;O�=k|�]Y�	'�w~�H.���[��_0aTI@�\��NR��Įn���^�85'oAӎ�%���!���ج����UF�9��h߰#u{v�7���
<D*:�0e%Ƀ+H�l�Ď�J��F[J��R^3]�����eP�I����lm�0�߰�0a��� ^������[��`\m���]���^�Gl9'e�V�Æl�PW��������ՠ�E���<��L��4�:O���;<��ü�UD3צ;����RE�c�Ѥ Ǹd.G�H�!&n�����~�#���ZSq�f7�7�t�g`���vÅ�͜)	�b�]a�Ŵe�Z�B;~�I�5|��=�Ċ� �+Q<FL층O����=0hۚ�E4'�����s�єd����B$#����
��·��hۚ�V�+/��9g��y���JV2��u0��*(��P��`�n,�����_P��۴��� ��:��~��NUj`�~ߞ��#�~��$����6|�Q��R�G�?-6Q�d���o�`3e1i"X�����d��x\'���޴��ט.r�C�BM<ȽU��|Y�9/Yr������!Kb�Yeˌ�y"��vOJZ>�����/�=�%�Ls?;�
���,W�ft6s��W�o����?���W�]a�<E��/��۰́�뷸�͙����}�;�hmn&@ ��-&W�!2�6�Eoj�l�is����P�߃���m�C%����%��������wr�M����]@`�G
�&����x����s3�U����}5���&y�Gh�H�#��4���f眂M��F�g9L������#ί�(���T���֜����wd���{ʃ�Rs��w��w0#��0��r�,X�)�pZ����c�ƻOR�@�q���aY;�ǞM|�!!���Q�~:���D�1!�G@R�Cr.E@��H�� �l��|��ds賿�G�	��&�%Z#F��(���J�b�s�}�렪!�4'�+�K�?�$/�%�
G�IFRo���{͒���[/9�t5|C�͝�y>~-�ӏ�[�n�՚ ��<�&�*���]��d��x�p˨���=��h�&{@���������r�/?9u��4�Ur��b�����4����wB-�|�]�l6@���_��h�_��L��J�E�C@����7���c�������$_��JӚV���QZ�vJ�O����!�[��"#a�E�"�s��B��3�B���mє��ӰE�%5ޚ ��	�W&�����a��U��P��/���
H�%���n��gؼ����҅�.[�:��qt����m���M���Q���3D+���Jd�p�9[����{r�>����? �zū�$��4���P:�*�Y�Ŕ�2�c�e���L���k�x3?Ō���;ji�:��=�_��*�t���),j��P�IwR���u���g����`��n�Y[ÿ�#���I
�t�?���|�1p
�uX`vJ��Hj����-͆e��T�1�.��OBe�T.��������@�HW{+���,�%����I��#���"D��������J��5��)�#+��@e�l�J������G�@����zٱcrc���P^�B�h���,�n�Z�&�.%"hk#����0O<�ɉn^��K�I�c�Sn�Q�;CS����֪�41u���0��p?�ƂL�/؂��7���H�'#�]�z���&�����:X���_ ��ĽD�'c|��I$3�$�)���~k�,��G�6�{�+�,#��pf(>9�����m�̑�b�J@"��Ήu���,Y�	�k@�l��=\�a$g��_/7 ͖�/�Ne����x��?j�Y��
�{Zԡ�ݑjX<�G!���`�2t����-��i��46�. ��>��г�K������X?�TG�b�k:3�q�d�v�9�4wn8Ƈ)������TC�3Ҡ�t�&�/�?�`�i���e�#(��a�������z��ͨ8sP���
W��.�+8H�g@�Y�k���A��:��h���Hg_��qT��v?��ū��8����?�Iw���./Ȼ=[��]"��	(��%jM��c�X��<��6�۷�psV�����LUn�a����İ�7)ď��� ���R Gw�	U8)��T�{�����xx�eG�$Q�ot-#N�j���<�'yC����Թ&y�2�_;_��P�	��@X������51s�蘫I�*:W��� ��6�ZH�XTُ��:b4�s��9�C�;`N�V;#�&$ZUUd�V<G�DW��	�]߀�w�\�^��9eϼb~Z���@�9U:�\:.,H�?{q��ʾI�x��=�&+��N��?���}��k�����t��R�s��k	D_��{J��VD<d��Bd�P�G0�F/f����p��T�H`P-'�@+�@=V(��f��x�#!�j9�_�j?�raNj�g^�+I�g�?O�y��^&�� WW^Sl���ɚu����d+J뜊`�n��0	��z��@T0�����Xǈ`�Ƒ^i��!@�*��@.F�]�(�Ӹ�,6�pWbY�$����,�($��ǫ��3FF<��	�n%[��B���0K}���5�Ֆ��?߯K�}�{�ds}/�sPh� m��x`<_�����!��i/1�-?�P��,Ee1M�������5}d�cN݆Bca��̾�x H ���0��yؙ빸?0��^�8h�|�6��&P�������u�	*p�:�8:����� ��c	_9�@KW<�'���C��������M�
�Wg�Э���H��X0`����R��̊���&
���NYo�j�Н37V� 	�q�n=+x��0���,qj�Y��;���POlu66�ksW�o�|ݨO���@���29�b�5�=���5Nd����C6�H��)=u��}�f)�B�l���h�f	 ���g�3M,�,W$�����oX�0�}�˩�����$5�{c�Yj��iMc*�%*���B?��P�P4�04��B�o���CB�Ç�~O�qk�ҳ7�y�0#U���
+StV[m`���`lv*����q�}��1޷/�!<=��a!�ή�^�w��3#x��ԸG[5d����^�k�5=�4�����Z���������H�S�͍Ƚw.ݩ�aM(��?������7��b�d�s�R/�-з��!�+���:�VKu����@>˲йa2�C9#���a�S���26�Cz� 7�F�c7�ݝ��u�^z���x"�������B�5Am�t
<�+9��7Y~�W�����f��
�/�h���aZ�FEsW�Wg�+��=oA������(n�p��(�������r�R܁���j��I,��z�_e�[� &M��i'��d1�C~����c��.��|�^�9����j��!v4���8�:`��\�趔
�G���uƿ�)�؋K��f��zڞb�a��T@��n�,���T�,��	&b9���Ca:G��qc��$EʗF���uW�ê�j�+�6��� O�F�i(���U}����D�sq��M��(c~���I�E_n�[nu\�f)l��"ߔ�nѲ5�ؘ��H��偍ͧ�j��_��%�J�!)�N$��8��X��x�~�BM�u�Y�JS⚿����|�qѱD�!�޷���S���ϩiqә"7M�KC�%�a�
��p��<'8��8�e��>;Z�ow�������]�N�3���dw�&i}v��َ���?�1ܥ�|G���1Ƹ4cf�'#V�I�4�հ-� R��%�J��5ha��*���a�~Fte)Kb�6��w���T��.{x�u�WR{�l���G��Τm�?F;��χ2�i>�S7����t��?JU"n�v��N�Y���+�9o,�&���I���(^i�X1�3����<ެ��=���΄��߳��8����S����cn�M<Sx$�y�,]4�;$���X��ߢ�*B.n������+ЌU�6�����!-��꽨�?Cғ<g����G�1b�����aw�����+¦���n�'��Y%>U<�_I��oe1[��m98$hi��|XQ�ǀٱ����iI�D�����4c����,琷]&	�9qB������U�i�|d*�do�ݠ��,c+z.M%>��	V��*M߬�ϑ��f]�뭥���̀��"�!��QS���Vq���3E2�gI+=&N**�#�wO��	F����e�:s���:�8ML�:�܏���B�S\�BU��D�_����,=���j�F`��k�A��܃4K#K�#��c̗Md�b�>��.%���� U�v�֖s�~� �貼�e�)M��ǻE�m���ƕ�צy��O�P�LW�����P!j�{���$y��V��EǆML^Fn��]Qc!I[��y|:�@�)i���z�jT���H��Z�e(Nx˰g��{I-3��5��{�mbя�Ј�u��jO�߮�+f��ŌA�7��;����t[N�8�]Βn�.���nnx;�%�9ԔV&8����k����0�
�TWK):�¿F.'�����DTAr�嵘�]%󓴆�p��z,�*?{����Ċ $�<l-(�+�x���QW/��ɔJ?��~z�캹�>ȭ��T)��+�K4OK��VzV֜�^��6b=��	58������z�����G�ǁZ�[h=3r��R�Lo���W8m�>�lY5Q����ӈ5*9�<�1�c�'����J���;~r	*��<r&2�)\��Բ���Ư.���K}���A�M拝��w�4���c}Ȕ�C��G�S�1($�dM~ջ-��WHMJ��<���_2�@�}��:��"��=O���|�
��N�`.���j8��!�O�I������'��[p�{Ӑ���N�.Ά#5���ܭ��R�b�<�M09F茟)h�lR�����ghP�Tt�s��Z �1ځ��@ ��N�z>Sӿ[y�OV8K`0H?ru�pa�OnL�T4'�� ��F�[�'�-�ő�W��Z�w����*�{���$��`��t)�������6O��(����}��z��"8�����pa��jd->�d$0�}B�`V�qq�(����[@/��l{{E�Y��֠�5�@��?����A+*E%x_)R�R%h/B���Q�,���H�1�)Fu��?������ɓ�I΄�� "쐛N�4�82���=�Pp��[� �i��}�?��!(�E��lK0�,��!� 8L(ny��~F�'�;Ңp�;�;5��j?� ��;zF�v�ר�D��6�a,����I"a�Cp/��G��xmo�Ua��a������I� ���@$��ġ�T�=,�ޯ}�R�p4#�q���U�|1�(A���y�QK/����#����qR�U��.U�(��/�|�6va��� ��V��O��@���~oxN$a/R[,+!C�U���ZYO�g�Z��u>X�5�pH�L��>����\�1�W�D�Uv��Y�)��"[��_�m��:���M�6������7
=�3ߓ����g!���"KǴr��Q���k�t��l�OC�iH��ݒ�?�C��!�����٬,:����QAejѥ��=�)��5�Z$�z��o�����v(���\ROb���OHz�wwm�i�-����n�����."&1�r!���@��b*�o���M,��p�	��Ċ���-i��E��4�OK;K��\z��B�OCt�rX�� �[�hL���#֖#0�,s^yͣ�a�L/7xE�\_��I�>���˰h��O����m*,�+,���$�j�L>��U$Rǖ����(_�Vё��<��o��uK*0na4��P��3���8����J����/
7πj��%��e)'=��G��aٱ��.����[���9��� �ஐg��JDoh}��������3=��5�'�;tN�pD]���-8�O�[d� �YMC�uB<�D��:һ�#�#��,�?_���B��4D���\��&�{"���%����B����Q���J��kW�&
�G=�M�1l#~)��j���@�*o��!^��^
� �~���d�/�i�-%�ߙL�g]&Q�����O���>b}�ݫ��M]4��WN��۵Z���ޘ�R�kjB$���D��B��A��K�sH�t)WOS�	�q�f�_�4��=e��{@^��ʮ�=!R��M8N1���B#�Mk�?fL�e��`��n�irVZ�iP�h���nZ�/��:��IU�C8������p���cg���K�P�SqD�]k��?����,;��k����Pt�w��P8�[�gQ���X�7�v�%�!`�8*�d}5�#�aHN�8p�v����h�]9���Ґ}+[���t*[�!Ћb���B��o}=���ҧ��ϑ��5�4�t�b�{�O�䵒�\�Ϥ�-I|��1%���u�r߮<i�m�G���I_�$^_�.��󁱪�����fy�x�xi7��Ji|���a�:\ۀr���Bje20F
�~q���Ҵ`)ųJ��
2!�*�A9�JZ���+��e��D�2���G�!�a��t��loe�9%��_sBt�b����D��~���ς7��S{��rj��5�oӓ5}:�Joq��w5��\
|�^S\&Wz���-���v�<���|C���p�A�!�+sy�*�xs� +Nqk\)"w�\�=P7��ͷ^�=�Iӧᕶ�,��-�+]�J�/nF�%��C����D#��j�X�w�'7���ݻ}eR���*09<ӣ����ڏ�K`6�9��SF�u�G8nE�ƺ}N5"������a�{��N�QGG�P&��l��۩�_d���K��Ne��(�����!M?�3�qHiji�`��=k�m@���HP��) �V�oFWW^^V�'�ju�$�`xa���+��@L͞bJw�>E�������P�3ބ�U+"m�-�ʾ�4���'m��������ct3"1FG_܎b��'�����'P��<�VΨ�!;B�v�o��J0�R�ց�oK�g��$���
������&�sK#�2V�gN�6�����z���*)��mO�;AW;��8�he�m���u�y���h�?fV���Q
����i�m���Z/��KבּG�xn�TA���8�/#�خ���92>�r7��M��c�C���8�	��s�H�.wO�I&z�����#�+mm������x>��7�rw���fG�Z���U���0nH���-��oⶵ�KP���M�k���ϐD�b��.���
>� �TWʏbÇ��y<j�9 ��Qh�(:�2�,�c��蹇=�����	m'@}��s@�B����O���о��^�,�6Hn�;�׆�`��~��s�����hڼ�d�("��)�Ǐ��v���t{�|�Nl��^q?�m��/K1����x�
�.�<&�1�%���#�����W�ʫ����Tm�����+WXlh��Y�N���[(K؟a�l��:��5�~����rr�12}�1Uv�8�����y�]��f���tp�=����"��,\�]<��D����!%��<)�Y�o���� /M��_�����ڸE����R�6����a{J�>���5�G�:=�-��'�ŷ�C��`C�㡵贷4)O�	C�r������P���� �y�[�j@��%
���&d�;�VҚ���x����#r�Ǟ�܎3��c���[�˞�>@���M1RJ+ᕬb햶�O�қ� �3igT�����q�ד�m՟	"{v�ۃ-�-�R�:㵜�p?����O�>N˱��6<���7��=�tt@2D�Bɴc��������D�c��|'�qM��H�Ӳ�RjEap�@S�z��$q���1Q�ʔ̴-`�P�C�WD����Hؖmw�d�$|��yT�]����(}��hڋ�N��D����!������YH._�>����2"��&49��}M���&���������h��I�F�#���Y�W�}�y?�۝yZ�W��q(�!�*���<&�V!�B�9��}X6��
H�'p �u.E��^����ŵN����\���ݖ���h�쯝�T�t����8�Mb�s
/���E��X�#��Z;�JV��4��M�8��P��.�o/U���
6��y1_DI�,im��QV*PY�&������^��!���I&�؏��"Xg9�Z��M��a��n����1i�ɯ�/�fJ
��ق���,���0��b:^>��+^�QЄ 碕�<Jv8����Ӕ��������Qv(ဏO`S���hS�qp�tdi9�t�.X� ����[z�2źp���<떁w%	n�>���K��8�S�bkŦdXM���NR�4��4���g�C�Q���K̕�*REr,^�;	X"��:��F ��B�`|_�P	�
�)~m�*X=G�jv���J�1"�fVu�}���@�a`>Yv�*A���URI=zES�A
�s��t��Iڃ���b��\I�����|�
E�)��?AIU;�ø.����y�5�)�#7v�9	E��Msh)W��������@���H���s��L)�pXf7q�
��B�K1��5��j"Gf����%�GӤ��f���L{!I$�V]#�*x�X�� -r)�h��s�k��';�E��7g���>ч�_��U��ZF�-u��WR\j�����x���x>�����f�=;ҥ��Ky;:�+�o6��Xf��u(��mQ�{����M?�)����L�f�K4��0�����5�EΣg��7�9L�b���"O������I�`���u�
����=8r�K��徃t&����2�&�\����g�k���zm�~�������Rn��il̲<u����y�8�{�����G�B�Tu�!��p~qǶ�D,�w�#׬��g���j����P��_�c�ޤ�]�������ɧ��/HJj��~St�N�s��9{%g�T��B�Y@2�ȧ��4@Em�MĖ��yr�Mi���ChxvX;Joq�UQߏG�s�82�^��oY���:7N��nTǼ�J���˺�S��@��OI���t��l	x�}S����@���k��5�ȶ�
>5�Kꚛ���H��.���C��\6RYu����	7�IhC��)��E����@s1��t�=i��0/a"ڥ���m��ܜ�U��h�w���L��CDk� �}�b[�Lӕ���b8��I�9�r��Y
�g���+��_c�KBm$,@��c�^��C�+���������q�+WAk�DP����'nT�'G�ğ���FQ�[�1�'�эC�i9�G8Y��s���~�MCML�cj�س���z�E3frm�q��߰�7{H
�7�w�e"�c6U��Jy!C%��, 0��zI�K�"=@Ћ�R��h�Y\�I1��r3_��#!�F{{�ٖ�ZZ8�ty�&ce��� >��u�ToR��r��v��|�3"���>�Á%�;�yZ��x	�����:�P$��u��|r���0��
�~�� �t&����SJ�zw�a�۩Kx�bj���^Ok�ԇ��u�,Rc�^�x6�RA�1�ң=�G����P��-�#�`��������-������a=��?�����?�R�f�7k�*�f�k��n�b���3�o���ܳ,�C�3G���d�����"3�h�bx�*�����y�NxŤu+DY�%�SHo�_@�U^J��b5X�n��M>f�`����$�k]vN�������TM]��C�Fp�����M<�7�����`7�W��0`�agoC�u�nY�D�B�z--D\�)��>��k��O={n(j�4���: �𡄈&�t@�2�	���":�K���� ���e�r}���T�I0��֠w�Bqͳ�k{�`��L��{��FG�(��-�>e��Z�%V��5�i9*�4�-���Ú� �s@Vy��ދ�������m������؍k�4IOAl��<���}�wN�_n�� `P�P씿�%���,cGY�Ҫy�R�n�"�a?��ףb)P1�_��W)ٱ�D *�;1�z'���C�{	��x�[%)�t�&�Jn����/*�0�d0�������l�≲Úw���'�.�`�y�6��,�Κt��{�`��_�� ��X��'c�7˧W�Q`�0�.Lw��� wn��nx�7qd�I�^{(�Әˡ'�e(�˶��mx�6������(�n๼��$��Yh�8�đ����WDNq)�0�J(��=JJ_z��e1���Kz.��˕�[�Ï�D����1�g�J'� �!ʁ\7��A�M��f�t<��an�aݓ�o�Z6���]�-d�������K,�0��ZN��\�Jx���g@~�[}}��E:H'����A�~�ٷ$���5e�˴��(	��m�%�5��9��5A;����W��	�E[`Jn����U��S�N��=���+0l�B��e>����l��ŋ|�?�nwWW"�h��:緉<�I36�cq�!��f�"����T��$����t0������}1�W�_ FQ����.D誼�8�oyi]##"�~�"'Vh�V�g����$r����7�����wO�Whu���XT�$�d��ta��b}�| ���K9��q��ypW�޸[v�nt��z�#RF����8g��;����0���빪y�7�`OU^�M�O��m>��:#��]�GQ�f5�Xd+ doyx��b�r��$чL�:`�@8ղ��)U��g@ڕ�!���,�b�	��cM�s��:�[/�YO俐�>���-��ʤ���t�CV��k��F!�����$J�z�.$tx8M�om�PH�M���A��:�ゔ ݉8w�4W�bz� �(/���h�+�bZ�`��i��}��9{�"���4'�y��#b�u �/^iZ���U4ȿ�QT]�Ig�|�lX-� F.IĲG��G�"$����v�*�Mv�!�Y�'�`�-NY��wZ5�4�y�q�#1aS��64�+�\�ј���cM=g���|�}js����u�� Q�t<��O׋�L1+ϵ�L�]9��ҙ1��[�|ڠ���x �������\���
tP��AZ$j����P�4��O���KMW�v��9H<ճ�ۯ�H�	�6Hh'	�u��8�	~��~QbK~�%ރz�$i�q���T�7�� nb@���� <�����>0��d�|P�?A���?s�L�ux�<3��u-/��Рq|.�Xm��0y��2����4 g���9�l�oY�)�x�D�:�$�&��V��d[����� �7��	#[4zH�/4
S�������(s��h�\8��dB1�@C���rT�5Z� s1~����j�Ӯ�P��X0����Z�gG&�Q�>f*?�*(��(W-�b%���;���֛��\���=�'BT^A�����Ξb�=@@���Fm�(2���)xg+�1�Ҋo��o��Vi"����&t��`�q'���"͚೪%�V��0d�o�:�^��%P��{Y�zCv/ �t\e��@m�є��z؞�8�͡,G�f����?y��w��|[��ۯ�CޘK0�,)�-��6o5O�z�7�,g6�ٳJ+V�y�5�O/K6B�� ��R�Q1.����3�����&:}SH�*���5�%W�(�7y�,����AUe��6ћb�8$fUM���.��l/x ƫާ�@_Xi5�C�	���6��[�IW��o�N��)��dw p�F��I��
e��q���(�{��
 *�����r0q�M%��ϑ���Y�Y:8��]p�<ǱW$����+ӂN@;hP0 AjS��{H���Э{�{�[X7hˇ���'Z%�Oi��Dޣ���Hs��hd)�_+[��,]1((��X�^�JK�:$ymIV�_�����3:�2�������H�=˽�=ja.$���3��R���_g_�$|Pҡ�a��69�!c�� �mZ{KrM���ͻF�J$s %���#FHl���4�;��Rp��Ǔ��hIU��:���1���	�xF��Ub�����Q$YcU�g0���GxE���H�g\
��1
�4�u��%N"B\)8���UQtM�h3C�Q*`l��-��� ��g3��x�����@L��­w��3���k;�gd���[�J׸Q�7#�q�鑆��yv�վa�8��b)6!� ��D�a"Os�_�ؖESP��B��.���e����#��'Rǅw�i?��q!��hBa��y��M$!f����8�0S�@[*�Q�Re�8y�m3x�ׄ*��L�]t��pe��_<��S�@{��D�v����P�M�۱�!a#��^Y�GOQ�H �!d��E9
��gX(�6�!���Vx4�Q��d6�%>��<x�j���j����Wv�<��Y������-�qU3��fi��	��9�O�9M7�.�l��8_"���W׬�F��P��x������T_1�*�̝f���inud�S�|͍�F�!,|�����B�Ֆ�PN�9�5Ч���w�"���m��ԉQ�W��խĒ*�E�sǖyE�%�oO^�̋�낥=�<gϘ{Y,�D-���覤�p�2x���#�JM��S��J0I�ҡ%+�c�A��3 �˨L�^>0�E�`ߦe�=o��6N�����h����◦	)�j�\�����3?R�H��B�~A���[f?yp-`��U�����0�c.V����� ����	)�`cFidw�/�c��}���s.Y��r�wOrh�wèA$���19�
��]]�f�#jB��s���E�$�,~vp���(Z2���"��c2U<}�Zf�fq���YJ���ò�Lu�sF��) _׬tQ�N�1�N�I.bS���'�=x�ι�=��A�7�@�g�sNؿ�#�Ѐ�h\H���5�Y/ �<��:�Ɯ\����
Lh���֓ܮ�6��~�;'И�oú���xZ+��k�����A�*���a��`��)�1�sm	����IVB��E�G��JMz:cx�w^���1̯ťi�l��Īm-��b'g? ��v2�i?�;AE�{��z;��&����jԱ�<��m��P��Ы9͵������u�MFQ�J���KI-�3r����)�ks��k!9lՙ7������7[�q��u�t�SU�?�<�q-�v~� �}:��K_s�xyE�vP+pi/�ul�F���R��duQ���� Q�*,�d�ZM��ѩ�7�@GT��*�1�?� �r�Y&�>v`���K�T����n:ah��<��+��6�p�Ң�gqg�q���*�@	���s������Ŀ��+:x�7�A�c�Yu�Y��L�{{�	��X8�����u�X��o�Hj����7�LS]V��]x��?��_G����[��h�h"cFIf4����;�C֐��Il�j�A����s�[���|�~5W=�%��<R��-z4B�j2�J��'&X��4Z��*�ڑ�ު�-j�'P����p��%?����`�z<훆�KW����\v#}@5����3�.DV�9���z�k~P���H�ғ�����Ð:�~4���{|uQ�r�"�`V�8Xs|	'f ��z�����J�Ep�$!jԞB(·��^��	8e���p�3˅P���H�����-��r\(�5�<z�3 Á�e+����L~�Ed���V)�,.e�.�%��gchul`A.��(E���C(�
sX��ŴO�Ɉ�[O� O��=���>}�ª8�+#1˔���T�:%�Wgpn[����r���k�Qr\r��ø�N�/OyH��zb�b��o�or�>/�rL S����ٴI��s�}��=&�J��3j��]�@�G�v�x��2�0w�����8Y�͑��4���Jj�@�|�(�b,|�b�*�������Wȁ ���(�o�06��dҵE,^�g��/�}v�:�EΫ3��I���CD;�,�xw������)��*`.��Q2���#�Z���Ŭ�q&�2�f��w�\C6zEc�*82c�袭Q͙h�^5�?<��\ku�>�/��l:7mi��*��%'\�1�HTyN=������O/��S�p��z�b9?E:>r��YM��뙵�X��P�)W�t�S#_l� �����K�^���#��I�*N&���� @�`�\�Ԧ���c��s�Ӻ\�\J��F���c-w��e7~n�J.�j#���>=�ǯF��?��L�j��9�t�����&A����, �
A�跄�m��dD�~J7����M�cdX��F�׍���LQm����:�6nP�� �X8�9��w��|O�~K�1h��+�w�~�� ��[�4�T�A^��ޠ��}��K��$M��ݏPյ���fm;.�AZsP���-pS@��ml���.���_�?��;Ҙu5�6C~��F�W/�;N1�Ҏ4N�*��m���X@���5,qq誺9G�࠱A�1��1|�ܩ���)-�����*�:3z&��������# X�.���`�}�ƻb�T�D�1�����>w���b�ңf����]7�
5�"r�������T�HP�jW�������i�T �sCǆ�6��u���9������)��EJ��������ǆ7���Kx��\%��f�p���,Ĺ�9(�!]/�b����G��ʛ��^�%])���D�hFC��@Bߙ罳�ޜQ���#�QCD﵁��A�n�w��"rvݫ��U-�G
?�"\�d��	C%١Xz^4�ѷ�����.k�H��v <w��v��Ψ����'�T�gL�DHe��l�Sr(���K ��D�w,��3@��.�*fHm��^ُ84p|�)ꓰ«V��8!��K�Ma�6�c��Q ����D��MJ&�`2��2��~ y�O� ���F&1�����@��؛�f�V�+z-�o�1�G��O�����f!�s����� .GKa�	E�w�]E�0�9`�� �t�K�fD��v^K����a
�?�uɩ�-�J��C�֫2.��0x��8�H�Kʢ��e�Y��@J�v�e7���V�W��ܙ����bqvԟzm���>�:����%1��O6?�$��qbcS� ��e�q���$H�-��
V� �JS1��s
�%BK�D��$�������-�Uf�rs�����I=d���Bn�������rd(�ъ}�uQ����+IQ
5F*[��� �B�ي+�Oe��N��v��c&L�k[����l��i	� ���<-�ʵ(����I�7�T:��'�Nu�y*=�7>ҟ �OY'ڀr �aڊ��F���1�C�o��Qϳ�d�M����E��kp��Z�	P�����e��b��
5��hΜ�hXt�w�]�4��s��=/�C�*]8��U��W���wi��I�mMWA���8;|p
CΨ.��sd��}��b�>>���8��׏��[;:Ht@�Zd�����l��#�^���ω�d"�Α��A��a���@�>�"I�$�\W5��k���� �۩f�&ϩ��`:�3:�/��D�YC����H?E!@py=�ʹ�� ���q�*m�����0��t�\�y��YP�P5ǰ�^��m����C����y�.��R�ׯ�h��m(�cx�k�k~9���z�`H
*�H�N����� `N�f5L��
�eyp��QiM�z#�,"���;��D�$zI8d~j?Ӛ���E�Y����ŉ$�:Ǖ�S�t1yt�c�!��_��,ĳ%`t��&~cD�Q6C"4&�
�3��p	� _�Bu�:4��s׵�*[y=�?��\�
7�.��4�Tָ�*)��f�m�&W��o��8.�����(�	!� �E4ڔ�ϸ,�Fh�>�ς�1�ĪX�|��- }��g��$��n.n�o�3�`,b"��Qw;�jK'�Kǖ�i�k���A�A�Y��ڰ4E���yP�� o�E��W6��a|���t�`�ֽÐ�楊cZ{>�i8霜������ڋ�;����������obf�K����u���D�Y+�[/ݗi�+ϩ��t�𖲗'(���Z� ;�yTz�Nl������e&R�1!��Wު�}���_�`Ϝt� ��? �쓜~��Am'�9��5�<Zq�6�I�m�d���<uڲ�l�_��kH~����xn�1bxzO�6�k �]j@��g�����L���qFnZt{����<���R��l=��N2��U}��n`���Ź�z��l��0�T {�r��=Exܩ�"�m�eV#���$l)X�� �������b��]%H�I!й&�B���u� �M�xWh0), �E&�3�rS�:�d� �;�� :Np�-��7���#g���.���2�{�ހӑ~��#v��ͽY!C���DO��R��W�*_x�o#�e�L=E�\c�˯DCRb����Bxue�ȧX�C��Q���*�OE�S��hx D�\�������䪜K�J�B/.6������b
�2WT�i�����x���˟��C]���0%��>*6�{��Ώ�x��M�7fh��џ�e�yW�R�ڹW�-&� ���m���ߙ��щ�W��r��B9�f���.ʳ8*i,�3Ё[�6�����!�Ӈ���Dj(��U�y��˞��J��:ĝ����(��{���,g��]m||�����E�����P���E��gWyb��~�H�����^���Q��cf�W�Tё=ng�������L�^o���*��r���V{2�q:)3S�M髉�m� W�_��Ѽ�Gv>�`!�źA�b�K��j��+xN���������doI�@ix����z�ST7��˶p�<뀍6?��6o0�17�9u���c讫�R��!lV*K	B����KF�kgM�,}�|�]�. �L��׼Q�5����5�������ֹ�vl�HL��3\���O,��7 8����>	2�(�g�p!5X+d�B�N�֐;OIN�m��5^��,D����!C�����T�cC��C"���4��R����<>�D+?1WVe�i�R��)�����+��l�	�44��(�$�2l���h>�Q�0l���M�A�>��J�+�VQin"�ӳ/���0@��{�����`�b"%�������ޛrI�O�+��@��-�K�)	����R�]�'90�aun��m�a�턬���Z�>�o��U%���fl\VA�����+L��4���	Ny��[~҂u_	����|>�T�f�軮��j0L�B�
�o��rO�y�f��2Sz,�1�$t2�vs#)�5���~9�������7�1�n�r��-���a%�-��N��v�|�ҖCw����[�����q	��y�h�8�=_5�/����ƾk�g�6��û���;o��(,�`}��M]6�������X&��M܅@��0�髰�R���D�����وnaW�����)����H���)����d��|�v�U�dOq�Ks5���R+֗��PΡ��,�;�2y�2�HM6PJ�oj�/CE6ِ��=�]�R'�L�e;_~���W{Yᙍ)�P�1؎H�[5��п�V�jǸg%S���(���(N�+�i[wD���E�7ᶤ� ^O��$P3���7����L#)Q���5��왓B��;o�U�o
 @�%/�!e�թ�\hQU�ژ�lB�EI�7���mc�/���,��o�`��Si�P6����K��<3����x7W�z:���,�Qni���:f#�cp�"b-Hs�L;�5�>ƞ�˺;��_������.���)Z�y�ڮ߆HW̱�+����?=x�mr�?��tx.{��
3�#�I�f]k���1,=����j����*ڔæ<�~��řwq�񑩥���{�/�X5�W�=�s�Ya����ۈ�m�.+a�X-�ξ�`�s�P�9���9��N;���	k�A����B����άy�$�x�聿�\�ۨ񤤫�t���,L��!�D\�ɳ_j�u:3�4:H4.���^i7�����^	xv��y��W;���j�o�Bԉ/��r{���k�I���'|J���'���w��Q��d��]5aQ7���>@��+����~���g����O\k����Ujv����OH�az)s�y�:�&���5e���6��\he��ֻ�a8�c,����c��`N\���A�j��qD�f�W%�ِ�Y�^�����(1~�p�|:F���L�h[-H>�͗�iÂ�f>��Y��S���E�ڷOԭ�4U�]S���o�˝2
jk��9j?�����	���)$X�L
_?�_5�9���E����U�BCŷ�^���L�U�9-J�@QL�r&$;�u�w�.���M6-�p��ٹ�.#�%||LG�=xl�VԦ�d�+���E&��p��|��}����/�F۴0�d8���kS�%0�������(rv�t�AW�R�br���|c�T��� �8�3v�Oݥ�C���Տ�� �/��1B`��r�Ee@7z��޳��D�0�v<R��0���*>��QE���B��j���P^xSW���U���;����d��.QG�|�v������*q�9� �G�cAW�7�ZQֳø�r\�}���Æ��q�ֳ�N������V�&׹t��+g�z8V�RH-}D��C�-��ث]���)Щ�)Qy㘆�h�ҝ~�3� `��u�?�G��u0A)�]UX�Us:�������<��
��X+����9����@�͋��}-Dp�o���z�K�3E]�\	�T�H#�3v��/jk��^Zf{�}¢� �H��q�~�2��&���)�����E��F��@"K5ë3t=r�r6��x��n ���QX�8��nŢħZr  �d�*\A�۬樯����Hb��l�����K�IQ��~ֱ�߈]���%�)�.�[���������*&�-|�l}X��_!N�ķ7�bK�,�I����akH��
� 6Lv��x!�;������t�&��Iݓ�g8�k����K����d���K��5�I�l�<~��S��
��Ǥ+j����K��oMR���	I�k��<���r-��/M@��/'a��"�}> ��5��[�⇺s��/�jD��&���Y{E�u���\�����#�}�����PF?�o���r�6B�
��܉;c�NG�!2�9�3O׉[�3�цD�����#�����(a���k�W|_���i�1�(i��Ťs�ڜru=t�GCv���A	���AV[�3�߃�Q]u�L ���K8��7��5IG?�5&Ҭ/t�nW$���/۩|Kߍm�+c��a,t��p�<�wz�o�� 5"���W������F����⯘�����@{���+vfa�Q\8l�?�ŕ)R�c���p�B� <�-�`�tE��|���C:�/�亟��¼Cm�'�Iw�J1ݪ��dGs� ��!��U"e�;Ms��r����c�f\B�ZT�j�n�E&��D�oȩ�/��3�O�g�*a+��b@�>U�dJ!��8{.���ؖR쨷�,˥���uӘ�s[�+e����3���Ac?"`���Y�����o�ci���";m�G����s�]�$[�ox�p3Y���`�f�?�TTm��j�DtJ���$h�j6��_�����ۅ
�a�)�)=�b��Ϩ\�V%*� d�w�$����ۋ�}��.�L�+3�蔐˂����K����3z��=�4��t�qk0�A�����Lz�S?� _���F$��+v�q�����F��ori[%�	(9Q�=xce�siY.n�jI�� H[���>>�.��%��糬���b�pX�Oi[��j.��I�_�ATb��JY�����l��a�9R��{�K��2oXo��������]��e��) |�0\�W�O�I����U�����"I�"Dl�X:�b&�Zq��9�p7t�L�)p�l �"Ҡ��n��~�P*E3C����+I�U������i�dV�*8q�ɕ���Ê��␔:�6��q�;��J��]m�o���S��Bx>�N�ܛ�[��:i��rF`m3��L���Ș�)9�Q5@'��=`����'q��]�߀�ayh~�e��eײ?�˥P�����,0��X�k���X��3��Ѱ�������>*��d�}Z���x'1���n��W֏.WǛ�?oDh����������N�9�a�E�!8�6�bSꙟ,&6˔�y��3c���{�E��|&ve^u���	��Re���k�C]9c���}&ʆ��N��l|��p��PP���c).��+�ٿ��)��U\�>t7ea��*��lZ��丨_��).�jh���U��׳V]�N.��
-,	�[��1:xhD8V&�Oj�+b�\�-�>�=�#HFM�O0"��HI8P� �o��Σ��b�6�8����+��h��<�ƕ�RŌ��d�f�b���a
9��D}�Yj���	�9�5��F'.���G�U�,�)G+�����J�r����ė'Y�>����4��T,&PJ�ZJ��jI�jT��z�f�����s��Y��6B�2��{���U���y4O�ĺ�5�3�}�^?m�'(##�!.��kZ� ���_� �+�z"ى&Z�Ĥ�I0ok�?�������j��>Dȟ}ΰ�x,ɂ���� ����y�����^��,����^��M��np��u~�!nV0��=�A��2��)��	�<�3T�����)���x�+-��
�����2r��ȾѝU���D��W��:�U*�����麝}r�U ���k�����O*�D�&m�~½iU�t�U�b�ń�{|�sA.��d�f�ظ��I�7��x�
���K��\�H�80�ZM3��=�^m.��#��V���4�(���D��b���*\(���'��������l��bű���)�''�A(}jW"m����h%��ua��1�azA�q��l���B[���6U�>����t00y=�.(p���^���S��L)+��űz�۶��'��ت!Д��1�2�w�%�u'9]���;>6Ll��I�ۍ]���J�Ot��AAA ���;���kR�q�fo?��y�����1Ȓ�lM=�{��A(�W�z;�d�^�l��͌W�#(���n��r4��
�$��OHy����iH����ǟ�fB�WsV�Q��������EW0�/b�"+�g$*�� �r��|�~}�}C��C_��bo��&/r����+�������{͒=q]m�~�o�:�������0��P�t�I�i'�����A$��D`���1Ae���X���U��J�
�G$l�� ���S:Ӯs4�����ofL�-c�ec����h�&M�7~yBU���ߘH~�c�U��}��r��nq��^,$���� q���
�PdxP��7cCf�=�`���X���
"b�N��-3���X�}�bXggہZ�ۻ�7>ذ�b�)e��_eR[X����
�Ų��tꣽ����2����T-�K��a�켖v@��ζ����ϻ��N$��W�&�`���F�l$���:G:y"ߏ� A�	a*c�IHB��J�ACl��Z5L���pE1����ü�|f��8�4�?H
>4����[-�9,si��AK�칭�0����
�k�s-����0�p)�p5�5&w�!J7������3Y9O4����5��������3���
����(!'y�������Q��tZp�����6����u�^�� �`��%#�p�����9�+*�61�J|0�l���k��(������P��+571��v\وa/��ˍt�<��K�W%�4���d���ي��!>mb���`:����vnᩅ�'��~2���_�8��nW�;��?Œ1y�5��<��on���.�˪�!F� �	�����o6-����2D4�x<<0�Y�����Fɑ��X����=��0mfH�X�Unx�ɷ�X[��M.v���x����_�=�W-��F�!W)�Lc+f��dp�0�Vc�K#�rTD�:�R�tA>���W�mJ�c�����Fq�s�_n#��[\Y������/�w(��~M���SPT��sN}g�/qo4p�Ɂ���I	 C�tp�����:8tu��0p�gV[� Ao��XU�MA=�
9:�� �4�J"�Y��f'^�"���A�=v��o{i��a*�Ӻ���r�ާ��gv��X0���q��ᾝ�H\(=��+��>�����L����2c?��T̚��mj�@��:�%2("?s~��݂������y_1-����$+���.��_+��,�ûȩ����ۍ��=YG�U�:	�["%"
�C-����^�(7�E
�~<	lݾ��wD�<�Fv�(4ֿ^�5�G�n.}����#�)�Ň����:7�\��l�e}���P��kE���rX�������Pȝ��&��ۄ+/�󤁖64(6��[���P)�}�&1Ӹv$�{�
N���t��<I3̜����fOw��A5V2Ty�����^�֟�wF�������׽�v(����G�#�����P�k��c�ɟ��(���L��7�w!aԱ�_��!N�ꏸ����c�RH�{����zE,�����{� yZ86�'����5�
�?�[����J~+�}!�s?��WCr<��ه,��fkY��CС˕3*qBR^[���N�'=gU4W�Bg*��ˋѡh����SL���D���]_Z�fqY�~��NE��μƯ:%�qj0�|����4їPQ�	G��\�6.:+�n�)O�@�ٜ8���M����� ��g����P�_EY������ �Ő��ݥ4��������n�������8�嚊/ϴ�n�B�-<�ql?�u����(��t9������<��A�aV�.�iXb��=x4h�N4Ȕ��=�J_���皰�^8%��I�P.��:9<��TF�I��m�x��c\K0��rJ����\N�C���Y����RqV��5T�j���e�ɼ�L�Н�lg�< ���1�nv���Ļ�R���!Oz�3�3�jn�V��+�w��J�F�-�=�[�$�ްw!k���~8Ѭ�w��/,���{L^	^��t=�H��`����* 朷M":G69�K2�
j��U���@��e)��1ޥc��ّc	�v�<�x��+���D�'KԈu�`'�<�k��a�Wf�}����s���&��9��ZQH�&��o�%�$��@�V�-|>WB'8��:�K�sO�@$�Ԧ�:xK�S3��VƔӓ�����d���Ȏm\�_��%hg�OjU�Е�}J�`GhF*b���]d/��8�IdGH�a!���>�Kׁ;��n�آ�#�4A� �T�:�]S��zHlX���)gϡ.������]=�>l<f�~�6����_rd��x�*��T�/���U�~;��;��p��I�p2���ebeT3S��r��Y$FAC�DQ�"���6q�P�e�����w��e��we�I1'�����񯅢h֊s�QԐ��B4�m���e������
-�|�R�Ěܳr���%3�%�^bS�H�~(c$)a�y���pO���'C��2���p�cC�L73��I!Z,�����U�y�M8��`�ēo�:��q��Vd�1�#��w�pD�%򬎈�0����x��5s�+yi2���дE���η0V������P��o���R"��Q��V�B�ޙ�&�H=K�Eix����2T�wʱ��H����ȹ�D[�����b�F�x9�p�I��yT� �"?��I�Z�@�2��I�8�{`��t�;6<���s�|��0]��)@��� H9�z����74f�7��捅B���x����u#�ڃ����>_w�r����`��&둝��8��� Hh�B5���|����Dt!�,��D��0��>�"�4�n��������t�X����M6���-�|J�ݴ\�������T�6`_M�)p���̴���*�,�I��	�<�]� �dD�w|��t�9��$�͡�)R��)��I�O��J��kG{�g�_��ݼ��4}��S\�<	�-�ee"�wPJ���3 I�B�L<J�7�Q�����؄�=����)롶�6�������S��P*
E�ґ߄�}n̞�rd��g�����%�j�����I+��0:]d�i0x�XS#'��p�������Yh󾅪����|�U/�y��`��Ӳ�T���*��`t�J���t���
JL��	@�<!;�o��}"T�,a���h�ݻ�.�� �B�u��C=���Q�Ǒ�8��U�>���f�r2�A�U�u��sI�q��{,QG�C�Rf�-ivX'N�Й �G��M��a��R������������0Gr�W!��5���,D�( �ws��A�� ���:�1��Z%ଯ�������rӑa ��9��8��W���J����/-�F���_�3��ꊵzF�v.�k$��/$6�]���1c%f|��K���w�ն�����jL'�_*�=�	yG(A����a��Sd�=\2���Fo�"���VK�ә�F_�{�t���@NI�w+ၶ���Q�5P�@>�کZҘSۥmt���v_3����o�a��CB��ضs.�*�t⎓���M�I��3w�� `.&��=����VrR�[x*B��zP�߷`l�E2ծ}�qh@�����{��@�)�<�;W�]?ϑ�/2͒��'+(?�B@U�+�����t���#�&\J5�`�Flg���d�r����oB^Jk��Ɂ�Z/�h~�z���6������re7����z���7j����I�8���0���30�I6À�q�y��J�L���9!ѧ,��8�9e��E�$�u��_�?'b�L�\��n<����?��l���9�7Z�{��V�u@M�3樯>9J�qA<\!*�ti�k+�uk/�ʍ��Y��d~a;��Dԅ�9�� ȷ�b����'�H�Ĥ�N�5��Rژg�>�n��T;�A&�HX���\%��FMM���n䗗21e�M�jH�pHl���5dI`{��.�>�%��d��NJ�j�C"t<;p�6AR��O���	��bo�	���B��47��;���<2�������(��Ԇ��`��ƌ��z1�[߇�nUtT�D�AV$��:� �p�p�xM��Y��,F1���Kg9Q%�k �A�b�Y�z��z���z���;����*�_�|��l��T�7~QF�"��3�����Ć�?�m`��*�7�ɳX�^r�F�sPn��Ԇ��T9�3$)�1l��3��|qJ�V+�}��K{��QK���v"����I2�[�.^�k\�ݹ�*I&�I�j�9��R�=�rHZ�Ka �ڈ��J���^{���LR�FE�9����R;dcM(H>Y�]�)V�E,�����w!w�+.�N��&��./K,�]!�X���~��&��m&���4K-�:��T�Ѕ�^}h��l�Mu\���&+�ټWIc��.Wn������vl�� I�����\����mc�8��l����P���5�e�C�����sj�<:�^�)�k�סY��'��{r ���I���_ݡ��9J,�l� |Ե�ACr��5�����%'L n�1U�w�:��'O�[{'��X�;���Ӻ���1
���¯���Z5kă��qLI���>���i��t�$�����g.��k)�k�L����`�.�����w=��Q8<Ұ[j���X5�V�+H����({Y�}N�E�H�^ᐚ#�?����Y�<L�x0ʷZV���:��FQ��?�e��k�f:y�-�%>lҪ�sh�
A:e��2.j���d��8�L"Wy��V68��ݝ&�GG�A��+Md��Z��Ȅ����)��.�3�@�S/$�
��ϔW�&���C����
e���ٍ$�����s�G��xg��	��6�C�	9Zu r��ï>v-]8)%J\g�ͺ��c�~�4
�˚L���;�ە�;�Ѱ܌���[��M��^��ﴂA�ES��e����0+Z>)�t���%� ��:h�^���a+�/�Z���h�M{ױg�;f��;�]�ۖ�I�L� �\��d�t�-�����;j0%���bm#�.r����h��h�O�d��P�=y۸3�[�3u�.���8�("�9�jH��]�4��%����s �HH��㰼`�D�*5b�-QQ��읙�U�邺4�U4��鍽w��E7P�؍���������%�M6r�B��T�:���>�R��uT��LE��Q��'�
��?'��Z�C7��t��9_����p�}�z�|��H,�V�^�����P���	��������!}��K�֣���W�J]���e 8v�ɼBQ`c8��Z�Ö�80���]��g�BF/��-��A��-��C4��w��L�}��חS:	�c��F>c]gPO�|<��U9���!3��}���Y$C^*��j"9�K���DA��J��s����W��sZ�C���C�����+8L�Gx���E��'	�n��q���O�z��҅ďU���E�A���I��i�\��sK,�x�F`g	F�W����^�*�^�ڢ�Q�g��f�9���&��J�;��D�x��Ey-�F���Drڳ ��6u M�;uTC$Y�%�-F�0�M�&�{^`�aYX�z���d;,�K�;\f��e��z��H�%l�B@���>�<���ˋ:ց}
PK�<�YL�㭓j�T$neG�Y�Bm�		@�i �#v���V�Y�3J9_bzZ+g�[�(�%��n����)�*3�п�����&-��fE'��y���=X�/^�I�?Uz��hYm�9&L�Sq��63�ғѨ���K{�0���_�*9�慉��
:2ZH-�ͺ B:�pm%3AP:Y��N�/�^-�ٵ��T��T�|�C{�`�\���_함��r�\а@Y�ќ�#J&�f�ק��9g��F�n������r�^f�'��.���i4��l4>W��b��=�٬bn��Mt����n4�^m|(1���L�+�i���#̏s��畈@�R�U��v��;�-�K{فw��#�RK�a���_�$��"������y��4��.���]�\�"�{��؂�q-b����y��%~6�9�����!	��Z��4�f�Q��q���Ϳ�^R����ص�q�V|�-�4c�[s�C��'��d�@Eą�s���E�J���y�I0�%�G��,޺������x�����.`U�m�-��̑*�szV�e��DU%r0��I�r^d!��<JͿ�M�yW8���?�A~+
���Q��Tpelϫ�Bq�l�>P�k����\����w�ۿ6�P,���g3���?t�\�9 ׀��Um[4���ռ�F�K5�=
�Ny��y�zG�Ԓn�:�KG�o9�e��A�b�0&z��������f��ڳ�Y���`G��>���λ�Kr�,�`x#���!��|=� p�ȣ�b;�1���n�[y[��W���e����<��(���?w_�=����@Z]���=h����x�_�~�z��Ї#^�c��>D��,y	`�woi��F^K��j��s:���F.�F�6�sd�����y)su�MMS#� lM�c��"O7�y;D��L�	�#C���4�7&PW����#��.n�]���:�{YEB��3�z����a�������דw��������������(:KÑj���~6K���Z1�����W�qf�V�4kj��QC��>�9%��0+��M��zdؿ��n���T� �vOg�Ů$6+�������;lN�g? �oDV��B�Pf�n�PU�����x~�4.� %#��#�D&�a;��hZ%
�f�����iȁ/O��������R�1��+��h�p�8L
(s�A��F��]�	��1&{[�PW��DmlpL��{^H��( ����X����z��j�"��㯉�t{���cJP��,��_z�E���-8�ˋj�`נ������nn38�AGU��ъ���\�&�K�"x�P�%4F�s��	'_X�&��y��������e�%a���,_�&�#��x?-8DhX3�?r�.�]�t�UF~�1fF����rW&^�Р#|mZ	�sm0�D���\���"~�T��?��J��P�LX� ֆ�`UX&������P���"�������>]ߛ ���s2�*|�m���l��ƾ��ǟ>�j��G�tW-�IM����3��Ș�Or i-���b���%���#�� 6bvu�+ƛ�wI��h��ũ �ԍB9<�>O���h̡9�Y�Ȋpʷ�\`���e}�K����Q���T�^�5��x��	C������x�����#�h*=�&$���DO��A��Vr���1�/�=�1y��=ijZ��9M�'^Uʶj�l���v��D�	���"ҳU�x�Q͙]g|Y�wn�E:co��t,�
����fS�	�Qq�n�v7�+GE�#tv�K�F��R+ff��d:`�\^.��T����'����h.> ��v�Ӈ�H��ЙG�|��|.@�\A+�J��g"�:��~C�$�ėU'��A�Dl�����=���h��I��[�m8r��Tk佀�V�_�]'�����}0��t���>+\G���ެ?*cԵ9:d���m �P�:�'Js6�3)���l�
�dюό�0oP�v_�>'��IzM�>��!O_�ԕ��j��N�;��`n����wI���Ry%?�g8�|����xlj}�#q����; 7E�a�ؠ��]P���RO�ﷹUOX�rpM^��*�TX��j4��:Vw��Xs���H ���]_5wC��	�H��:�֗��-O����X�4i����ǔR]/!�EnFݘ�YtqK��ؠ��8-gUAQ.���πu�^6�K��'���Q�'�L���-�yUC��	�j��acnn��I�j(��O�+��uH������Wg��ʺ���H��<�B���k��.TP��Ŕ��EV�I�R�qA�C�<�3Z8�_y�*�U5�}�3!�a�&���g�(X��S������Z��>��d�E~G��f!��^�
Ϲ}C4p��VD.j���	 ��#�|9�J��ja5�3��� ~j*";�X4K��i�e׼�'@Ye��+f��%U7�R�:G\�q� JM�&n���Ӳ�w�E�;Nٌ�do�?,����^���L9|K6A�3�&�늤�0x�Ľ7@t�3�0�3�pa�����$j~LI��A�C�~��Z���q�R���;���=ґ�ÞOE�~Sa2-�:h��M|�0#�/��A�{ۅ��z�$�(�؞��D/�*���c�����ˣv<ňNT�\7���β��ι��O�|�#��<SS5&����ʚX����Z)�b=���9'6��3��&�R��MQsp�t��\\���u����Yrn���b@k)�x$�Ĝ�w��&���&�ܶ�Ֆ��
^~�yze��L��-���r+��À��}-&n2S}9Za%>��S��;|`H�iW7��VU���y��a�������ȷG����C��FS~�BՆ�g��m�v���3����aY�8aSM��t+�ǚ�{5�p?�������OZj���V�n.[�� ���_8��(O˓O�g�D��un�>�8Y����ioQ�	�*G�U�+`(�@\���m�!�$��X�d�
\�B�W��Ew�JH����1�7�.M�b�.+��kq	������� J ����L�J����=��:,W�/H�\r����1����h>�{دs��p��DoY�S0O�R�H-���or���Bg0�B'��KT��?	1�~m�0�����O�)}�s1хɗ���V�=)��W~�1{��VH.�B�7]i(��9x-���&�[si��d�upW}���������T����	LQ-��gu��5�g9xk��TČ�Dl�n�XRJ��+3�n��ap��4�� =�@>qe�s�<\@��[.oǻ��wfj5?��I���l ��$�	LU�.&��Xݠ�$}T6��*ؔ{+�/jTZ�[�3�^�jI���*��^`s��o�xǒ��`QBw����⥮�
�Vvژ�)��?�0���*�?�{���N��� ���S=�c�ϺP 8�6un]�OFi�N��ܮ�"�L�G���Y)a�1V�
E��l�=}����/�c���;s� ���U����/�
�1�84;�}� ���Υd��10�{���z~m���	����>n#�-�:�?n.AXݺ��u���o��N��C��w|LZ���~5W[�[��FV��!^9;S�F�0Q��DO��/G�-��Ф��	.W*iH��B�QW죷��bOI����3t򩴖��흭�[Ϟ[�"ȝ $�����x�%Z�9�hp�9����Tw�[z���ؘ���;]J����:����W�w�^h�����i��Ȟ��/B�@ʕ%�%?�Њ��9U�KQd�/��	��^ޓR<z�O�yϗ�~�d~��Y��*ɉ�=�N`OS����4X[�ݻ�օ{�1��w��fA�52ȗ��nz�\1>�dEgLUEf����pÈ�k�
� ��B@�ܻ?��2;�y���9]���yJ�q�|%V�?�׹\�r�3��ñ��֥�=��`�𻽰���\[B�+��-�h���	Ga_k%'�8��X��>2�7��@����|���~,��շV�'�˻
a�e��j��6)R����[d�Kp[>�c֌Ʒ����ڲ �ޯ
{����y���`�V
�b��Q�Y�r�C�*iKm{;�sԜ��x�5�̴�!�������F���KjKp7��%�y��w�����\����֖\(��><�H��g���v��Q��p�6X<�fk�?�\B ������֪�I��I���
,�&�5v`��Eo�L�DL�,���z]c
jP\�5qPj�:mr=
K^f���,���f�<u��&|,* G�X�O(�4��Y�W?mLf�Ϯv���{�x7�吉)<�x5�a&�g\��h�	8��5l�/S�%�C��ta90�����'��*�5���{�v���_w���,Ř1�6�D�i���B��R�B(r]c��Psag��=}�F�bUPa�B� d.U���+b��GN�)� ����`�3�&~^N ��L�&D��PI�E��>���P����:��K�$Y���R>�?��'��-�T�p/�@�f)���i��@:)�3���ٮy"U��j1��,��+�9�x5���Xv�7���w߿Ԭ|wǆ[�rl���� #���P:&��a��1w���<������}a��(*�9L�~�F���2��@℄E�W�˪�@��n׳@���{]�n�{
��5���w)C�ƘvN���m�M�Y�O�W������`�ë`��l��3�,�m(E.������vī���@j���˸��d�>�ù�!!:(P`�@u�I;�}����9�U�y+E�����4�(��\
g����;�LV�Z@k03��^J�M޹׎��h�����5~?6�_�
��	.�K5�ZՀdV}1ĬoTO��ul��-�`�H��ھ4�|O�����`��LGS�1�?�!�B��L�|�w�ƇfQ�m\X�5����J���d�9a;p�p��'ͷG���DTf�+"h�ޮӱ�
!��K��%V���@$d����B�.?���Lc��U_^6f�܃E��{ώ6��=�ML�U\#�m&H'a��E�^@)��s�sZч�g�"�"%0&�9u��/N΂����%k>S|Yc��*��7Z�~�U�I�uW�5"4O+���VGŵ@)lmڙ��W��é�Z��A}�ᛞ��$j������ԒŢ��Ͳ�Qc�f�����@n�]D��#�eL����tNp�!w%��h� ��<�V٘`�(��~y�k�$HT�%D�d��Wc8�`K��j�:�o�|��|�f�1�� А�/����k��p|���5Ph�ѽ� |a�{: (gW�_Ygu��ʤ�GL���0]E�l!�T���F�&y�	/Ѵ�+�+֮�`Q�\n,V�%���#�Y=� �-�	�N�p<4Ni��s�Xf>* "�sk�(�V�R�_Kp�RG f�d¨�Ϛ~�Ls��@��m��ۏخP��7ʏ�B�����@B�p��fu�$D����9Hx|�b2[a��O������hvA�8f�3�[�tS�EV��lI�o�.�=�~�E�r���cj���'��0�+�[tt����ɒ��� z �����s��]�iĄO�U({gY�֕��>7�'K3�..�h�j�sX���.�/7;p.u�+� ��ʆg�\�b�(�x�1 :5���;:�$��57wt��/r����]s�LC�z4���l�!ߴ����Ho���J��pzRA�V d�����tH�Kp�5!���C���O�/�[Y5�=��[k���rQ�L`�k�J����T+kn��UR?���/.8�D�6��IA72h�2��l�C<a�\���%63�}q/�
�M��VK���9���i��J�V��'\mi����fU(v1��-KS>��Jg����Up|� �����|=Ikˣ4N���<[�3�좇�ȧ�:��&�1��}�aGb�J��U��E��s���6��Kl5#ֺ�S-O�����bZ6�އ
�� �F h7a��Ud5'�E)d[B�ft���	lH��
z��N�Y:�c�I��$��zOU4aoѭ��	�/tԅ)��Q���wb礛Q�֭A/I�J��n�i;�s{�\|���Ҽ��� ��g{ټ��R���\QY}ɠ��Z.R�
��������;��xfn�+��W����A���i_XMLG��2�D��F��PiB,?+��ݙ��G��*��O���G?��D �	�ٿ��^�Ve��i��?�)�D�HɌ��e�ʜ���43��e�f@Y{����PJ�W`*R4k�lo����#L��ԃfU#cە:\��̩h6Ż�!~�f��YJ
rfzq�D��h�w��_�⡴ށ�U2�����4`��W|7_���ú*�IbA�)o2p�`(͚��qx������/�`���*�ρ�>*�����9� ��+�cTzV��jsF�J��{�بqh�C;��M�7�0	D�sv����R��%W�ث�^a��Ё��>N��_�����M,/U�Q)l��<�0)$m�f��Q*΢8	>q.b��Ovɂ���a{�.�j��Ԥ�o��fN���qU�k(A�%+����"�cY#��6�~�Bx�!�������j�����4�;��C�H~���+���j�6�H�җ�
����U+#M��3\�P�[��I=�66'����J�Wl�S���mC�����ٞJ
؁���pdh�!�F�P:4b��Fy ���trO�V(��I(U%�M��Yd�Jڭ��+���/ؔ/���>�Ghf�y��Ԕ��CP��ư�g��]�iU/t5������@���} �[�V�:����,|:פ�1���vGG)�M��
-����RmAs*h���'H��B3O�\>u��'���0�^�:�&���@�K}F}��_\�(���>|��m��_⹝����K߷�o�EAڐ�N] �y� P}j���Jq�E	�mV4݄z=���@C�7�
�mϠ�cԺ���+ ��%�q;M��>�O��:�<�Ӹڙ�����Bh�ѩ�qW^|�6s��@�R�-l1vӯ$|�.ʒ��V�;0����xa~%�T,�g����@�oiƨ�Gvc�5��� �E$�����#�񝯌����xGq�5��{�rY� y<&1��+�����NO��)��ʅ$���s�7�ݮ6%H��zO�ح)�T��u�S1X��F�|��@�0"7���T`���>���ьs�I��NgJ7G�ȐWrݯu_ӟE?wM����6���×5y��ő
�� �C;�,�i:��,�џ]ٌ7����G��x��X&�ܘz��]� �����
|�o�R-���W_X
�9f��J��3��Mn[틒��!��5(O��<�ʷ�=i��B}�z^8�c�H��R��B��(7i��}�0�yʮK/Y+�����ŰT��i:��t:��\wӶmyq�*��	��9��Nt/����lW�=Vrd3q����6=L�/�u�}��h��1N� 2��D��F�'��6��h��$��J�xȂ��C�0�B��qR3	�ȗ������7��7�Ė/ߐ���s�$i����=x��J�A�NY�ര��'"�3�W���rC�_{,��%)�a�W�q@eaDtC�<z0O���2����^��ď�K~�N�*ĹXRF}1�z��0��J�)j#;�yt�w݇����z�v��V��j�����:��BK��;�׌�09��Y���lg���M�E�}�Ԃ��^S��Y*�4'���ey�!u�89��6#m��x�|�QsMX���m�r�9�Hδ,�s��Vܥ���S��SM��8��2���i5�����]�+n���y�6h�A�4e?ڞ#��M����4�Y�QX�0���Vj����&*�-�Q��8�V�r�>��y;`Љ�%��ܟG�gx�e�����A�~�w�M;�Meo�-ɭ.��È��	�!�cĂ];���A0wP8��pk�jn���&> ��"�L�[�١����2��$)fy|�W�f4Н�[�c_��S�d%_��)w�q�O�n* � ��5��p��Q��Z���E7�ɕ!�d��G�-vo'�$��+��Od�c�q5+Ёl�Ղ�B���1�n1�"� H_J�����4^�9t�G9�yXS=�|ġJ�s)�Vp��"F�m,�9��Vv��B\�#����k\���?�>����S���	c)A��P�f���U����.l���a���|�Z��i<�\���+�����Uۓl;1�5�P�n���QN{.������-T�{�.��[
[ʢ�qd����b�w}���Bū�Z��hcHs~�:�� >�W�O^�5���R=xI;<&�P�z�%�(��Ǚl�^[��ܖs~;a����_���l'�C�W}�ON�a��@�9"x!�r\v�U�������<����,f7C�Y�G� r��0:�fi�)����붟��)�&-����R�#�Ӷ/�H(a"@1;�ěs W�?�����ޛ���5@ ��?.�@EC�NA΄��5q{#.����Y�G����-�������2s;t�
�� \��Q����Ѝm}�3e�^����yvUw��/p�7D�-�!l�T�9��͗���x�n���߅zv�<X����m���7�l��Lk�Tb�n�j��D]%��ۈg���{>��
� 
���^�#���<�"���v ځ?&=�ﭜ֏5���^�=)P��<ض~����z]�s<ˆΛ�H'�2�X�d��;����5r�SJMm)zb��р��S)D"���1'��T���T�
,̟$�ۆv�K=�R�?�)��� ��,��#M���א�ca�	����n|���C7� �"ƨ�Oϝ��RD!W��q D�{9'��Fk��3YK�oS��1����S��3|v�É%{�pI�XK���}�y 5�(��8�زh����^3���T%���n����9�m'q�����w��M���v�W��_7�%����rH��_�zQ�ev36��:;m�!��Fj���`�TM���"
��[�Ts�,	�����ajV=>7γ����I�w�׭��_87� ڴE��(;OzXi&@�������=�i�n��۵g�����s����A$ǹu�
+Bm>��u�>�O��B"{~JD�h��[mm�a��-J�PHX��@�Ɯxʍ�D/�oAR�"Q�����,�xk�9�Iΰx���L-���
䧖8�l;��濠�q{�V�O�1HS�[CkWQ/⣡
?�۵��Xb'�\��:���G�,j���b��۷����V�L��r��z�dB�>P�/��H���~҄��<�aƎ`�w��N�����aӃΚX��j�7�����j�����?�nk���~��J�(�p�!z�P|\��0C���[����M5�̄O2������!DBHt�x���4ԝφ�%)�tjX�l(����d|?�X�\��kX��`�=#�4s���>���.�9'�9��E�G1�ۧ+o�P��X�?�r�9�ٓļ��&�D�KyAP�H��5gCA���NKi�H�"a ��fY���ք�B�o��#����p������٧��P�Za��Ǡ2淾p0T�����'(l�_�r�6�O�M(�x����?b��n�^n["�'�X�`�5*(��>P�!H�3��x�^lZON�J2&�HԢ�����e@�v
S+W��� D&p]]��:�Eಯ��^�!�<����1׽\��Z�u�0N�����i��:�W�6���Y����4��s]��HM��ZCV���?��7�8a��N�?05��?��	e�#��b>�B����������F��W��@L�>�0?��ͦ�'��ϕ�<o�-���\�U��U��c�����Lo��dL���A�3Y���jʕ�����7bS��墟&9Yq�
�6�\��\B�`�jT�5�C�uzEJB�J9��ʏ�NW�E|��n�j�G.�|&����{�I�2H.���U���=Z`<jk�If�P��87�˦�m/J�ѥ����.������LkX=�9�0�5����^Or��D.:v��)Y�0��{�3���p���#�jԥ���=�8H!�ܿ�o-�YH��E��|c��|�z��:y$C�^q�N�MU2F�͚9���
Ů�BK�! ��K��`��٧>+6��K3c�aݸ�<�Q���D�	(�c�p63��/����W���o�}=�[g����e���·�q>�#(}�����*'׻|�~S{T� �í���\TZ�+X��@��?E)�f��*e<�٤Xlh!���A��Hh��?���܋���]�z�_[<�������_����̀�"�M�?[.b<�ZZ%�ebI�#���F��)Jmk�.�i�Y���3s���3|�� q�/C�;t�\�a�Å~/��(g��,yc/��,	ˬנ����0��ڣ�����E�S�A���-��5��\��T@���w�v��;�0Qk���8�M��U��-�0��������p?՞&�,�U��W����8u��TV��p�k�=v�_
L�[�[�b
S;Ҧ�2�o�P(�P�y�j�0)�t���
֌�F �,1"#���J��*rV$��GT���V�|��?�����`�,)x7���"�1�h���ԥŘ�7���W�T%�$��T�f�i���)
�P¼��"#�W�3-O�tj}.ōR}�q��5�S5h��c9x���"���� ��ء1(�3��M�E�gq@�������I�1�k�6����,ӯo�T��R����o���ݳ��U\W�d.Ah�SVﰔM9-*N�K:u;��u!+�5xZ]3Dr�D���	��e���]K�	�#�C�y�	��.,N�[v����S,ArU�*�|��軳
`�h���g���1�D=r�L���/X.���Qa�ؾ:���A�>0s%:N����_Q��
�t���ةU����`
v��Z��>_�����5���,2�y�Td��k����K�i|�T�?��D�ٹg�Dւ5$���W�z�ɺ����,�?D�>�����۝�"[����R�rDH
��.&NZ�\O�������Q:���/��R9�����Iܸ��
�g�Qoc���}�S�ߧ���p���ے�y��}db�d��m�D�oTR����3�s&H�nXŮ���DIՃ���։4�C��*p�����#�&ND�*���D���
.^���.Iu�{.�ÂΒ��խ�aL�����XV+�6�����W�}^i�-/LM}Tw;TN+�ƞB�Ϧ�ȮV�o"kzo��������_ĮDȑJ#��`L�����6_[���P�U|�s�ӖeD�J� �� Y�fA��5/����j�\"���<& ��/Hߠds���Z.�$�z_#����L8)r�@*`bi�r7�f�2�vl��J	Q2��I�%n	�]��@�ǬWغ��m�{��A���}3d��:S�?5�����'3rѺE��!��!�paW���@��ŷ��~l���s`Yf�ɾP��>�J7�Y��b��?7�)-sDH��8ɻp��V��
Ii�gv�ChI[m�z�^��$iZ���l�ܹ�b��6�ز����c��a��8?Yp[��7)�㔌r�50��E�&!D����w�+X��B�=��8Pf0[IB����������������+3e��2�1R��xБ�Au�l>�E`�S�'�P��RG�k�ۆ ����1�G�ʗ���9� f�R����28���jV���� jc<�mW:U��7>R��Ս�G,1�!:�G^
��;�8S���%Qo��56!��6j�k��H�6��u�d��ks��^��I��M��[�K#�4����i���&�#_����S�$�����辈���ޭ�5��|3E�D�"e�#��B� �W����ާ�mwڿ
i �*�c�uapZ���C���\J��v�Y�
^J�gSHk��~���?��3O�%��qk����|��p��C�\`q[�޽ru��J�{�Eʩ)���	{�حl��*q|/��h}��$\��%��L�k��\k��p0<d��a�]���P6�ؗ!���4�#eU䧸��[�c����oP�)!�3�qH�Ip��+�F�l��ųq�m���"֥!�K�zK�L���^1���V�)�?�����|��Lt�D(#��=h)Ɛ(y�Kir������vd"(8p��ح��qyŠ�ޕ���v���ň���Bn� ��� 0�>u��q�K8�U�<Kީ8O���F�ƮU���&��WݹU�>9�0��,s�4�h�`Y?���[�A)&�-J1/��@�p�w���E�X\;k�Q
�+3�W ��~˼�LD/vTN�9����_��2�{�_�&��r�#�$����k�Ńt�c����K&�v,��W;�s�z%�PJ����y�����6�l���>9{��^komB��u�S���: ���D��� �?:�)!�(�J鎎�EV�aײ��Z�¹/��/��*��BJD�I�wo�E�\�~��+ٓ�aj�V^s�|�'sڻ-�3�z����Z���ԡ@Ax7��w�'DD�y/\��xH��?X��~X�zN��6$B�o�(0*�l�vrN���� ���0�}�f����a�l+�w�㼯����,2[ᓔ�ח�)����0���(�hU&��T-/{?�V���E`�ކ'|�B��'��J=�#2���*�=3Y�����J X�	�	������� ���>&�m	� ��1إ����L��r��#��� <�.(ɿ���vǤ����!�ps:���+�����8����v4��s��,���s1�*2�����Ƕ�����NAY�2@}-a~C����Cx��������jO�����C]�Rh��y���e�#Ʒ	���>h�]�}u{L�eޏa{U�l�����9�fF�����6��O9I^V���n�ԞI�2�k��'�[��8ן4��z�Q�Q��F�/��\�?W��6��]��S���DV��#�=�
��]�OS�� ��ž(N��bP���B��� ������j���	���Dة��� 4�
��/�&�08���T`���u[>���I���]x^)s���+:�j��{ψd���YحQ�&��?���e�<N���P.BcF��ޱߖ�Z���?+�>���6��9m�C�??�q2�:)n���?kW���4�4��2�����0���mȠ�s��j-��9�Ó�����`S=�ߢ�s#I�?j���}:F���O���X3r^��y��g�R�P��N��h�1�0��96o����xk:�ؗ�L��#�8��B�������a\/J���L^�q�����}VU� �+�n�+-��������k,P��$��A�׀�KٗaDE.��=|�{02�x2���!���̻'��Po���dO��'I({71���~^r뤗�cnS<���We����{U]�}�Y�Bo�S"G=�M\��7��Y����|1$E�'��^Bn��>��Em�Z �%�XK��#+�r��dMU�k3���-���9��O+#� ��
B�R��u1���C^bM�1�B�pH^^�J�Źt�Lz3Vp��3yO�����?��F��V�6}�e�M9`�k�9�� �c�ٓ%��	�?�0͍���Xy��>36���#��g��|a�*�6;�J�ɛz�>p_ �]��4W{�@e�49Ly2.�k���~�t�*����\>�	ux�D�Y�)���3����]<��>Z��_U�=7�ǽ��F8�p�_\ft�}���Uu#�����2�^�E�P)rm��Q�~O�fR�N�% /F�=y�-g�o�2�Sm�U1}���3B�%�M��Ȯ��U�����d�QB��L�+h����jTd�h���e}ڱ`$�<9Mܐ����i�E;����R�ڀD͝՜0%�F�fG'��ebN��3B��`~��ʉ?�qDH6[��m�����:��n �����b�����z,����f{��`�@�������s�Lvh�35�5:mT?C�� �W����Oc���숻���>��+������CZ��紻s�8�����n(��6�Q��~�o�g宵4�؋;z�y�r��
���9Bڟ���
�'�ՃI�\�<��!�D��^y'�1Qɻ�W1��D+Sey�&je��َ�&-�hC���)��f5(^�X,� )}X @T_��8�`�זh�Ke�ަslM����rK
 *o�8'�s_q�2�"lv{�ψ�#{�)�<��l�q�����얽�p||�+޶jt�pI�E����l�8��S�^��56;.�M�b�v		�� ���^��3B���-������sfZ���iyȣ�b�G��{�+�g ����g/���Hr��͠]cD�(�h2��@S�ڄ�,L?��!��1�_c����u���e� ��>�9��a	���K�Y��,*��>>X�w��,!!	]� 0H�+OC'�Vc"�p1/ٌ���p��o��q�uz�ec%�z�$�÷9�.��(�߶2@m �x�X�G��A��Sm��r�^���д���/\�=J ��߳1G�\��{���mN�O�k��4|Jx?�d���ݟq�W��]��lv��J������[�kb���N����f#����cI�r�E�t�SXI��M�����L���Y�%�
 ?�Fᇮ�O��?\Z��nv�_d�J����Id�b:j�����Xqh���>0��{0��Hm�4C#���8��?X�XD�Gg�vRe���[!��̘����Ӥm��UWÓ�����=\8۝��❾�K�g�s��4�M��-�r�ɐ`^�o��N�"U��<�������F�V��iiCA����w�fU{oE �ӎe.X�:9���u�^�����7{y�!xֺ�nqS��qH��`��Lĕ/�&?�4�� �N$"o9u��_�{�EEÑ\?�1Æ�YŰG&s�nZG:g�\n*Ǫ��~���A$q� .x�o=���;����j��SI�1;z63x2�w�I8p�sz��������ĂϪ��:�]߶ 薐Ű0H~�< ���ԯ��k͍嘻���س�m�!v�M��j���.����f������0>B���:d�c��ZEVg�z�Ɵ��rD�v�EEY��a�γIgD�� )�O�d�p+����x�ԭҺ�\J�B������`�q������z�ћ�+1�*�~ҭ	�m08��J�r��}wY7��.30	CJ���&��Ϡ00�ރ��\Ȍ­� t�"i�ѧi�x�q��X�v;.��7�5���h�6�6����tf�6�{�4^ʰ�Z�h�\��!3�i�|F���@���GUA�4�R^S�Ҋ7�}����o Z�S�!���{FY#������%N������b|�eY�,�t���d;����J%ъ��u>P��Xr����d[� �^�7�׈��ƴ.h�:b�<�������O�����y��Y~,�F��qHqye~�v�i�F|}n╶_��x��nY���$������T�N1�f�� ��ɑ���6~�n��[l��7�aK���;���6y�Ⱦ3}�$��R��Q���z�d��8� �Ť�ˉ��.���ںS6��p�%��� ��{oO�jk� �2S�˫�P��8�4�����ڕ��=�j�!�]��8#�^�U:$Cc�#xA�����Wo�!�a�GG��<"Ћ���ًJ��֥(���|�2�],�I�R}�EC����P��.�;t���쓒��C*���f1x0/
��uNtJq:2���f=0:��?:s��L5��^~j��pg>Գ.��6
�,��Р�����@��%�TK����Va���և�D�@I��p+kQ�������c(��c�4Α��`��:�z�(���C�rR�������6&(LY%�sS�*Z�|?�OCI���U��l��y��%��������D�H��dR�q؍�Y���>��.\������i�Pg�A(7z�.Q!9]���fo,3��b�������
q��S����ńha�����ۥ�l�c�~'x}�B��oA۪|���ч��@φ�`l�,�E����?:�
�tw����X�r%2t�J{8����%؊��j�B		�̋ߑl��l����{34>�}��l�}�9`F�cG�k�$#�6ھ��~�U��6�Qξ�,��E<�U��1E��ob����xI�KƄ�����rдd�7D��gUO�/���Ote_"�Ov�r֮�-P��t��@�xD�:�<��f M���d����0]��T�蚀��G��9r�=9�<%A���(��Lv��M��1�&���T��/���yg�1�Q9��L�{h�+���ÿT�P�J`#]�~�YX�Q�:g�zY�k2P��f����p�~��$f�$��IY6���]Y�~[�M�-!�����<�܈�"����؋n����Z��q-��o$�j�@�wp�[����O@�p=�Q?B=����c$u20a��~|�6�|۩{ד��|�ә�d#;���͎X��;�i��Ҭ�C�(O*���4��#bV��m��DT����RV�/����s��j`�%A&d&oS/)�E�T���t�Y�Tlp�|	�j �q,<d�֮&~����:2Hف���D��q�+2�|�G������P�[���}w�s'�m3ςh"K+[m����@���̌[��t���f(p�g�Ns�����hK�EI�b9m'�0�ǥ��L����N�/Ж�%��[A�Я� �����Htq���:��k���R�L�4��l��]<���(n�yG��(v|	���tn�����-�=;���%��<�6��|_ɐ< �3=/�mΕ򗮥�L܅�7��/��;�/�q���&���r��	�wrC���BD���F��b�2B�z�K���_�������1mE�۪-��(=�"��06t͢U?�'2��˴�)��+	�g�B�Hi%r��I�8ܙ�/�O��:ٕD}Z�)�E|�P��*O����_�w�#�>�/�ڋ_f7���Lճ0��|;���*b���ۘnL�]�yV�;W��~T]�0F	3���!�] 1��5�������j����O���+�����^�8i�<�`�rG�ʹ�/3'>�\k[�`*pg	�X����OԬ!���z2Au���s���v��A+�R���Yc�FEs;��\
EAj�b~U�:�����7�a,mi�F�/nnUE���	k>p�"$$��P�U�O>6~�����e%eD���n�G�b!:#�N��6<y��4]�2�e�eqo
߯�H/�tH<�+� ���l#[�U �oa��ZKs#�j�d�B�*��s}{k�t�{��ă��v�U�"|,q�d8U���u-�h���7����܀�#��� hR ����'Δ�qTX8=�0�YbG�>l��Ô������p>ѽ��P65��6��ǖ=����$���#��[�o&e_/2�_8�����$٭mpa-\(���.�9=H~��Ob7*�5����ؔ�S��Y����;�C�R,��\�z7{�s.D�u�ȑ����uhyv�H%�c��m��3����0z"A_�yG�4]�.�����F����	�M�V�m��#¯��Lֻ�2�(`��}zW��1W�]^���RK�Ľ��{/�Ȇ7�����Y�zVl@�]Cwm�*���ʔy���5/���^�[��xg�;��5��3:q�����=J��<�����nQ�N���wSpR7h�(�$��-KG�ɾ^`�_��U�/T#��<�)�D�=��Т;�@�Ĵ��Fiʸ�pO)2_�&y�=)�щ\E9����v��$��c�_����}$9�l��SW�5Уi�� p��c�
�s鼋���r�rJm��ICAt}��'�6��;�>&{o+ =�x�EJ���� �����2�̎������|=>`�w
GXʱ�r�Xre>I�%�na��3M���;�V�����9d�v�pB�&������m��6��^��V����120��0��+M^�|�wX ��Fi��I���&�N;�!2���?�P*1��1z�S���kj���T�ŋ�٪�����'��TE��;Cm���|\��)i��l��4��V���a���%XC�^x�b��Э=���٭�ۮ���\	���5�b��^��Dצ�}�q��C�������$)ʞ�#q\���� ����f�h�?����P�����o���*tH�X�_=����ͅ����ȵ�:�[��R�ʲ���Ӄ����OpB�"��Vʶ�����>F�M7���Fx�$�S)z��<�rp}5���S��l�E�r���_�!����o���)�"�6�֘�U�A7�����;"��Q����
s�X�?���20y�*\d��U3�dΆs�4�%@���b��l�y���騋�r������fZ�0���)�������	��۲'����9kXդWh�V9�oA5��{
�I��8h�k\��1�).9Bd}�b&�!�w�	����^Dgd���}�����7��ߧ!����9[77D�}8R()^���	�܆Y3�G��o�[��M���"/\qb`.�sZ�i�g���T��RZO+�\������`;⥼&4�������~��O�$eO��.*jA�����꿅�C��^��}C�Z�8��dv����KiUL����K&���O��h\� � �4�x�Ӻ���y�=F���5�����zg_X-m�����m+i�'��R��\��|�mI�Eb����(vJ<:y��	���S���|���j�ә�ּŒ_��/O\,���!�ɺ�s��6�I��r��oJp*��#.��HgH���pL!�8��Rļ�7̶W�M���zx�xn: ���#K�_��=�ޔ��5�n�73t�e�B(��VtZ�����m<w�{� }�=�tr�7m.PrZ�>pr|�1n+��РJ�s����셲"*+`G��a�c&&�X��"�g֩��1��
mK\3�ލ�l3rL��u7MB�����^���(Ш��:�`*�E�?�-�Fϡ��V�K�hAO�Χ_�3�����{����h�U���q�g'��ǖ����� ڣ<2�-l��Z,@����Y�%�R�k�%�ܺK�R�b��gD�����0��R�����ې
<�B�>�L�^ '��_�҈�D&��7koE��:ỉ5��d���'�Wv�8����J̕`�~U�no9Ct�HE?�4�h���s�AGf��j�l��V!���<����ٍ�#~N��su;�<V�jH�/�\��ܙ��R�b������4l�Y'd�e$�ڠ7L�0�-Z1���w�s���.�}<������եT2�(W�ʊI�LfC��		��ҍ��N��>�Q���P�U�\�'Aa�1�0�8�����P�(j�GC`��c]�W���RPI���R�#�-�\k����K��������i2@"P1����!��V�|�at��ַ�$d!�[����Md�UfD��ReC�6컪���Ӗ^
,12�u�#�Gl����"���P��Du�����4���AV�S�OɌ5�������p�l����S��-t;*�C���������U���3����Y�V�!��F9��y\����	�̔_T=�#u{�1x��@��p��M��:����g�O���E�������p���OsuB�袁���u®�L'���u ��u�Ї�Ad?��`���w�e�͔w1��&�O��I�$XR1+1��J�ޭ�T���5���NǤ�Hջ�.;4ʊ�i����#=��(I��:4{��C��aāpٿL��ފ���$�@��L�r{I樈^G��g����"�C�3�Z�k�U%�G=�Q{�A~o�c��FM��ВT�<"��vf��t5X5�vd�*B�g��o]�NzI'-r=���N p�h� )@���N��;�Q�� A��%M����i�d�6��,��0�s�����Ll�"ns�LuQ�\�������c�0]��-��ٓ�Z!�jܰf0Y%��<A~�1��O�l�&͢��W����%�fIW�:�~����"�p���)����k�+h��y�7F-04>\
�F�>����$Z`��×���?�&�7aW�sq�^N @ �b��n�Zf�'0n�?��`��Q4med]i����u?�%&�4����o���3C	��穃��}ڷ'�F/=Z#q�x��K��"F�%�� pwe헕]|�<�٦�����od�v�)|꿋�ls:rKE>��pJe��<��-�bܬ��{8���Oc��r�mKQ}�q�& �W��o�	�9��/c�SR�~��u�[����K���Ȯff�+� x��p�0qwz�<g��w�=A�h<��z�"q�k�o�*3)���#��*u<ʎ����(�����e�])Bt�p�Y�kv!�:k��ΙZ�	��{���Jh�Y�	�RK��bHZ��5�
J�bDj��˹b7L�(�H���aAjS���:�l��c��
�uW"q`�3}����F��
q�hi$x�q�qѨ~�?4���j���`?�t���-H�r3�������n����ܸhly#�m[�~4zW%��C�_������?�?�FZ�POD�\��A ��cͤ�*(EE�(��r|��6�X(�[eu�b�@����M�*�̆}�ܰwX�� y���ؕ��v�t(�R�Bީ�W$�MKF0�I����+�7 p��8�./��@,!�w�/�'���z���c���c+tj+J\>�������k�Z֠m�A=_���WӨ*��m�=�z&G�,1�=��++O'��,��֠����b�� 2}�r1^~�q=���
6D�qݟU�J�~_�2qݜ7�'��A}:���N��M�����p#��Y����J�>o�����n��-u�h��$�a�-�+����5�d�rN~vQ]�qр���+R�2>���*�b_��2R�%/݂qn3�	ʾ�F�
���[f7�a����i���.��#+��c��0~<���������Y7v7�((�O4��kU�,nN0t��U)�NE��5�`#�ϖ(�2hz�)*T���+�TɿH���(zN"�N�B���a0�a[�.���v�1{x��{�=��K�Z1��0+���f�����Z�}#��¼j�M��
1얳����ő�O�l��J�ɇpp-c�M��Y<��"�L�5d�̂�-չ�'G��X�߸��6�Q,7�BSZ�b/kl#�*�+�ƹ�퀆���"�;��Q2*�j�7���{u����}Wh���e���i,�>��:u�� �#��jY�!D�taN!��� �i-R}�����| s�O�����!�*�/�Vo��Wo4!)+Yn+���'��5����<�o��b�-���t��FdΝ���Vk����I��-��} �I�B�1�rk7����Vv�suK<`p�.0�R�"W1�=d��0�r�s�����I�ê���!�D����@sώ��oķ����e��UӚ]��2�W�%#�0g!%�0�W�EU�Q��
<_�_Lf j{醦������]���1�uwh.0ul��`��G��e
cF�Ϭ�F,S49Ԩ�}H�d�R<2�|���_�\�{���<�G�M/A׮��r���ڤ�}f�����j�(�@�a\����c���Qy��]B
^�5	�.̉'���)d,�!�چ6���^�aυ�j���Ҍt�7g5�2̎fH�v�|V'gt�8YB�͂�a_vr���t�k��\�i�R�O��A�ɀU�6:�ܐ�rT2k�6W��$�������M^�._ _5��o*�"&$M���g���=���/��@�,����B�Ѣ���a"��<;�Q9
�/�nNp왞ϥ���N-�Q+�H�Ђ��A(�5%-2�W��[Qg] fЭ[���̿<�LS�/KŊ�
��C�9T�,�O�~Տ�(R*?�d&@��5L����tZ����Y�3L�͇�ZNMY��i��3B��P_3��kV	���J�'��1lKz��(���vݩx �����U�����@^�����@h���6*!H>�77S������Bn�f�2nh��a  �!"���돫FFu[�UIʾ$��oU�al�����������Jp=i{��@�I?mӯ���`�<��g�㏻�Y>�eɕ��_ww����`q�L��*���x�:a�\g��r�ȥkjh�%�7,�W�͑�!�1n��N�e2vH��X��6g��D�B��l�V�[bP��E%�=�j��R;��8@M˗`p�(�`+e�u���$��͚4�Fn|����M>I"��?՗�Z�D;NyZ0 �K�A��������<1jU �1���BݣZ�̼g���!��F������� 4��@ ]�Q�\B*ȑ`���p],��.ψ!�x����,Z~�P���d�h�6��U�^W0wT/Y�B$]�G�W6�@����W�W:�(NPq2P��ӱO���k{>�,]oQ�kt8�ǆ��M��V@
�\��[��ߜ{H"R��򡅙�U�5��贀�Q"�����Ueh�I�޳��0��������oö]���Q�ᜄ�LK��4��*�*�]VѶg�>���֚ ���߁�?�#R-�u�0���<�I�_A�
{��B�3�j��wr��#��8F�����.���rR�t���|c8I�IW��q'*�07�j�ۀ��Ǹ���.,�҆9=*pda��}���w:{��3�g/a�t�Y��]3N�iZ�l���|$2��T��SNǚJ��{��6v]*���G�S�'��i���L�<¦��G���`_��\����Rvz9��KQ�rE�!��3�%��'�O/E�fx�F�V�!�K������{ҙ�R�Zv�Z�(ٹ� j�9y^$ ��j�]G��I����;ց�t5���Ԡ�����N9�I�W\.xO��{��C��<q�D�Ma�e'5�����MM�J�h,�}�Źxi�6���� O��H��I��u���՚ߟR#4��ŋ�*r$Y��Z_DOd��i0Hwu�%#2q.����םُ�Լk����]'[b����>t4�����B����q\pr�_�,
l�iD眴$��'�C��a|Zzp�9�,�@�D�	�;z�B�x��u��	O$1Z�a@
��(���9���f�zR%VI��l���\�2v$Ue1�[/kaC�n|0'f;�MÅ>��R �"�ua�(PY[��<���w�������d�[Zˇu�rљ	��Eo�!��Bձ{A�x���FL&�Ϯy7�!b�yv'�[wa�Q�LpOoR��D���A"�o�Na"�r�+�W�c(�Q�l�Tӈoj���o�V\Qd���yzeⴟ��.֠{*z<"Z�H��0����q�-��k��~x����X�v�i���MZ�Ϭ�26x�o���97��%�� <v�A��K��B]]C�JR��P�-�8��eZ�}ú��1\�������<�J����[jZl���_\eQ�}��l�PF:z�Y+6ڔ�Y�ۣ�ߙm}���m��p3�9�HM�[8����X���7}W�� yTz����c�whfBY�>S�R,O]���ua���oV��*�����j�47�i��y��T�x��q��0~���7I�I����n�0��2�)��u����KA5z�/\�� ��������r4�CnB������#i�0J�%��}BܐfK��Zi��R%"i>�>�f���)���l�D�ve-:��C��8W�C1ҳ3�$�Ob����&�(�JJu!]Ɍ��ޕA�t�o�����1)!+w���� f%�rG�N��挱�K�2������������)FI�p�t�x�0�	����������!�h!����@%���C�_@�ai��O��i!n�8�ƞ��^<�VAȷʚ�^w窺�����.>y���b !O5�>AZ'��i��2]��Z�!j�/��>���V�{A}�]��Z�X?r��D"'�j��/&Â��?�w���Vu���1�O�q�y\Ĭ�a9P�x�hC�A���o8��u52��V�3�G���Z��<��K8P$^.aX����~ȵD>��-�G��NS�)UO�ױ�i1MC�
9��aY�)�+c����u��.1�cU�Z�'h'[�mk��;Z[��c&����W���z=N
?0?���y��]5����C#iO�iq_8����%	�l@�B&0�4�)x��l��m�b>�\�Ʃ�Z��k�?�W��AR�LE�mWm�	��lO�:���Ψ�YNE��,@�]XT��ξk0!��^H���Fd���JED�Pߜ��.DIx1"�B���I��4{�I��mx�3?,[��[�ζ'5�VfE��B���
GC�%������Æ��H�K��In�x��l�ǣ�w�<���WW8��8Uq3�r��H��q�����.����@�Ű4&E��y�R���y��.����:@�
���g<�t7�R�7U��UDU����˰�����2ũ��7�orL��8qC�}c�����~q�I;mx!w�Ψ�nI�Z��A8��X�|U�����-{�_�%��`ƃ���@�g︿<RA�?4�1| 9��iH���F 4+ 94~ �-���U�BʹnU
i8%!ģ^����MC���A�M' �H��s�6�;I�����m}{��-�.s��&��)!�����W���9J�{}��,��畯S�������-=�ʛ�'���R��jM3(fzӕ�=L鱴�IQ��m�䶌v��r�
D��K�惂>^yԬp�p.95JD�C-�i�WηMAfQ;��6�,��	j������6]v^�[��G�r�J����ƟS43�e:JZ���~"�a֭ɻ���E�<�����2������T�0�$��c's]�c�����Z�)�w%b�n��ؠ��e�m��cL�{���=%>��T�q*m��b�Q���o�)��A��Ns{>�<�������bjt��0>V@�e��I>���i��J�շbu�-{��L�`�D��q�y���y7��[��M�O:���|�O;e��/��$��.��v���~�p8����6����M��}�s�Sy��|7IZ�T]M�A��@ �}��f��f�Є�D�б̕BВ�j	p����Q�^޷�2����I�$����bws?�2��&jf���*ki6݃#E��4pFR��=9#{��hM��(��:��^9Tm��*�H��k�V6ge�+�i�4D1�ݍ�߲��#
��C�@PU�����_��l��嵖3����h�(7C@����x'�e���#͘��-m��dyM7��f�Yn��> \�v��m����C��a��גP�q��j�j� .q�1���^u0p��� �)O��7�ۑ�eP��4Ľ�f�,��F%P.�����W���9Ѐ�z�Fb��O�f�،U�r�3�~�;%x`x_Xs��Hq�T���G���5g�_��ϱ�����Lf�h}��4��� 2�m��d�k$M%mƾc�_���OLqd,D��ġ�I��� ���k��t2��]�擘��1K� s F��gcց����U���e����H@t�_�Yx����V�`��%:�IGH慺!&ة�]ނ�g/�bݭ^�>8M���2[�O!BV8�n��uW����ɛ�	x�b�oG��j�ћo���_K��t���f5!�� 6F���vz �ɠ܇u��ϗcy�)�2
;���6s�Vkכ]s\�B4��Ib]ݵ�7��;P1�����J� ���_���qg�>��k�V��՘��M���C�R%�;�\�׋k$w.NU������胁��]��C�)���ݴ�]�!��MC�肒�A`���r�����S�<��{���{�Uz`�L��k�Q������hp:]�uKF[ɰ��J�vhг=��aݘ���6Ǉ�u8.����p�A����Fh$�}�hE��XU+ԍf����J��z-��b����c\er�ى��3[K9�<vV��Eq��к��-8;y5G7ba
ܛ�-O�]�U;���Q�Z}�1��I1�0g3��n]/(�z)��CVr��%��@*�md�@��� f��h�ZU^�K���C5�dX���q3�e]Y�;%���2?Qȫ&Z'�EV�Q���u^��NC� ڀ�<�'~�m�t~eO�,k����D�ڐ,)�-ς����e}�=�(�nF�h3��([��^���S8'	j�2��BsU�������g�Ώr���3Ul;���n+~N�UE��
n8�0�j�cq9��l_Ϣ�4H[��Ig'&�t������}�($�B�Q�V��=:��]L��=b���)P$���|kKqĽt��|�����u����ĉ�3#V2��6���;i��](��椗���p��p�����e���H@|_}��}<W� ݃I�u��}�b@�[�:�˃�mȜ��9���k�=����j�T�d���:�eȵホc16�v܎�("f�f��ǵ��#�yus1�D���Y�w��m�s~���F fL�����(ۇ�e�2\�Q��x[�����߄�P�7�H8�S�V@?+E��7�1Fg3���,5"&�[�� �`g�_��,f�
  ��*���d�Z��{�K��;�m2�,1����^/-��rO[�l�!�����^GL_��l��mN�%�d'+	&ce�����輝f6���_AV��\���#�����K@�D{c� ەC��ʙL��R��g��͋yة�3�Jt`�=�9��)�H�si��������a��Ĵ7u��[.�bN����@^��?gT�L� O{�&�ȸH�|���Yi��1�!cF+_놊����2�(�Cn�sNP(�7����$�0�߾9��7X �E4_�::MTG�w8?Ԝ/���_���M�oؤ��9]L��H4���7�i�8-�G�h����Hg>�!�
�!X�Q��t
&Ǿ������Q��'pkS$f�'b{@9��٪�i��Gڼ�}�<�ڎ:�/�*��D��(8���-�qA`Е?�����V6�����y���ɹ"�tbE�P�c�nT�(�o�NA����Q��}�4����� �U��hc�v{U���EN�7?&�N���-'��G��nΆ	���7rL�u)r��I,X'�n��T��)�):���(
�T;��C��`�������<͸67�@k�
���]�}vl�߲�j�h'v��TuKd;[�kywc��b����gY���:6�]g��Gd}�jfx �Kf=\5k^�۬%*<�QrA�.d~��٢�BV�~��'(K��LIh@��	�$�^2s����%�X����r��ɧZ)N?��7c�"1(� Ga����tL�$����ѽv�*F�ջ��݇;,�^y[ѫ���"���ƭ�W/�7�k�F�4�%�E\�r8�K�ygE�asetV[����/�hG��7��e'I�]Q��?�l\��� ����b]Q� �Z� Hq�3	��}��e��]�}w���W~;blT���k4&7�\l�x�^�@k�~�I��T<o�){���Ϡp��̥A�`�W�z��_~6�`��І��'B�@z����wc�����.�Z�A���2��.�M-���Ĭ��&&$t�_)�|_��)�d���w9�{���n��<�8�#u�ޮHX��r Xl��z_aOYgǬ��g��]���^g8k{�u3#&uM����l$(�2"DkC���Et���U����[`��X|?�n�4pi�Y��O�'ύ���[|j��\Q�������J���h�}��7�s�.�(�E�~uǜ..2 �(��x({�����<r�4���a���)�0O� =w&��\�[3��iL�l!H55v~���ɟ
ڽ���T@�|.%�$�9lh� �$>z�mױ�I���K��$���B�*��Ƞ?L��CS�I'�T'�f���F�\u(���N5���hƘ�&���&�YI�%����e�O���P��T����RC�L���P)�M�TD����IZV?�,<K��eQt���i�[g^�p�w���$���g�F�[��4
��9�a�s%V'o�C̏�"���j�ʝ��E�/���=h�}���[���
�pL��ja }��:�c���jiN�:agO��hiOJd��4���F#�'=�n���0���ϻEL*�Xpp��Kp�?�io�֚�_/Quw��b�y3Q�10u�O.��ԝm���jq���M��6�(	�1����uٽA�)oJV�?l+J��pyi���,�`���!㌧�n����]Hq>W�����{�h�����1*�F)��l	��v���1Hrޱ���Ws��~������|ء������d]��}a�gT%H98m6@�<t@�!�	�,W��7�è��xR�!�yt])]�M�Υ�g5�R������, ���U3+J7��jڦ�k�ƒځ8�nm��mZ�cKbi)�p�JI1�?�7W�*Z[y&y9���B����x�o:o�ք�|zO��>���&� H-�9����� $LI��ո�����t�d+b݈-$#A�&���͂&��$b���z�R`3�,dx)=( ,�:�'uݲk�D@V�r_��zMƋ|����d��W+XuY�S���fx( m����I���Y ���5D����?|g���/��P)!��g����'m �!M�.H�U�pk�52 ��=���]�Kb�š�	�uíP�_����2w����uRizI|���G�E C �Tњ<i� �ã�,�Be_C���u�Y�?Q��s��ťO�����'����8J�H��A2����)w-�j�@�Bâ��l��3�c��I84J�e_"��cJ�c�yfE��h򁒖aP���|���,�x@�ld3�b��DR������^6�8s�Ч�E~��q��l\� )=W��ޚYX�Y~@�C��6L�^���I!�qɽ�혀�����B+����-��Z�Ȉ��I��Se����*8An��H*l3�z�s�: �c�լ�o��!�ºz��.�ؚv:����1	Z�Q�+0�6NIľ}\i��(Xأ=�=^�ia�	�A�A(�hkc0� ��>3s^^�[J=ۛR�I��m�jo����FdC�\� a��v�p���t�W=���Ka�{��v_�J��)4�7��=p����m��zC ��(��a��v����I�+�R�"���oػi�3��Om�9
��s��йtp�Ug�d��z�_7�<��Sۊ)r3E-5`�^'�J�e5_�^}>����� ��+Y1�DW��~;&&n�Q���%)$%�<��̗^z�'V�DDW- i�مX���H�Ƴu,��m�w�T'[#bcuZ�1����m0G�����"X47����){Z�ڑ;U�~Zӿ�eA��z����W��2^V���#�&���۴�o.=�keo+��I�>bN��w51�p���%OmD�v\To;�ͪ��Qs( �X}��O��;(g�W2�^aM��S	l�0�/�)��z`�fM��HR���1%�<Ի��/����L���Pqo0(	�i`�@\�-��,E*��Q��K� Ɉ��}�E3`���ʀ�	|�^=�����Qt.�/V���OW\�L�l�c�#��mTQ�/g�QL���c�{g���>Tm�O���ـ.vBI�K:�/�Zw�7�LN$*��x�3��Ϭ��à�_Np�R�J�M�/�T( �������U�"��2���0�ɮ])��X����n�zi3F�=�}It)\\�6o�b��J@�t}��X�s�++���Ga��o<`��WV7�� _s�$�>f4*rj�r�]j�;�!�bލ>M�@�+��_��;��%z�k�^E�ac�{�^7����������GD������W#�ݒ����c�jسWi��*�n����5.�݉����.�Nk�q�c���sY�?%�ґ�7�#A�X����׺�;fH)dV��=�&@����%�e��ѣ�qLA�S��k��U�S�p@2�#��$[嗠q�d����u|�@�=�ֈ�=[0Vi�eg݃6k��z�2��~��� �r�	[���-cΞ?�+h^=>����dC`}E��"��KK|�"Jao�!:p�|ͤ��R�q!��s���u��p�Oww򎏻!�Ka�L�\5΅Ō@r�M	ޜ��l���8������B�m� ���U�������c���ƫ�WoT��1!�h��:�Ӫ1A�}V��d$@�S��X�_Ҫ���B��ȝkMM��[)�p1�Xb�����*=�uv(G`d�.�?y���B�@˪P$�9�M֑���ܽ�"��TUՂR=#�)7�uj�Cz�nK�b:s�jl��Q�b��c���X	��\_�j��9&%���_裣FT�8�6�h�F������Q6�|8��Zc�R[^��p�]$��mI�o���K��s�����-��E�`1@�n4�N��F�_��2(�Z,/��1q;�H�<���s{l8e`^��}Y�����296����aN�+E�����%�D=��~ɯN�z�C���c�3>K��� �����'�9��-��myk�;���a�̆nn�N�JK*6���<M�nCfّ���c��}�Ti�����nC9q�:e��$u��+f����`N�*��+���Fc���W<ov��]d��(���uX��YiA��:n��jʇ�[x�i�|�,�����܄�#膣h��b��Y&�B���Xؿ� {�� ��_N@�\C��˜��x�B�IW\��;�F�F2�b�j��,�.t�^(��o�����'+k}�s����2�~���G&xs��}(��ۓb��/� ����B�[�{��7̀(��.#o�V�DI���_3��0R} )�@N��]�T-�D�r#0��f,F<�)PI�Vz2��N]�pў�,%l�e��2��[�f�Yλ8,�&�y}]���Ffa��ы1}8�
�N:�����uن|͇4�[Nb2�������o�/�|��lv��&O9��q��d�W�Rbd���=��M�"�@�*��@��������ނ�9���<���=}*�����H?��*ۑX���I��.�2���b$�Um�A�q�*����r+}%�1;�h�~I�&����)�(�#I3��*��t�B'���-�Q�>yU���$6�P�`I6����R�"0�>o�4��<:'�#yn�r��Q�z�ҟ�L�܂C��p�8��`&o�ʴ�Ű?��,d���;��x�ЏZ���=)Î�1���
���1�{ذIm���QV�L��!U9*��Um��-:�1]��b��7`��<g�.͙H�)��e^�=�Q�%x�BV�ʝ����|�P��1Z���@;�l��?j��gbAH�U(�����.�SD�Pn��K��BϠ�ͪ�	�`Q��K���=��b����rsM�(*k���jEA6}w#ڪ�w]����#c�z-2���y��<�z+oV:���e���>��'�������8$*���MY]Xv�ab#�r��#E]�Ǘ�v��1�G��G!6�)sK�b�ih�����*�	x�L|���]n�N}�E�Kb���f�J�#I��K�f�GU���v�gn9��5MÒ;�����<}&j�S�ڦ_�}����j+J]���T�Xq�;�Gm���/*+�/��2��~d�*ڔ�ei{�Y������)��Me�|Wk5y�1�W=�t���S;�&��L�#�OL�Kw�����_�����A*���yk�O+�rQ���>3��Q����׳�u�x���[KGW�wx~�E�1�����;�"�IT**�~x��9к��1�'i�1"�u0N���П䵓%d ���fj� �tE 24|ޒIk�F�G���]u��$e�_?�w(]7!J1 5#���+ �8�������D/
!���Xɶ\Y�޹���X'
sJ���WWi�^i�`#����Ԇ/^v@���;J{p��mC_E��;m�� ����@H31�j���ތ��/r�Rfju��^j#�{��@uN �Mo��d4���3��  ��A�����w�oF���p����T��]hK��beÅ�5�z���������ӐO��N���ѿH�d`��pm15��1a��{�C�mOx�9|L��f�Ԃ�ApU�l�97���{��>Xz۴0���eY%[V�Ce2tEU�`��U��P��>�:ޣ��f\/�be����]Ƚ�I땭y���:�j��nD1E�_�2C~� �ĉ�L����RW?F���QL'�>�k�i�M� �Ȋ)fpr���rW�����맱��-�e+���Z�^��+4��]�	j}N�Mue����)ݓ�]��[�ӌ�m��H��bBc�-g\@-�ídY�ن^��5F⡈�;���3nN���;$x:������(|�nʊeׯ��[�苽���9꼌�B� a{��o�)���,>�~��t���'�7b����=h�u��_�������>��s���m_Xɋ=7��dUZ���<�_�n����mX�_!��V+37�7�v�^|B�u��륝p��]&�c7:��ǦM߉n7~��/�an�`mQ�[:�8�7������P̄�~�h�G�����u�A[b)1��;��f���L Y��{��t@'�gT��'$�&�`N]�����7�_iJ�@����g*,��`��(�V�K21���A����?.X6|9��[<g�Xbkb������trm�T�+�\�J$���#s����t�	��5ZfM���x������Me^�eL ��h���L�)z��/$>V�E;���	�S�����[���͑���� ���*��+@+�(�%)f��w��!�J��x�kh����+�8ϳ�κ�?c�T\���,�V�"d}��=��Sf�pTI���4��:���� �Z���~vpd@���A��p����Ě	!���� ��>j2P���H��q����,� �� D>G���j��*+'U!2��6�΢H�ͭ�ދN�c����[�-d�Θ�5�~6������tjz$�8�d��]�Q����\�=�^tk��k�]�o���r�B�=��zN��q�}��)]��Må&O	NNQ�r�9�限
O�F�6*����"��b������\U��g��{3�����r�{�F���Ph�IvL�=�
���.�c(���&f}���d)��K�C��WI��O)>W��!4��lm$aq t>ܴY!�h�3�}������{~�Q�L��@���	l�[�T�}��賆�+�Y�&��5�9�%O�Z~�Q|�^H�P���
��t��i�5��ɱv��Ȋ��T<���i&�W�n����2���������� ��J�G-Z@,�\N?��.��`���Io�l��S�q�eG�S >���9F;qض�h˪!��D�˂��N���3����\����L����~	3ʋ}������a{������A9�]�6����R-�.�2�����J��O�n�o���.z�?�|�Qv��0S*� ���>׮�QI%=3,�Z�@�+�����I���n}V�^l�-6vN�XL#x�����6~�H�;�b�ze��|��R/�ύ7N���>#yߚmA�r��]���l��:E�:G��1�PcA,b	�xD��ߝg˵���N�1�^�W�(��{��$?+�����S��k���4i�3����ő�]�պ�&���*.�����|���� ,C?���~�ϊF��3w��ɷeC·�#m�vaޓ����[��uQ��4+�I�D�1��Od�������Щ���#��a�becԀ��}���V{�r�2���*T�C�7��|]�S��tF�?�lv��*�D:f����Uq/� �g��p9*�0�c��F� �G��@�����0��;���oK����k�gb]��qS�y���.�)�N�o��)����Д���P ��2I�=2(%�SM�sB8��w���W_8�E�J1�{9�i�%�t@a Oh6��Eo�y�l�=/mUgٔˈ�0��Ψ�ҥ㍔�g⬾�={�9z�GK���&�A�ݙ,<3�����Zʿ�tj&�p޴�%�:m������	qWd}��7KQ�p��5�Z�=���*'e-r���n�,�_�!�Bs:T?
P�R!��e��<�.��;3n
P�J>���͓�EΫ"t�-��t�/ۇz��u69�M�$��{���~V~����MC3ԛ��[-�@�J�3��/�8�)�Ѷ"^�t�0�.h���,�q��	�#8�b�G�pSBa���g�5�daK�N��ʣP�<����ڲ�k���_�ez��
R����le2;M���}��z�3=��nK�Ik��ZG���1y��������H������<�Y=�o<TxBR|�]Eh(��ܾ�y�V-�o�RA���;l�`��6D�R̓�P�|A�v}Hf��ứ�@b�� �)_@�SC�͆�{]6B��F��3���O�5���g��xn���)%�/ʕ��m�(�N�����Ӟ�v�С�^&�
d�$H�N=7�����iJ2�Y���̱��z�i�s|�wEB��_�+�� ��M�3k�ý���K>df�b��Z�fm��l��ֲ�G�r����g~��:�B4�jo�Ap ��l�j��@�s'�ϡ��4���-@̺��Ha��I	� uS	���GPӵ �!u���B��R�-V`�L_
�2�D�s���?Or˳�+���c���c����M 
0��G�H�X���H��'���ql`58Jr{l�����Ő�e�c;�X$U������t¼I'�;�]�|��y��(�jM����$�Z~���pW���^�N:ɛ박;l0U��s�W5�q�nR�D1�t�g��� W"�	_�frU'��ޔ��ܫ?"��|K.��f_d~����ia��,�u�vq�Ɠ�:��5��%(4I�]`ˬ�#zVp�,y����T\~9A���"ow�"sD�b��j��5nɄX3���������ڡ�S��=�����e��^�K��8F~\O�0{�E6O����^�|�3�m=$�M5��s2�*K�t����`�ls�gg!L
aJ�y�m�4`���M�cl^�6 ��j�v��Jt�fC�>GAz����<3� ��nm�A����r�����jwve���~n�G��W�������p:T�ަ�T8x�!K�PL� �,P�t�$L�N�f.��t�f��4�78�9�v�y���[ø�KA�t�ʽx�r�Ζ;)�R�p�T�,B��g��, e~�h��»p&�9 �c��']�Ú.j���v��	�M���(�(�خ��gޅKC�sX/i�����4#�\ �cyU�7d=V�O�)�H�i"��g�F>Eh�D|��Q[o_�?V�M�?`L�6�>����Vj�K6�|��N�������E�s�k��0�z��_�L�����,j���@��
DA�2@��_j驜�s�E�N�x��S���9�熤��V0yK�c���?� v��	���v��2G��:�K�b�=�1��]�$��_R���P�Ƃ���I���]#����GeI�����*���R��QeN~����
�W������ �I
.2g�.�0ܓ֛2�SR�hoj����$���?���������"��r:\^�~i�|ԕ��
r(8�b���	��Kcl:��H!��	ga�h9欗�-���)xM@���H��R��0��$���F� ���� ⥄��^�Z��¢5�J�K>[��~�`��m��*xבl��� ��������S�7�����WF��*�l�1ALgFh�� ��k-����nj�<}�^�`��_�5	dT�`T�QgP8SP��#��.&�>���F�Tk���=;���ߍ�re[�֑��M1:E�O���%�վ06�=/�T��Dw	DϧT�M��e��q;[��w'���(ώ1����r]��&~��u�:�� >D��Jx"��szV��1:M��jQM&�_9�38W��FR�f����s���i�H�$�0����-��C1��Y`� �닟c�iT�����AL@��`8Ϡn�5�Pˬ]c	�WÆ�?1.F��C�}��>��	*G�gO~@ �c��E�����k���4E�װKԗ킒c���貂Bɭ�2r+4����T���D�G
�D������0���=,�VW�9R"��M��5��}@���7`�?�<0L0��u�ĉ�}�h���`N���7��Q�9�f�ȩ�#���@k^@&��v��5�Z�i�$AD���`~���F�Tx����f�����ט��#�ՓK�-�f���k ŏjnt��2�\�X����Ȫ<�����}��G j吖Ǟ.�Tp������-1>z�cu���X;��G��/��5E���'j�l��˩�n:���<��o�I(DO�����3�*���s���;��ok���� ���S	��<�b��UWh\�Z�G=���z�-�����~��Y(D��7��K����y��������Z�5��j!}0ȣ�'�qzκ%��:�t�7�������n>4z�(��;��&�P��Z܋b@*��RN�ҷ����|Œ
�SF�=��J|/��G����|����>�U�f�8�e�q�歋͹r h��
tH��i��9��-��Q��s����}�Zw�9RW%"_�������~�5;V���D�O2YP�Q�宓�0A��v�a7:ܚ�.��U�^y+�y�����٨��)M�R��6��ݰ�����T���E�!�q�����+Zq����1��@a���'�J����r��Q���E�ģ2�#�P�f�8
�_��wԎ���M�c�>�ƹ��b�֣�J��"�*��v‰� ��@�� d�MS0?柌�8w�4 �0���#'�F��	����v^$�y$��dz��?l�;�z��}(̨i��y]c���Y�J�7;m�-�B���$X��s��Y�a�ŃJ7<�MM�O��ʎ&�J�|J@�٪�uj�^������L�u	H�ֲ͓C�kKOa��ޖ@�Cc���T��D�ܡ'����q�ۥ�h옔AL�4	������>��y��Ui�xc[�n��*B*�����X�����l�Zpo�k��?:r�9��{�^$�=�x;����PY�A�k��p �tqK���H���?�\�w�P�DE���p�-�A��Җ����bߑ��LQ���l��=��JB
Qv�{���� %u�Q'�՜4ٍ����4��c�B��OK]�>�vP�V�l��@���}%�G{��e�x]85�T3�z[��\�muH�U�Ƨ��R�FH7瑠RW�6��`���r�Ս��B��fw�r��\��t�+޻��>��hd t��1
_���g����a�(���b�r���]HX|��b���p<�)���P�4:����G��lڹ��53c�-���Xi���L����B�g���a�ψ&�a��m�SE�+>�o��օ݆ ��m5E|m ����-�3������5�H?'�nݣT"WUE�T�KgQ;���Qh�Zjd i�1���� ��ۉ�ݶG�V<�Oד����sw�G�Wlb�
ݱ���S�C�}��}q<7���ah��)�]�M��+�����n���B+ф���'�gIEo�c�:#A�9�8�5Zo�He7��÷D�T�%�SI�s��T2����I�C�b�r���w|�c}x��u+�Yz,��\��_^bW��CYC�caF�pw2�N#�Ӱ5��J!�|.� ���ss�n��������|8��N�盖eQ�+�L����g��ߩ��:<��{�?�*��d�"Gz�h���=����jD��W������zp<��?�;��N�z���Q�Z�.i�Dͨo����v��c�NAc�@Ti:���x OWz����W��[5���u��\7C����>���	;�}�ڟ��No`�����x^s�Rv ��"�w���
���RN ��DQ5��b�i��)�:1D2PH���E��zDO����J�����ȗ���x��H���Gz��:����ge!6Ǽ��6-d3��v��_����ƥF�Q���aaE�\w��Q�u% �x��.��d��J���ъ4�X��A?�0���2_�F�f����H��Ӌ"��%�b�=�	<��y�������D��9�-����3蹿������^�7��<�V%N���ҋݘ@U���Peݷ��cq�J/c�pۼ�Qj�~��5��o��!2��⯒`�7#�䞛܊2��\7��z�'�w�*
g1����-d m�Tׄ6��h�Wc"��C��]-��Q��d<D�G�"
�С4l='⚣�4��{��}
yt�PT�C}�L�l��P�Y��h�ǰ�
�����k��m��A�*������R���S�@K��Dkcm��j��u�4���ٝ��=����%lŧ�8+pFDtr�+�
�Cًx{4l�]�m��:|Ζ�J� Dx�B��I�T*� ���J��o������?t�M�G�oOjц虒+�Z���;s^M����]���#,x�2���X�x�f�/y���xq�T�Ԃ�r������ �@	iirx��(Iۄ5�m��#�B�9���f��Q+�y9����RV��lL��ڄ�Ŧ'�����NV���Z��W^6�����U7.H��*��0T�ޑ��Gj�NVǥU�Z0T�ѫ��~M���w�U ������5�d�����@v�S):�]~��:��61��o* �S��%9���
�o�;cL��\{���#���[��|r]m�1�����2�g�s%O�޶��+�!�.��5[E�� dd��c\O.R��9���W�f9�*d<l#}�����ū�����gs���Q�UC(q/7`�����ѷuJ���P�Ʒ/��i5�D�XO�U'	��[��q}�F����s;擑�ؓ�6C|RU y��Q����_��Z\wH�ٌAk ��"=B�ߌ�Q:��m���\t��퀶�]o�
c����ҕ�N�P��E�֌�0�;�z��i�^�1}s�\����p���U�0�UA��<~��ϷyT���O�ȏ�Vr����~m����tLA-"�U3&ܐ��u��hPgx/Pzli L��lǟ�	w�'���ֹ���r�E-����񫸐�F�zhW��	D�d�����>'�����Yc��vG��6K^&4�����v�P�&���q��3�'��}GZ�sb�$�& Ce��0���"��*i�ܟp6�߭��X�.-ݚ���F�Ma¸�}�q�̉aӦ4OyW1�a,�r�P���ND�xWE�]��}�8x�q]%J��v��+ݖ�)�э��_�|U�v��H����ռ�W(.�qл�/	Q�s}��|1��{	�f��T>���b8v%���i(x��;GZY�kX��'�M��o"��,ֺ���Cc@�d'%��¡�:�np����-mv�H�<��(F�n��Vd!��Y��g֥of���N,���]C�� ���_4��iC��L�|���ڽ	#Q���1�H�[\&/����%_�=�^@'�?vϖq��FN�����>�TY�רZO%L]86Q&���E�v�ӄkZIw�V���r���<b��kA���G�a1μ����Ti7.h���
�uK���ub����>ʜޮ��]��l(�b��n�o�s0�*᝹�ˑ�v_�x1��b�d��&�������n�����W���~jS��z���f}V |�}�/�XJ�"�3��-��T����T��
���P i� b�.#�X����4f�8G�3�&7ư��JX'�5 m� ��HZ��V	b�Yr�72�R�}w*&fx�Є���df-4V�E��Q~��W!�(�u:�w
ط�L܂�߾MYG�t!�V�L�♠���۞v�z.I��#�|g�����
�I��B�o��� d5��\�K
���~ʕ��f$�ev�M!��e��6HU��l��F��u`�Q#T+�[`����M_��a�o|k�Z��\A_�3�,D�2��U��+b�kʯT�M�'���E�s�>.�u�r\�Ć_������u�4'�F"����z�� �&����b/�3�ۂ��؂�����Q���ďq���}�����q�be�뙚5T}6o��f����X�?T�PŹbN�5���L�6Z��|;�� ���mw�T�C[#�ui���{j��������'5�<:b���c�����Sx�!��(B����ޢsm���m���,K�x0���q�U!t&�C�is�O�h�z���G����M�!9d�/^������?�GLH:����|�>�M��ym٘��"�y�������{ɑ�\a�U���L�Ő�������dk�\����g��s��Ⱦ�r�R�os�s��U�-_0`�iAdo��=b�x"����4��4;@��9#a D�
���;��er�ALNe�ZC�G��/�{OC�pԝ��2Ǩ�{�cB*�ܨ�#>�ó�Jb��������	�#�
�fQ/O�Ï�;��;Q|��������"�->����J�����ZN3K�����'s�<5Y�ƹu;w��A��=M j���`g�E�F>��?@��T3��W���A~�x�3耖����H�!w�&N����D��?V~~�_֖,��}��~u��E�MM��zT�P���/��]lau<���y4W��95@�[	*�]&n�b��Y��VB�`�o�)���ύ�*���/�<H�d�+ �^�*O<W��l���	}vnh�d�|i�'�y�
�em���y��{�����+T�eU^�FAՉ���FT$��d����(�8F9礨`�F/�M��]���sK����P�\V�̰������;�ϝ��`���ɦl�K�~ Mj|z1�Ғ,0���B]�8��4�b�55�������(cR��:�l*M���3xnV���qB��	�C~u.XZUD�u(p>�*��,V?p��Ν�.:��Ǖ/���#�_���%�C߱�������K��2F���o���R���'�=�L�K�n���2�;���R�!M:��tn|���b}���:>T��s~s��sN�\:���<�g�BqJ̾�V����2$�|;��s��>qe�N!\�V����B��+-o�@RE�卵R����6�9��,?̗�ɔ�B,����p����H �����ma�ԾG����(��S���I�����Z@����S���b�(�����dk.��@h;_
�zJ>���R$5�\��0���t�^�q=;�aK!�Q&�m(Q�D�N���	��
G}��%!�|��9w�l6>��)��F#�H@���f_N)�~�L�1��q�M� _#" \����\G�D�ھ-��[0p"ސ{3�#ʹ�M�/R�e����Y�L�G~z���ҥ�fT���C�#%��m��ƶ"/P9Rĕ}U%��ۭlդ�Jڱ6s�-	�d�(7'jsխ����*����X�ҝYj,��ݒ�l�<��i�>�NY"�A�=tkx�0N���0��G?�(::��XM%h���g�IK����ڙ�9�T3@��U��֋$�xU\�������i{2�`�1zV,x�������	»VxY3�0��0M Ѽ"�?T��RƩ�c�W܃�d6sʥ�U�V�H~ֿ�[�(�NY?.��s�P��㉑)��n6k�2M�������]X��?�����Ww����bh�;��h�HV�"\��qQ0�C�pɖ̑�xV����U����I4�z�0�r�`���*�M�G�2�Pg��	`h�Q �?ު@K��>h���Ɗ���Mc!��d�vN�I�WA���`GUӒG�����&+6�_� ,���}�̪��l2���X)�J�)���Ɲ"rn���= ��}���"t�R�Y0�>.wcB$�
�*B��1��Q�I����;v��N���*ٗY\�0�%�P��n��48\ ��
��pc��Zt����a㻹�9�1EɓY�Q�x��V0`�O��ϧ�RG�+�V�`�ȏ�%SS�8Z�b��%.ǻ���T��I�(�3s������h�HV�LR�JX�vari�ҨGf�en���uXM�Ny~U��Gu����Ygi7O���+�q��=��1�G	��??���л����Pb�t��л:SI�{�� |�X�=	/��39��1�{��ٞلh}r�	���������1�� +���O ��\6I��=
i��gUr�O��U����&;�J�Pª!j>gY����1��E�O�#�7� �����g�������k�9�h����[�ZE�ޘ�k�7��dnH���&��J� �C=a�b��V9C:�I
�:���lļ5E���s�wt��"��^�XE	�x�$�A�PAi�fw�]�-�*$B���.��kהu�6KN�֖�'l��ѡ��N�7n9l�%��q C:� th�|�F�T�-��1���8���~ߟ�cO�9	�����p�N�ь��#(=(��*�M������L���pqUz�vr}=�3��/����tҦ��wׂ�1EY�T���&;��B3at*� k>�?Gs&�&���x����d ��ƛOn�&/�_6�Յ����8��V߰pҳ>����{*�/7��,s:� z�{,S�y^c����/����	��U���L�[�)6�$3w"�@���7Q3E+ȣ��:�M@�Ԃ�7fiz<#D�4E�������K�Sš������,6�p�Sd#0�!�����Zm+G��"����~��E�s����:�>��\՞X�!Wy��!���0�|��[�ᘾ��މ/X�W]��͙�e�a
E��]����w�_71��$�d����J�ع�<Q��H��lk��U�y�8�}��(�T[�����HT�,y%X}��"��y����rv����W{�#B����xd�G����`�j�E�0��z'l|���~�@���L�/v��w�]؏E_ uw�)�����:Gl��Iq�;ߋW��<����wϿ.]AeV!�K
��^5;��rXc����������wl�#~�~�l]����oX6��#��'������Z�|�����3�e�GE���2�������o鈉)n�`$U_�����?�c�0�`c�_�0:�z���i�=I}-��Pj�2��hD�,�[�r2��^�e�_�[�]X�ä���C/ٌ��M��6����X��k��s-���I��ߡ�_�)�>�hN�
6���,F8$�S;V#�鵤	u�?�Z�I�3i5�j�&h�c��z�TwqQ���o(x���f��MB���$߾>��9wr�k�P^�b���)���[��]#7�]���'M��(�*�8������n�i1�M�l-�>uGW��M�le��Y!T�$�a���/T�^ԉTh��ԮY(j2�T3w����e����6.p�2����� ���4n���\_)�"sn�]�q��h�N�rB5��W׏��$�&u���Q �������Ǘ��Z�>���'٠�u<��N�]�!D8�!=H?��&�&Ϙ(�R�B��=t��?̇�c{��𾣫�ƽ!���NM�D!}ձu�<��G6���;��Z
�- �W8��'t2��bW-��DրNP�f�H:�co��*������Y�t`fu�c����g�β��3�s� Ϛs�I���+%� �b�:���7az����c)䓥$�'�&i{5��:���)�{E���w�[����h1�aJ��
z� �A���-�����ECׅ���Ye;^����QD��6O*�y�aJ��`�2E�|�yI�L�Z�E�2��vh�AL���c#�p|��l˴8U�OG��ys�N	a����G���WH���o�}+�����N�$�d�f_��?�*2�Ev�jhb\	�Ыm�����`$�02���4�S0dJ7���k!�ؿ�c:��_�BV�a�t�<b���P�=#�Bk2��\[��6�g�ޕ�6/,T[�C��V�'�exH4ik*~H��K�1��e���*}1�8WiqV��Ƈ�-ZIL-���CSgo �܇�����M�hRRaxƈ���dsn(8�A�\��Tw���wc^���ң�Qvuqy��nI^�Oр�j��u�+[�1�'�(��Z�ˏb@�'~�D��<lo`�8�Hng1o��$ �hL����^�	����^pp)�S��w��9_I��X��m���Ѳ8�*�f��.qv[��5�R-���>�_�K�4�q Vc᷏�Y$}��t]
g�+������Qm�J������(��7I琻5��e2<��|ٔ��nY�sY�N�%���i��~	L�����+F�3XZ�f
���OC׬�)���Qi��҈S��O��G~��c[� kQ�;�oF��h�b��Jv*�lӼf{��mՠUJ
�c�+9�@@Tuw� �-���!�N:�(���9���?����MU�1+�5�����сL����сx�P;5��t�4*5��I���+��3����"Y����C�N٘�c�D<:�\���{��@P]����CY��?K#_v�����o��{ϯe���k9uqo�b
��1���ABھ��|1�]�ޘ�?!�3X3*����8�CSĮ���3��4���͑#c��"M+B�1!2��5#s=Y����37:����0��d���f5,r���c�J$^j�l��0�B�}93J��-/�_�Q-�K��X��%��PL�Fϳ�9�ܼq��T�|[\n��QI7!ܿD����A�b=zCm�UL�9�J�k��N�=��c�t3���(�2@N�̣�CH��RKn�F,�r��Y*�2SÂ�D��÷x���dWV$x���;!�ke��aNmڪ�T��`\���؏dἓ]�/G&�B��S�_�
�=�z%�zم�:.30R1Au�SA�D�4�*U�M��loh�G������i/�g�s� T�Ր�����!CA� u4�d�\�?xF�"��?{M�e?�:�BL��j�bA��lN�q�����\Ux$f�Nm�8��bw��,E��5ϖx�r0l�uo��:���;���ľ1��Lq��Sݞ��A6T�I��/��Z1c���b�@���L$�� T}\�z��}�K�K*�W�2%��M0����
c���?��8�p�,^hӁ��-��RW�*`�Wd����V��l�Z�� ��%6BФ?�r+E�͘S�0E"� ��q�9���̤p@���$��&Ӷ6p��
��L�����է�e�D/ŵ�:�z���^[��lz�t���T艤%�,��'�����|%�ūB�jM]�k_@W_��Ϣ%?#�Iq��nTPuOW�-����z�%��%�g�[S�d���t�K,Fe��9�� �t�:R(�R��5ek,�>����6OK|��������)����unV�$����_�bf
%��s ��S��{�zj��i�K?���򉆔�\���e�$���O��������������^e�]�B��E�]g���Y�� ���s��=��F���/Z�,�9f~�����22�!y9U�^�ƻ��b�2�s�9G[,-�{��s��Zi�f	U�ou��jNý^��w@z�.�q&�ڭi?�ʐ�c	2���#�!+u*Ƴ�t�e��T���z���r�|��"Ћ�Wf�m�l~��d^�X��R�Hy�x���[��T[!�#� ۟�ʛ���� �֦"��m�*̽�a�wxC���gRE�P=����S��7��s�G�)����Dul܏@�����Ig�Zq�f�"�]cA��Ւj���\�M���*��E$����9�>,��/.m�?s��W��u��ʎ���p͆��-���-4�`�-�t@n��`�(�[a}�cCXO�|�`n|�T0�d�y�g�4`t҄斧� ��Zeu�-��^B����sۆ?�Ҙi�4TX�`�E��������j�*���/\�0��N�.��!~�0��ی����WRqַ�� h��R�� �rm������I4������F��� x��Ͷ�58�Twm>4�ѡ�3Z4ş�i�˝kD�Էq~ѫ��(�҉�`VF3����U �5�+�91�,��o�F���w�|E"y�C�TgF�d�=U�j�� ~+Ck�lv��j"+QwGD�:
���'��"[i��yUD��1��k>������b�0ke$$����_��(T����f�����Zs�y!ŀʿ�E��}���9�B|�P�.ְ��ᲂіүdu�Ɓ����'�-ӏ&�6��Ϡg�nq�G�Y�1��,sk�7q�6���E�f5�����y��u+��J���V�wce�*��<�CM��mI	[f�K��>�ܷ�6lt�����H`ͣ���&tT���J��!\/XM��le�O�g��0�h�Ť�gY"��+��I���z]�H�)C�\T�t��;zt�Y�$�@�OЉ�����7x�j�C�E�zD?���A_�UG6���d��C��B3�6Q}�U�1`I�|k�;_�a�?�D��Y"Hr�[/�D[Z�B�>���+�OE���.�-��p:����"�=VQ��J[�������!�lS�ʚ=�8l�z�$�����&�t�����i�t���0_�S��n�XTu����Qބ����������A�E��e�������&��%�sb�Y�6g�S�J�&�)�z�
,V8���f��h^���?��A�4��6�i��J���"8���7A�d�7�2��B̍[�|�ї�̇Z&��W�]���r��&w��D$�	e!�ĭ*������ޙ�_�Y�[��伄�	<��m�KbG�8� dL ���@��ˊH��NJ����[����+*@���.Y������kSC����1�Dn)�R�j@0���I+��O�O+�[��Wz2�3�:4��;��|I�8���U�O9g��1��9�ˈ+o}]`��q�}G�{�ރD���M����c&�����6���ې�$tA�o!�W+*G��4��g���)8X}����e�	����d��;����s�P(�C��)U�A�s\��j��i��p��Ҙ%��#�����<`�{�dY�e���oĚ�%cxX��h�0R��y����G������w�%q�*�9a��o��[�>��u�ֶ�v���W-���}�U��=� &�+�N<1���|��
��\M ���]�sP�.[F�g�s�[b�w?S�&̅��B�,�[�>/u��>��������9.�Ȥ��9zO�j \�2��m�<h��}����w��U��t[�9'�-F��v0S#Hu<6g�"/��;)����t�S�R1�����&��5���;j��$v5����G��ϧ��&�3�B/�N��m�ۇ�S`zS���Z���,o_ ������+�'���)nx �|��V��cc}��H4R�0}فC�vg���DZ�8��Ӫ�Tßt�:
 h-T��G�)B�\ZTl}m�5tU�M�_�y���\�����\!��P h�iY� ��x42��!\|}�?�'*�'�"��z�1�'b��)G�М
��D׌�V5�<�����G6��$�N��ֈ=j��֙,�����%[B��C�M�OW�w��h��.�gF�*�87 mG�Z\+P�������ܬ��`��N�V'�y��)��wmS�~�K?%���1?�tx�j��ǐYQ _&��53��H���==��V��a\�*�㘋��j��Il6���n�Q��H���,�K���E�=�ss?�����m�E�j����[�d�M��ř���	%��m�~u���+���6��0���<��{>�j�`-Ǭ�4��Rݤ]bޘ=>��\������S��iFte�]7��f��ޏ���T�؇v��C��TaC�Ţ��u�H�`��t𶧔�1���J��Ռ 1��A��:�`$BV[^�R�oC�����"ѹHa.m���%��d�^I�k�Q�Ն�0^
�-"Ƥ����V.]7�A���t$�w���W�N�Ud��˶��!���m�Zg����_�h9�h(�M���f�@�*����{$=����_�95UNS�1D>FeZ��p���=@SQo�ٟwA��J���U=,ypy���Ӌ���q�WS��
Z1E�mU���x�k
s5[|O�Zx�|�DQK3[����yS\��Y�OJ��%Z��SW.�@������(r`(6����#��=��S/���2y�b;�{ ]5�8A����FL������Տż<� }Չ��hjG�+���k����`��}�����m�g�ѱF�QK%�)A�bP���+�>�� �i�?��0	 ���W\�a�@Jk���*���'rX5a����ŷ��o�ˏ���)�B˞?�`Έ�����%e�>y�Z��_#c�³"i���Y99���,vE����#ޜ�{v��� 6�5��y�W�l����)�Ȭ���ѩ��&-4s����s�Z��np�����)-j�2|kE��`5,>X[�(N�S�86�`R������V1�$��3����=4j4�(��V2�V8őn�3��$��0��ߊ!\!�x��ޏ�B���@C�� ,����P�_ qC�Fs�<�Y&6��#�?�(��0].���ȵV����p �<���h6�*O��-g�-3}3�S>��;��]��d]bcA>���&��$�o)��jy.�o�Ѝy���*N�!�F^u�OX����v�ZY���Z}j&�J�b$D�6r�#�f�Q�^�=�:r��;��Yi���>�H��d�.��Z�>�^��K�}���I�!r��y�g�ͮ�>�Yܼ8\՜6�r�7�Q(4�&Ѩ2	ž_����/�B���ֲ����}����0�Ju���=#ǆ(�>�HIς�-y�iږ�����V��(��A��5!:����$'p6��C�kM����ײw·��8����[��%�g�<Ǣ��Z�_��h�Afi�m	S�%mڷ9���T��=Q�)։3#V�"���3Əs
�>U/,�<qفo�`�s�ٱ"��O�%gRq��$�}ٞ�o,5�A�tK������I:&�N~�>U�qg5y-1~��ˁ��-&z y0-�c��O��H�qu cO�p㗗 �Lű�V ���0k���L��L���h�E�c��_c�F�gme�+��#fy�6����(ʓ�.\���:~Y�SϖOP)�υ��怢���𰔘j��E˫��>�_3�OA S��"�!�U��s �f�l&i�}�qR�`wû�*w0�f氿]��4>G��F|�l��"I[��=,�Q(*kW�w�#
��wD�[Ȭ�yZ!`"��������]!d���͇��f��Ѻ�G���g^���%(��	�O��Q��|FG���V#�Q��DI��;��E�A�di�����5�g��LP�@���OeDQ��-��h��p�S�Œ�x��t���FR������U�I^3�;�i�?:u��k��Xo����:�%�W���m�����߰��4� �_�i^?>/e^����@Te"�i���i��������VZ,Bc/�����8�]��\&n*��},�9�$'�4$�r��Y����4I�r��	 kd�� ))��>"�Q�*��Gp�5;�����:-N�:�1s�7i� ����17�*�+��2�Sew�n�cg�
M�3ʖob�?ȘPZa�j���	Nǰn���S�6p���xw��C�}k�� ����
)2����32�g�:�Kr��+�8�B[ֶ�&��P=�M3&��+��w�:�H#-'Ü _��J~��r��;�FF\	/<���������Րy���۔"�����ܙ��|�3`�fĬ�߻�ԫw��0�2CP!Gzun�0����%1,�غ�bcFU��D���դ4�u��|`t�i��M�Vqc�(�;���4�G�E"�#( ��'�ЖG���q�?SL��R��V�� gqF�v�L�P�+`�m���&#}� ��O2���L�-n���ҁ;��ܨ�q|����o`��a0�pV��Z����+��؇�q9��l�لc�L[;*�渴n�4r~x����0g+��^g3|�UD�f;��	9�%eG�U/=SՅ��!�����H)�3�Y��Z1�N`h�Pq���Ӊ~�Pv�g��~^�".W�Q�\�e��~Ä�}.Y5@KE.�0��2"m�ECE��_�_O�_�!�̓N���5��ڻ�䗬�:���X�U�:��l��]f���p$v�E���o�Nɨ,B~���?��;�Z���ׂ�ض���M's���;�>���x���y�\Z�4�>�n2A7P^@�0��yl<�gC+sM�0�Ű��U3@�|�C�]3�3�Pl͜�u��˲YP��);X����F�ϑr4��ᇓí�>i�?_?��t��fk���G \*_ȅ�P���vgy�+�I��J����+��l7ߞ�\UB6�����,��Q��S7�P7����h��8w2��S*t�]����|=uy탥�'2�
 ������$	?�Tw#y���RU��7���.�r��=K��-L(�S�Bg��n)1ַ@�����3�_Jt˗�N��&T������w�1��u���O�_�T҂��M��8�&������Q ���t�q���	�
���xTє���%��[�'_�/6��6{Y��]�s���m��j[RR�ݏ)������T��������[����ռe$*3D�'=X�>��D��)�Y� �I��+���|7#$ÙG>_}�]W+�N�D�[Q��z@A�Hw�������9��A�}y8P�y�1VsX����c#�*x����8�2f�t�?��^�~ɏ�/����(�2^ ����5�E��x�B�q�l�c0=z��~]P�\D��j9�Ol��w�Ƒ�>蛹B�`(����0,s��	XD�=�Z��hɜ�8ܷk�p@��}<=C6���v}�ď�_c3���1�50g"��#�#��*�٫6?f�}7�v��S��j�Cp��|Ɲ员K�穜�l2l���c�TnM	��#�u���jQ�uU�(J�q�#�O��]�a/���E5����՛����_1J���nm�/&���4-��x����&}����F����j��'�P���
<K��L ��/����u�&�|�N��W���ˊ��/F��Zx#�z�n��r��J!�c"��������aߊ�a��3�y&�`�R(9�@o'��?�qQ�nN��u��k y��������_t5ׅw��;���aK�a'�-���e���C�����y���e_v1}56+��S�Y���^qw4�t�|F�M�D*#dDP-�y�u9�J��aH���4���H������n�^N��Bnt��v�ShdD����~.���V�;�=�X��X��W��	�{�<f@���G��i��XO�^d�d�{L@'�� V�}��si�9K^
49r�`:.B����^N�e�B|)AOka��>ƕ�N`Xl�A�>�ߚQ�e�Q�=�t�>aVN�6�V�n=��fB�$~�xd2��!ӅXg7���O�ϲ�lrT�҆�ܒN�%��eEA#�#�,�J��}����t��7.�ܣ>�fb[��U- $\�5u͉�mEz#l�G��j<�%	+��
nK�^��j0#ϩb
i��o�r�l���07cI�����g�,��a�ᬩ�o�&f�FR/�/�<.5���i�F����@}���_�Q�̝AC�7l��D�FI!�mc�x@��/��j�#W��nq��UǺ� �cg����Ѕ͐�LQ��k���	���**~��౤|�!G"��I�����J:�lOs[$�t7�Z׊R,~:��F��O@��*��F}�`Q�x���c� ��@f5������ޟ��K��V��5"��l�f��&k� �+ȫZ��������u3v��g�%>�ܾ�].�Z�����mFژMi=+O�w��C��S��b�A�p�+�*�G���:TYȏj�gc��tH�͡��
�7���9`�y܅ �+��X	�:�!��,�*]��5k�f|�w'��:מ�C�����.��(U
.�"���1BBϪ�N�.SrG�}ٿ?��ۃC�w>&Ȑ���� aѫ*/|Z��a���H��g��x�}�˙��e_�=�3�Ck[����\&��r�} vm"����,'�v���uN6�j��Y��������[U��n#f�8�����	�
��'�?Ҽ*���Ɗ��NH�׶5P���ȶ������1�b��3ɢ�Z���ˋ)K*g�OhbC��G@H���1��C��R@`
�n�K`��&��#����,3�7p "�?�r�~����2>e�c�%t�y��
��dE�ږ9�ǎ�f�h>�{=:;q�Y�W&��i�g��\��6`,P�1J��m��v�
�൙80?L.��������T��}��~vD��3�L�.�;;D���j�1S��1�����&9�ɿМ$�k�S:��$����[���3[����9�����j���k�y:wF��+���{�.�� �Py>��m��r�oc2:9JbS���ڣi����.nN-�k��Ͱ)��2���Q� 4/�����x)��5�xŘj�BŲK�GM�7�t
�D`���Dpvc0'����)�����@���,���Ï'*�hI���DPz�X�P����1Q̞e�ELZ:U[�&���C�����e���25�_As�z���M|�rhwޔ��Tk�Z�r���K'9�ɎZw�挭}wW.�l�~�jD^�|lMA �}H !<��"��tŴ��s�#�+Ω /3os����m땺UöU9Q�T�{��9�-zi��l��$��^r[M$MG�!1g��=�L�;W�/Rvb_�U߮�9 8\Pt(��,����ej�e��6�PΌ�έ�.U�5&��ȑ�����qł�.���p�0䁆��sZ���c���ksW�1�aeS N,@���:��ɢ1����YP�<��F���[aNYi��86~�J^I�2ί��h�pC�g���')�ʓ�!(׻���~�7��i�foG+/��\?.G��7M�K�n��+|������f\Y��z��Gl��-,|��!Yn�7O�MRAgi����8{���y�-p�<'%��*�x_Q�m�Sa�����+��A�O���2��Ej�-CC��K�۳ZʐFb�CW�����rr�X�;2�{��Zl����ܷ��w�Bk�%��dzjM�Tץ_:R&��I~�{�����rɳ�V���W2��A�m��W��O�M���zj��k�6U�r��4޺�A�}hy�ͬ����3��0r����sgOW�"ţ�.��Ny���˒N)�i	0���w�Q��.�ig>�t(t^
����_�J��-O�@mEZPDdL�W�a�9 }G׸�K���d����>LqƐt��_�u"�ls��Ǐ�
�U�*Õ�Ov�k"틭��jSϴVf����mOm�2���w��.
�P�J�"����g��ͩ�,Px�;�Ua�G�<�a�k�?ҙ�tuE�d�ǂ5D�?J�&��*w�3(�{ˀp,e��k?)��3I<�@���ĩ�J���/������g�R��xM�0�o�ђ��U�Fi��-8��\8���4���������|$�11(ݷ̘V��=xʋ�e�+�^$,	��
��^	�!�.I�u�a��8�i6*�"���tP">���G"4J�̷���L�塢0?*��D���5q�y��������N��y��p!��MYLn���n��M��1%¯I\�D�g|�\�:��Y�eX��Ӄ�N�#��(PC�o��d��q�F��X�%�N����[��D$� �!��f3h���^�v�}}4�%Zp$Z
>4�t��#��F�����-Z{|���`�k]��(vO6�_,���o�ҽd��.j�3�n1����b}�7ך����ڶ�-�V��Q!LѶ0�KA��1T�z���
f'���D��j��7�pa���{`���1SǖP0�?�t�9811W�Ζ��ݻh6�	�OwV�v�S�<�$$G�ؔ��:�x��=Ȍ�N�2���4�;Lpo�U�6��g�5��{05�v�����V��</e9[�P�"���c���;�n��MN�L5��o�40.��!A�K�p>�0��߮����+|���Y];k�������QA^M���;�5��G&|��%�Ց��+��"�=[��,�E?%�DڔuaR~����ɣ�A�F��v�-��� %���3?-d�Al��BY��.V�`�A�o�Eϼ�H���ηk�j�T	 �h����C�T�������Rs>�/pI�m9��0}wSY��)0]��d�sl�h�؎��E[��M�`e������h��$�3���ܟ��ݐ����p���P�3R��a'��MLW\{Z���(D"��ҁ��e�m��\<U}8�E�-4R6��>��x^W���e�Z���
�P���c��\P���<�n�6,���Zox'��w�}���`���Wn���Ͽ�aư�I]R9�JFm>�,�
�:A\��
����ͬKO輹;��]�?j�ϔ@�g��a!޸ L��$���dķ�5�)��gD���b�0z�+��x;C��v��Q�~�Q�����$,�*��`� ����?��.Vя�v��s��[�	��y�~�x��b����FY-���|�,X6ḡ�.�;�?'5o��v�3����{��{�&��q����/Z���6=e/���2��F� ۨ&��4��0sz�YF'8/�*%Ǻ���n�]���b���؝��̘�R!ِ9��\a\�Ҋ_0��ٿL�*�F;dzI��i���k`D�B���(�p������Ix>��_��n^�a�U���֞@��H,��3��-�l��v}[����t�aO��M�Q7J�����Yuܻ��!�3��Flx���3/$�NR�. ���O�E�8KZo�1�=i}�.�z���ivd�ǋ��� ��>>]�C����ta��ūk�O��h66�/��
ViY)Z��nYT�ײ�_�:�����E�Ƕ�,�D���'��f��^����m��f;�}����������(F��<
_upK�g���;���E<�M��@G{@����P�V�����l~o�x'4�������sh[��3���R?"O��M�/L�����Z��'��Y�f��,'/6�r{�FX�k1hp+�u���/B����Ԏ�:�ӻ��)fH>�k�.8	�!�s�?������ �S�nē��:dW��!o�%��(EU�x�w�iۯ`�l�o��B�ᨫ�%	/�s� ��h^%򕭥:��˲�$m��
��p��U�dGH�����Zs���o��Ը��u�<o��hk>!����"��y\�R���x�o�l�v�ʱ�T��~����k�0s��k�X�u�(�椫���Q��=�];��/��
���@dDu���3eC'���F� ����H��x��@Ω0i-��l �dk��L�w�1�b���9CP�T@��I!�=`�W��R��y}���4�4`*��Ԛ��t�/�ڎ���/�e+�]�����*9�N�M)�����d1F(��|���6gi�mK��=�žƍ�ʣ:â�1P'q���d�9�����P��Z\�z��Oh�C%�`���:W�J�(�����*�J�/Q$b)���!��qQ>RD����׍�9��Ö��{�SҢ;�q̀�#�T^��Si�f��s^��A�<��$UU�~M����ؽ(Ab՗�Ʃ�͊K�Q�2��h�q���ل��Ivy�Uz�4Ahka~W���G7�&����X2��er{���db����ߐ�M�*ʤր�(G<�kެ&.u�3��ڪ勞�z���j��oA�����j�)�������wֿ�r	�5�$x����|m�[s����C����Ў�o=�E��x[״�5Ⱥ� ���o}�Ј����V{�&ϓ���[j��a��0H�"���O�R�ZS�H���H�m�bU�d�Eb�؂�`o2�D+�3��Q��~���}��[rT��a��r}I��*�T�{�k\3O�,Ίn'h4d�"F��ɟ��9>�ȅ�B�������ނ��7$�N?`�&�����+�i�W��P���!}���K蘈��xC�֙�X�.�6ߕ�>ڿd}QW�I�K9Sa��U,�7ke��}�Te�\rMqG;+g������>�b�Dn���㗡Y:H���~	XJg��}C-XK�wwQ<Fܴ��=�y��@髾(��C�T��R���t�,z �
�˲�-��)���}�=��~,L��&?��m*�B�W����X��0J�X������jG�{1�oF���sT��2�k{�*_��P�������K�Bu|b�,��B=N�� .V���������wF�<g�������~������@!��Ք�	�<��uP-�}1B��5 �K���/�k��a�[9H��72�>ǰ�EN|��6�w��l;11���o�n��xE��W��B�s��,���ֶv�]��,�����hZ��ߐ�ӿľ�:Ǎ����Ta����g&�C/;@u�uR����n�t�K/�3g�g�~��{������]Q�C��Q���ě�ݐ�fhM�2S�s�z`k?񼝍�D����˼C#c?�l�5l�ж �)bm�}�Z9��W�>��vSq|g=��ʯ鳔�z��@5�vso9�Þ�`�����w��0�v`M�yZ��d�AY̐���co�U?�[aٺQW��#6E�ĒGJ��/�~�������~M���Oz���Q��^�� M|�(>F����%!�.ύ��l��|y�X�"�ENX��"k��*��?m�Ȧ��V�)�Y���I��фF�*����$�S�����|<'^����C6��	�VK?����+d��I��;���p�*آ�x��.�z���I�f�x ���j`��'$v	�Pr���t�[�;�i��}��"�B��B��Z�0Wd'r��:?�L;��H��S�)�B��,��Z��JAf������q��jE{f�r���o}�R��>�
v
�w��(��Խe�o��y+�0F}�D��P���s�r;�%t�$�Orե���;�o���8��8��%���ye
nJ��Gz��-&�N����'�	���uu�����%C�0�n��y�o+d),r`(b�i�:�t��Ju�,��s���qC���z����OÜ+�j��E�.�R`�kP���~�jx@!��H�Ȯ�T�)�;Y�[�,�#�����╒H�Z�@/�Bɽ9a�C��4u�yIP�;W�����+Y�E���wV���E=̑��P��&��p9�'�����OZ����1�a022x�8��V�b")�}���8_E�"�}Hy����A�>���O~Q<�a`��e�Z5}rrZ��I�PR��>�/31�~��Ab�*��
�����Z�H	m;�|$���1ʘ�jp�jҼW�oR��ݭ����I�u ���DXd�n�T�ˡ,w�Q�ň�{�~� h��o�GĒB|s���7�j+qQ8�ک�TJ���BMA�yV�)�m?! Tş���l>���v3��,��/uz�ɕ��{�<�G�-_����δh �+�"h�����'}�K�g�OX�;��Qz�Hˊ%Z:��P�;F��6���Wo@�Q���ɵ�M;����h���rn	�a~b`Xtc�����E�#�siw5Y�A5c��|K��g��ߢ�r�ר��c�B�3Wu=��U���7M�RQ�;Ly".�^3&`���C�=��Y��|�mD��Fi1�'DEY�q��Egy�i�#��F��e��bYKy�|a�1�r�������٤��At|^Bw����?:=*�����I�.}�������&�Oz@�ȗ�V�p{ʫ۟	��z;���Oq�{�������,�6Q��)X>�I:�UH�w��Qw�Cdw6g�^&/NY+����ф�yS&�/&/t!s<��V��{-�!E.p"#5_3GGdUܚ��L{�B5���Dm�H8��9^�Fp��J�%�aX�WI�b��] �๓q@]>��=��g��b�v_W"=+o��0W�l�c�Rl� |c�pC.�Ut7,1�s�.9客 }��K1��L��s��ԭ�8w���RnW�b�����{B���w^�Ѵ��ݤ� ���A��^�74m��1Q
\-��]�ҞZ����nY����>�������ǇBpd$B�5ˊ��΋+m�op����?��BC���Ӊ�(��򾑼�ƴwj��\�D�r����eX�[�23<wiz"�0*Z�)�nzL�nH��������,�9pO���S�~C�|̸g"�P�QU���HFO�b��a�SS nAٝ?�"����I���������<��${>j�>�K�R�����'C"Y�Ϸ ��D`�ĩ���u�t�}���Psk���5�E	iɑx}y��~��t�f��y`� )�d���3Kq�ҁʿ%����~J2��V��ëa�Q���$�q<�2tR��4Y���@��)��(T
ǃm��HF�`vYe
{ Ԍ���N�����Kf$]���Ot�N��;��A~�lZ'��%�H�S����He�m[cye�dm�K"f�c�쿕K��_�X�5��\ߝ�	��`������s�K�/����n�
��(��]Z@���eΣ"����9a�R���G�U���/V0
%�^�|䌉��j��E4��5�"iwK��m<L^���L[��uUZup��2���1�0�
��lk��"�7��$Ҥ�� ��?�1�n֬�r�׀�`�H�E��-�@-�����C{�wt������߰6����������&�y�7PMoZ� 2�ϩ�R�{���G�}ee��=���:�nbxBE�:�Mq�e����$|��y�۠���O4]��SK���u͜��N�Q�͂�	^>�C��`;��3�g'wy�_��Ռ
�!�(�ϋ��耿K�F�X(��Y��ߡWw�{���։E��Y��˧7�`�/3���WkZ�����:[$��q5/9b���y<��7���w���t��!1'm�4Os9�o�x�G������8��{D���k��i�AK�:tk@ƥWbx���E<����γ��T�:��2\N��J�r@�RB���K��R���2L�}��N����|9��}B��|Yd�I�O�A�
=!����8��yz3��\�Ѓp&Y�M����+����ø~�d�B���5��?6xg$j�o�w����;7q1�r� �����y��w<UX#��Ì�0{��fN�G}F{�[0+�K
�ٻ0��S
�����z�I�2�\�o�bhA�2�>$5y��Ջ�����z��0GP��X�v:�􃞥x�5��L��[I��՜�+�	�H���+G�٥K�L�H��D����$�z���S�^����`���9}���71<��1⽪���$�d`��
[�j�hY^GB��#��T
�93�2�l�(�H�#�Ѳ�	�f2p̮��I�A�}F��F,b8x��	��,1L{�~I��j��Զ���5��j��N��[//6',��3VӢ�C�8�v6J���;�;�):)�᎑���`R鑺Ip��f���Ms�)�y]JhVC�T�����Q�����lV2��ax2�+<��j���Q8�������.�Y";B@]a_�D�k -:xt�e��A��=;:�9�/�Y����)���o'o�ۂ1�'�Ӧ?&j��r�9{�q�N�o`�ʂ�H֋F���g#�C�{�L�|��k�O��eb�*�.H>`[��hx��;�4�t��bBDf�F�����2ћ�F�oX��:�޴��>[��w��< ��b7c16��ДW"[F#�x������t˽�q���>�V��z;���LX�&P/���w-#�
��?���T�l��*���k�gxW5x��{<q�w+���:�άyX�>���30��@��@��r��݊�7�zf��h?x�Y+�
)�!:���Pΰ�F���
�z�#��b���_�6o�	�)�������>J��XM�3�LA	�jH�b�^�EYC�9�rI�O�ƌsd+�ŇmeK�.��?
O�i&���)T�^����~śυO�[V�d�qG��}�u��H�C�^��!�G∐�^����|�R�5u�v�
��f�e7GR!�|B���Φ+>�.DbT_��h�,�;^�AM'4D�1q�zix�3S�:R}]Q���ן?LH3��;*;��K��q�0���C>�G��2�Amf�Y�-Bsd��B�m���z�b�:��v��|z%sP|c��F��͜X������>��^�e[4r�Ub8��#C�r9�G�s����Pg&�E����a��]��J}gŞ�ׇ�6�]8�Oߎ|�֕[�c=R�@�֠h;�E�6ﯟx�k��F�/D�[	j} F�kԠ8�i�R��V�y��7���5���������[�A��Y,��gg��aب`)@e�A��w��BZ4�$_�s�k��B�sH&|�#T��m�zu���A<��J�0�Ph�&�է5��QD:���R!<��ؕ��o.	�F�e^�7wb��m�d&�SQ�JCm�{��{��Ì)��n[�;�����;:����Ǫ�L��L�K��;�|e�䏅y@f�o����K����{�\�L�������GCe#�ҍ�� UMhzam�=o�H5n �E�G��e�w�$�Y�<�gG�:r�X�,�y�w�k#�|�W�s����#N><���f8���ab�6V��`F+K+HV��<^L�j�E��VO�y.Ƣrw�&���]<�a �����ՙ�+��r~��s���gi,s+	�	�Dַ�fj�iVŋi�
+<P�s׍$V�ovC�"���W�w��O�%W��5/bCI�W�F�å�-�Aݦ9$�t�܅7wd+j������	�D�6Q9���K��^��B�еZn�I�;� m�)ۂ�\�ŭ�c���%9��؊<S ��a a����q|��a��/��!7�p��4-�q���H;�φ�އ%c;9BPaG/F�J�]��!�<�,�5���I�� c"3B����spw� �1	�� ����$��\OW�-�
���{��Q�/��0���|FlB�lp+�qyߓ�aB��6���#� Y�:hͪ�+�j�k���U��8���!�7���6=|���
Z�����r#"5n�eo����=�6��>�b��\�n��@n݄�f�����s��	_�.2��V��y����O����[==.���@�N��������������Nl�8*t'��m�'�����ϛ��C�Y=�ݶ����7y;�W�-2reaqV�������S�ʩC���0q"��W5}m�hHf��ԑNu�	������Օ���RXޤ�����/���mJ]w^�;�з��L?y��ۙV/��H���-�S�_l�mf����$v;��@���+��2�i�I�+, �9@��J��U� h2>��T�� �c#���dͰ_Y�1�L�m�|up�mD�"y�,���$JW>T����:�v�me��go}09ɴ�r�>���л.��͚b��Gb��[U�n�A"�!����<��L��L&>�����p�6��;�3Ҁ��+6ol�n�ROZ,���̅�9N���%ҋ#)š'��x[�i�;wu]�@L]'�i���jp��!���κd^�<��T����Nڽ����E�ۏ����.Z�}=�ʕ��|�$E��'}C
.��99��m>�5�V>���g�/�v�,ؕ:��ڬy�]@��n‥��	< �]�'[rHi5[�a�ΘÁ����SL/j|2D���a�qo�%��1} ׼Y�Z��w�F�|�a�qS/h�������N�`�F@I��Fz�9l(���n��{o�&BG�'Q�0�6FY�V@p�LhL׈�@������L�`��C���%
;�p<��7j�V���?G&���6_�>���ED#P�@a%&1�=�����uj�{r�lkLk~~l~:���1������?�`���_p�6�.@��c��z��y�rU�?�lc!�ҷ=�B|y��̢�)�AԐ0��9���x��J?�<~+��A̳z���c�f �����Z6�W���?�<&�|�-��`)WT�j8)��r|�6qS z����l/��Fd�ax|X~cw����v�Ϯ�(*k�Ҋ�"�#jGc^�+���v����I�л�4��4r&ݫI`�X=���γǘ���G�Z�� �5��+#�Jn[�K��U�ƈ$�U ��2B�:Ym�^���q���yzG&�*���U/=��,T�D܄�j�H�S�Na8�"�
(j�C��)k��,pK�eC:�KD	X��}�����k�X7��=":���s^���/���@�Í������,ދm�
�k6���|Ķo����������1�q��;8bc�,M��8�J��+�o :�/�@v}�����y[d��Kf�Ja��<�@��be����mc�e���XT�m���#����õZ����ȕz7=[�]���D����$�D��)���zf��d"󾴮}�1�6�E��hr��̟�����X�Dy3n�!,���-�-z}�l/�s��z-���fp?l6
Sx�-��U��I$׽�ԝZ�0����.����^3��� �c����q泱�Y���cX���m3$�}�j��2q�l��9;����p%�+R.�%`nC���ho�	]Ijʞ����^���Zf��2�"������wI̕�I�`���>�N�Y�=��%�t4j}��/tX��c=�q�A�ľ�ī#��U�,X'H��IQl_�f�2r��� j^����sha��26;�6������>�YtNٗ��G�Ç�;5^-EC�p�K(L�������"Tz�E�?�Z��53U?��K9`�$��c�;��l�pF8��_��ey�*��u�2��:�����WX
~M�'�G>�Z��r�!3�6����=�����I�vNp#�����N��6������-�P	W
��_?��2�	os��]g�_��n��ͨ��2|p*��N�l�����Q;�x{�ݜ@~�����Ms�.���Y;�smKE��u�=˿�0Ҧ7����VB7Mx�L��_����D'�"���+Y���f'z��NEj6j.����^�{�/�G[Buk��ؤ�7��w�A��lq��^H<�Lod�SP��^�o7�d�W�r�P���hfκ��E�ރN3�h�� �f��Z����,�P��{��!bӺ��}f8�6o�1W �K�ɔ�ʤs��{�6s�H���\������\s���)G#I�`��o�y��ߩ��߰4���5s% �Ȳ��F"���a��i^;��Ů�W�(*お1��O�l�ê�9���寖?����m����R���Q�������Z�M��r]���G��������w�Rn����R�L��{\�r�$N;}� ���[t��"(��g�6y����ҋ�4�n���O#�tκ����jG�p^�Ü6��M̭���'̫~#f�p�Qd�t��8m�)���j���|��Zb�w�ʱ+�!��T�P�뚑8 �)���3��@�B�3Eȡo�P���0�q��Y�촷�8ٙ���z�.d�ef��D��� ���,V�>������>E��� �&T;у	�&y���zZ��p�"�A� 2�)�]Oab���B[y���#+"��c���{�Q�7[RB�N�1��m��B,����k7V��E���ȝ4S���_V��B���D0��cxK���%M< ��(�v�`�����r> SP��w�Y^�:��VC�1z[�#���zu�����u�><�A�c]��y}�Ü3�>h�?��Ph����Oi�,Jv���q�}��k6j����a	�؛k|�#�/`���3��	�s�XYLs�b�2����l�;�o��pn#�<-S�Y�L5E�go�T�!d��$�����S/F#���!��Η?��\�<�T���,-qI�įB}�������9�����G��䄧t�: B�m׷��R����9l0��k�.�E�S��O:� �L2Q:��z�6���fz6H"�#���h �wku�W�嗬�y��gV+��h�31�=�cju��ə�5�����_-��\�G� ��,�n��r�����Ԁ�m��t�����0��X�v�zEp�oO���V�H�v���f���4Q�^�CZ$<xIa���3� �8�-��6L���.Q�������ntb�.ձ���KV�j�~N��a5)����3�3<T��m��̌���ܤ�^�� ���>�\�܇�OS�*��C�Q��{�a�f�wY��#m�ܾ�����'� ¦'�*hf����w�J��2}��u9)5�q&��N��om�¥��i�T�90'�/�X�iCuʚ�a�B�(,8��{������� ���YxXEL=�My�Z+�Đ�]� ��I)���#��m������mXn4K�Gi	�3����Y7�C~�J�k5�s���dpYM�I���d>��Y*�F�"i��{����:��4{EI;{pUyQ�_<<�[�A� 2Kof����/?G�;��%%&<�A�Zx���(|����Q��<�f���帨�O�/�LX4cV�p���Q	�h�a�qL�����<�7��\��Cdp��ޗ�D���֔r����Ek���ꖃ��2�g��v��Y����|� �D�@��FO�5�OG7m
#�V���@�����~FGgkO:h�����Y� ���3��>/z�J��DNT'��������f�,#1����l'��=5gF߬��\:N����`�d�l��&��g�c��KQ쬥��v�A
N{�b�M�� �a՟�4o��gLx�l;�A�	U,'��9A"�+V�� _��Y���h���j��+���1ƺP�Ieq�n��
���	�H�"2qg��Yʀn9(eëñ�T���wr�q$t�C5)j�s�7����׼?>���<m��~B�,/�V��u[�we��|�aGˆt�e����
������$���������n�����ň$��'d�]��	�U~S��X|��a�)���� ��U�ſ8���-$py�;�'�m]�*9c����A��6�S��;S�d�H̜�B[QҹH܄?}[�!\�R%���Jx����C�X��^�)���|Mp6�����<�i��`#B�^#��rĥX�`���9%�\n۩�P��W	+֓��u{�,o��˾3�p���x�S�fBY�G�G"-%Y��Д_�� nG����[�@։
�0� O��*�;��Jj�0�ԭ+*K����H
*V�Q0ܙ.��hD.o�,^�=����"�$L^[�z)�#�tTG�k���4�pIy�,��#�3�u~��-K��3'gE�HI=�M]6���$�vO�č�4N�ة�t79���f�fJĂ�%�0���2cL������Q���.�d���׺��&�h(&"	�l����4�)�"V�୻	�n8�6�t��Y?_gK��#R�DyF�"��P�v�o�0���̽��Q|�jڼ��c�Q{(����8��Y���m�r���`* T��H��9��n��U[��֨�G4 1��LW�����}F#3��ˡ*; �L��d���yٜ����7ZTH�s�a��6s�,����SQ���j�����k�X��a����h�\�)K�w�]yh��*�3��菖����jZ�=��rs�B��(�(�^Ҩ����a�mp�Y�XU%�0��-�6�y0��%Al.][���r�Hs,�Ӵ�&+��;�^�x:$�0��Qg_�ː���6-�A ���P�nA�Խ�/��|�	�����ӌI��U�V=��[���:A���g�k7���PZ�.���2	��n?�she��g��ܣ�H�H�P�榄h�krV���N��M���Ѯ�5���c��e<pֺ���%��M��tc�ٶ�w�/]�y��D�������7�;=�NS��� ��\����p&R�����Nd��!	�$*���J�Fw��?Pg�^���p@�$��6�RU$y�\�LR�"h�B�E�7�Q7jZ���Շ�[��=MeD�*8�^{��<� N����%�l�n�qOA��78�����u����X�����}�Q�Ve��)K�Zu'o������@��m6��v�]��%�������VA���cƁڕ'�f�_0��N�������$�S��Qn��F�� ����+Yλ�[j�Hҩ�#��Dpy�t����>�u^�(�B>��* �}��/�s6L1�Ȅ;27wD�_p����ˀt��Ƣ>W�/����c�v�s�u%����E1��D>-I۞�C�{�`hJ@�X��ܼB�'2��|�YS��9a�.6C��W�BSi�!���΂'l��Q�je��N�"��+����S쩽�Ǻ0���>i�H��b>�V�$�%�Q��\Ya�6nd�o��0���<N����󷴏T�����e�E�M�j������n���TXn ʜ���U��C$](�ۈӫ~��Q�E\$9V�&�w`��?sE5�v$�r.��?��Y�����,Ƹ���"��I���W�+:*2T�
�i�̖�Ñ����G���V�)cW�З�x~Hic�W����Хߤ)rā�"]��Tl>
Q�� �h��0�i��l6�Й�z+�+g�ͅ�r[)z����N���� enY_�K�ʒ��{\l 6_��Ҹ��1q��+)jLh7�u̯�]uDM�^�M�v�hhtn!,0-Q��Z�3�¨Q�KNz�q�o��y�����@oS�}M�&a�ח���Q]�<�PanְJ����9�}��1ǋd�J��}��n�]=.p�P���	4k����2=x��M�k���Q��{�0&H��mvEYm'��1}�J<t�e�6��ʁ6K".=� 詡�d�6�=�3�=�ggtr��ȗ�O>ݫkg8�Kd����9[_�+������r��[��>� <���y�2�-�z��۪�TZ�(9���M�f�ÎP�l�YOM�.��{���m,f���z��4Yu��7)dx*%K�x��{&��:��n��^�����}��G�gO��Şam���UG^Qԅ^��j��(��p�̈́(�H ����\�[��gj�tF��
[z'p��h�LɎ�\�{.j�x,AdU�[Lo�4��ZZ:c�Э����T'�G���i����a ��w\}�%��4z����L�ʔ�2��L 
/ڗ #*�6`9� ���f���)��Qi�i��'O?3��>H����i�Y�I�V��K�ղ�G�_)c�e��WG^��&���׮�Boi��]�Ci�Xg|4�J���eLiαb�8����F6;�W��uz_6�H�-f~�e��#9NԋT͊bt�9����3� P�Ѵ7����@��Y$-y�����P�\w@��X6�u�#�H��Bm�k)z���vR+��h-%]֦4wN'�[�D��ʁ�G|Π���tQ]�:���@��*W-���S@S�����cB�u��(�	�a��OP�`F/�x���+]����\�> E��17]~˒��O�Z/�pĞ�<�
p�\��v���#���P��M�/s�#������0�����w�J��|�c��s�*5y���4�E�ϜxR�8o[Q <�Ģ��~D�����p��D*,�5 /�R{
��i����r��~x;~��M��ϏT�'2��(��.AiQL�l���y�%':⡿u��[&#��1��p���D����v��ZԙJZe+��F�1�~�x,#8�<��h�6��v�s�ZE�(��d��)��:��;8ا��->�U\�Ҽe�:S�N������}$d�����6o��������,��O<?��r`����2􂹞,He����cYn0�k�fa9x�M���>�Z����;�o���+�k�]�	��0��0�u��ZO�-��^"K-S_�h�򨞌�����1���§)0�M'bok|o0�v�22)L�]�1����k_.�)��D_��m=�BVv;����BV�K���:��/�N�(5��fZ�CN�w�%����䨇��Yy�Oua������?�ó3��|/O^��[-P!V�\�>��>Wjboc��Q"�l�1B�`[)�AL��_7�F�!:���\"AU�B�F�_��O�X�z��A�2��.T7[tv�������V�czY�3U/��4"v�AEͣ�*V���EYW�E�+��'W�����w�M>�!��y��"8x,���^�@��k��u�_�{u�zW�Y}����:-��3�!��)�	�!Wc�~�[2�[����pB��8YA�� ~�^ ��{4_�س�o����`��Q��C�'�%��� �'���h-�fgl��|{�A�4\e9#����b�Y�m�m�W�',mUx��e�'�C�&Y��x�z�����=�^�Ǆ4kZf���n�0h-xi%��VC�}��cx�v��يk�J�q���F 0p.g�m���ч��s���B�O���;W~bc5 Y�6�J�u���R" �N�D��qa?m�f@$�[)3�o�[��#8��Ϛ�nՉ�I�l�GS�����D3}Ǫ!�\�>�O��e��*��%�ɛ��Gh�;KqN�譥ߒݕZ�w��:��k���Vzo�8oc/tQ��HZ5����S)��a��imE���p�:��ӄY��uͧP���Z�t?!��J��/	65�YW�"�i�(��!+�L��u�PQ��`P/�){���&���{5��K��f��[SL�e�MAҀ5��۩��,C��׉�k��}��jO��}�5f�|�I�����v�W�0M�KZ$�l��`�J�m�� q�w�T�[FW����]�vwp-Z�'�ns17�	��\��T����-�;�yȲEU�j�/r��侤����ME�@UG֪V��p���ND����kp��MoG�o��3*�u)�i���1�B�f-�Ҥ��^�wV��5��]�=�~[j���y�<�o6�d)�_&Oa#Ce�*�;����>���CX;4j��ߞa��<v�x�a�c�]��"����/ǥ�ү'W��y��M�(��3e��6XBD/�M�(~�X�6���M�ֳe�ؼ1S鵡�_�3g�nrZdX��c�ݬY�n�&����0;��㤻�7�M]�i�+��gat���P��T�۬�t6G�1&�].����wS��C����X�X�PG��
��)'*�=ݲ	S����̈́��)�M\���{�7@0Gp�-:(������oHFI��~�2���!tq��fMf���)����\7��_����S�d��~�	�q1yX+���a����e��A�@E�����4�
��`�K�3��㞍�IJ����<��7.�,�+��T�V�-�DRX1e6�C*�t�"�LZ�~�4>s=נ�0��:����L�L��l9��93:�����!���AuK���9rY�1�$lt�B��o�g%�|��69�+�ʁՋ�-Y��	~h ѨK�upT�I���f��ܓ��%sR��2�F��O֡l��ĕ�F��h)�Z`��d�.T_�%��Sn�����ӽ��@�Gr�}�\�����ߜ�-o��p�n�8��I���b��;��t=F�ޜ��1�8�I�,!���"�yl:�2M��^�l�������[E?�/���5��|���`߂a��tu�^{�vprtpq���|�dˇ�n������xM]�
���փ?����K�L�^�&2r�y�K�u���u��&x����5�bV�^(�9��0�J�*��|c'��E�=k��:IR���@�u�B(oRF:+�q�p�)c�>���K���4[�e�ק	]# �SI���2��J����0�J'~�eb҈����it�g�{�:śyQ�Ǣ�����"6�������Awd��'4�'ZY1�����K����֝��X������i ��J��A��a�v��t��Vw��jP��B��|S��ݒ���;��W�xX%�'���B�53���J�����{���Z���]��-EA�/�����$��は�󉓀�H��ڸE���u��K���K���?���h�vKgA�*�9�l� 6�0�0~s�ב�z�`�%�°������@3��L�����$P9�I}sS����\�o0GKP�5\�`�;2�z/k�3O�'Ɏ(��~�?q���z���7�M��?q�Z3~�e ��1�[!0B�����dv!r��Ğ�e0�a"\i�8�����h�`c$�	���C�ѵ���m$��\n��
~��mN�׃�*F���u�[�mN�-<,�[��ZrIa ��͎�Ϻ�[0
����>��tUb�X���NHy�^�I�Wkj�>/�nF�fie΍�{}��l�@�0@D��_xz�&�#������]9�`bt5��;J�������@���e��X�3
�̳��%��o��Ű|dc����Y������yg}`�� ���k�	B��X+
s�p��e��px�w>քy����k諅�K^�&��9�_�>M���P�:*6!9�x���C����س�P 2�%;‌l(��	�3�l0B� C�f �Y16�y��o��I�N?'�
�l����J6�)�V����A�Z��8D�'eo3�@�ǘ��XD�0�&xH>��)4Y ����JN��L�ۯ,vd�C�2�ru�L�41����m.��#���׳�ߌ,h��!!�'�1#��`O�5����L0���3�1Ih'@��T"��n�/�zD�����l�L��)Ğ=k[0;�����^�'���1�nɊ�l�	s%xtk�}X��J�j��\�)���Yk�|~�j�ס�\��qb�=!'2��~�Z �E��0����f��m\��/j@Z��*��ߠ���!��L^-��`P�}��K�� _���q+���i����<����q�V�U�D�uriW���~L�ۺ��$��^!��:�X�� E�������}R&�~�X�K���	n.e��u="dZ�O���:�R�A��ë�C�/��Q�A�"K����UPe�@E-ȇ������g�6]��-�&S�sJ��x�:�^8ߘ��E0�H��˨D��b�Y���ѳ�p�������o�Oj��ʐF���я:��n��#=��h�h�O!���o���?F�.Y#���-�#;��s���HQ�b'yEn�I�nC�..K��?�=m��>f�[lù0[�O�ވJ�"Ɯ;��KŻ���5N<����1��3
îM�����  >G."�Ψ:ݾ�JK�(��U�Kxbb����h�k�&1���J�e�)�Ŧ�D�~-`��u�6�Ҟ�IFX�N�� `�?4�tZ��z���˲M���|qa�������m)J��฽�Gh�" ��F�x��E�f�c��h/�h^�<�w�~R�]�.!��Le�&/��U�V�7���a�j�%���C�ci-�pO���>{1]��`�>��e�Z� �U�5Y{5h�*�a�F�B�W���&���Գɣ��k��ʏً�1̹�F��u��v֫ʀ��� �j_K>����:F��)�ts�w%p`��7�.a^h_ݤ	$%���]4r�`�wdm/�6����:���~g˿�����M>�ˌ�U��<-"��Y*�nmO�ʹV�[�� ��rdޖ���t}�V�n`�@Ԧ�Q�F{�,3c/�!х6��NH��a�U���8tK����oË��&�uǘg�ItI�8�O/c��-��N��8�)w���R�S�"it�&5SyQ���m��O�E��v��Z>nX��Ea�*-!-�G�����r����y�r��Q�'G������<����>D�oQa	�1�����jr1�QM�W�p��u�������>�V����'�&�y��#Lq	&� jz�� �^�"�������3�V��>�1M]�j�Q�����[�o�j-�$�|�#>���u�����ʑ��$G���)I919FUH��D}m�[����2�����CGk��j��4 FP;�9*����}K�Т�!Pn�n�!�3u��Ɍ\�F��em ;�Z\����B9AD�����n�j���X5��վWw���m���-�t��35�*Z����3��Df�2wv�H`��~���f[,���N�E:��^�����7�Γ}��:��04����V�6tX[��p��}����sU���r�T���B	!��k�:d�q/r�=J� T�*%��ҋĝq��#ϡ��>���@y�6�NY������O��K:�t��m���:Z����w�;ű6S.1����(�6R�^�Vh���h�^4��1�ׄ[��� )J�M��H����*V_Yy�
pCzX�_�a��7��~M��Ds�
�z���ͭҟ+n�������$1lb�^4n��q՝�����@�׍�lg/'�<3�����Μk�݃Ĉ�`� ����~pp-|����P5Do���X��^�TkkOq�/�����1-zl��\�H��`��;r�BP��@D����-e��*(���&����yo4@x�C�
�E�0�|����J��M�<FR�}l?{�՘�(,k���p�,�P�ǫ�ob�
��#�K�C�0�9�#&g�_1�
䩅s��|���C�F�b�ңo�γΙ¡PW��t�pO�p[�Fڣb�Y{�a�z������{ נ2/��Ds*��;:m]�t��q���_O�_t0b�c�ᓼ$����i�F�D-�|���,U���"3�F%F}��U&��YI�H�=�!�u3�%�_Ն�uH�oЎ;� >m�$k���l�5u%���;4�?AR��>��]�يs/�so�4�A~�G�gF3\�]~�&:hܪ7+�%��?􏹔7�`1�wSCC�7�o=↞��{�&��k�3Q4Ê]��2�嫠yj�y����@�7J���%%=]}8J���
B��x_�^<�K�s�$[D�\��3;E<ϡ���jq����Hߛ����Y�Cxs�aǸ
����	t���v>�m���|��i���Ҁ_��m��@H���g��!�*�����]L<�TzP�uLZk&�O��-�&����8�1s8h�7~L��Wc�~<��wq�G�ϻ
E�A�},�!�"����sA�D��2�T�H���'l������9*Vį��<����z`Nr�G��I�?6�?ت��|zp���?��G����螱g�Æt���i�/�A�yY�2Tii�>SkY�g��κ���^���Uv]�'.�X��a�*�G�6��b~G��P\�|0�����wvgގIC�s�
�E^5mͱ�Q�Ƭv8��.�����IZ��Fn�>�F,��K&�R�1I����d��$JF�ŗ��h�8���[�lm6"s&�YR�Z�뮍��%�-�莟��ʮ	-��Z!�A�o.�9s����t@�R�2�m����'=IEGK	9��C5��A���J�?x��A�����w�siF�U��j��s_\��4�e���bk ݟf�v)ķ�@hǨ�9�s�@M�������e���An���<������M�$v�����@�Ҟa����嫄>�i'����:�}Or�@0H/��y���p%-X�����؉ ��C�s38J'-����F��kG�� /8��'��]��͆�{�G ����n�:�ʟ��2-��[�̵�M�Xŝxy:l���y\Ւ�tg��k ��V�V����}���!�&��PL���>!;�#%��rh�-CLUzYsQ(���awB2�A��?�EIAD�ǇQf��M1@3��E�����D"\��j�J�5�T��C?h��'qQ�Ti��Q���]�v�35�H�Dܚk���$�A݂2��؂��ְF�kS�f�y�;m����k��4pO�HnO�:�/�Tͤz��Gl߄�=F��j�����<�1�@�;)qǕ����q��^�_ �	N�sZ%*�.����R��T�|tP� =�X��ő�U�&r���α;p\�áp�>ҏ������������F;���-il�(��L3�>�d�����;�hYT�6�1$z�4c$�Rt�U&��X���,� ��K)6ڌ5+���k���Tk=�t�j|�s���3,����C��`�ḽ��~���/�"����_Ib[Qv�}�[����9	&����h���X���{��~Q&z�/���4�e1�4!�&!m1��N|ڭO�[Jbˉ1G����S" �>���\ջ�4�ԁh���g�X��KR�@`�+J�5��ӝ��<�d�������a@�o���f>�X����5TF{�ӏ��l"@N`YiH����o�vU0d�[#(�����+�j���&����dHD�y��|偦�,��}��R����o�T|;Av=�N���F��:ų0�S;�t���@���+5���)^$v�㜋x)�@ry���}N�#��|@Б��Q
X�,���]o{@�z�\��N�Q��4�����WX���b
�(�dH�@���!��K����}%\q�r&{P��U;��;;|l�~i�?�ح����l�n d�PD�0R������y�Vy-�9��5
~l�8�9�A_Q�e�]��/w1!�E�M��N�%TfV���Y��i���`pe	1�](<���P�r���QW���9��)
��?*��(�Xͤ�(�X�!��~~vv����8���������?6��CsZC�Ax�d�W���,��XS{���(�8����E7J��P�A]�m����J�$y�
r�D�ְ�Yr��ƞ�K�e՛�1����K5��Z�����Կ)w��6�~��a��g	�ِj����׸0��d�uL��=b�m5<�77Ol�{ƫ/D(�h��揭���Ž��׍��M;�[gפ�}��p�w.[`B��<g�(;b6�,�#�,�>�v�9�*�l�%��4��gL++q��f��#LRCI���7�g�t�*y
�q�fv�JA�� "hNQ%��Y�u]�#��2|Y�|�!������x��B��� ��95F��(�D�P��ߑ5���j�`L5�R�Q�+C��j�ޢ\�m�	�ށ>�nqs��mt���c��#� xH(�İ��M���	�yY�}�3J�iS�5��d,?��X����O���d�������������R�i���ߪS�a0��H$o0�`���b�1�f��a��v�U�G��
~	���k��b%�3m M~�VD�1
쭻���pP�惡C�06'��[H��@�S��ğ�&��c�W�GN`G�a\�(���ɔ"{���m;�/B>ދ��/���1n�sH��-#�\�rP.�u����gZ�w�x8��p;W>�sO�aӏ�G����o��L�ϊ����Ö�+ba%���t��{�RN9?]a�a܌��N�Yy��Z�>�����Gav��veS�#]-�%�VO�m&��(O��a�>��[����b��a0`�S�r�c9Ar0��7���_ �����%[:BT�����>���R_�}(�˿C�g���o*��0,2�A�쵩��O�R@u��V��K��B2�m�#��X������e����P�������7`
�tsf"�ۼ����,��`
������Ͻd���_�R�s����a��D�� }�z&��sWA���oZ�o�W>.�ƾ�|(m b�[[���4�Ql+��ѠV"�1�.I�&��m��54��FDy��V����:ȹ�+bZX�������֥�u:]���S��K[��\;6��"�{ vQ(�t��8�F�4Xt!�;(*����b><|>k݁㳜� �!7��˹T4v�l=O4 I� �B����n�BD�[����j��a�V� �Iϝ�߿�i��n�q4�cB&�W%��ƚ��np-X�vGT���.R���=F�pM��؎.��o�3R�3����K6�f�Ƀ�������k��#��x��o<��	n)Ҷ3�Ι��	t���ue��g:b@^���.X�z/�����Ǆ���Z��:e�������$�<�/ĦD3�d)D�U�#l��j�O�O�p�P��}�XoWRs�� �I�b�����;(�:q��ye�-�ʵq^���q���v��`��0�� ���y{}(�a�T����bV��3�A�M9:p�j�,��ƛ�=����_�:Wv^�7O.��l��Z���W�{œ�J�Ň�����f9��X��Y�t�d���"iuL��)rӃ����J�P�����`���DIF��1�j�Lt�����bx3��\�@��D�A�ᨕ6���C���[�<��<�:�(�{�۔���cB���i��Q�qz�ֱU�S	�?m���8q��*���q{�J���h�A?�?u����+x��6�kƶ�h9G8m.hļQ|��'JO�H�:/����J�	$�����ǡ�����P�ۜ�m��+��5�#.�e0�~UQ�ݲ�h��Y�0#��Aa�g��{!?A8ԧy�Yyb&�S_�2(*��T.�~XC6���7z+樑E�O����c����~tyj�u�e��7�͸�����67U.d�W�un�.��4O�R�y����[�����N�҈��r����xo��I���d�}Ƌ����Gw�Ŕ:�R�#�E"Dƪ�8C�����5e}I�"a� �bx䦌vfG)������ǧ貈+�ߨb��Q��(���v��R?c�u}��c�"�y.�x���kvP��߀����&�nśU�𛧠ѭ�%c������6v�*# "���>/�q<����X�]��Xh�s��n��Ĳ��}�p�^�;A�١��5dg�Z>-�h�QY�)��!��#�漚h�@Lm&.���X�ܝ��
<��1T_��	�u�����ɉG��y`k���y�{/l�W���� �G6eN�)_C
��#�-�?��,z����
�6{�����}w�֩��wűH̀�=�ӑ�hX�E�'*΍+�Uh`,3�KeX� ��:�A9&��\6`Kf�FJ�`�U�?q�ɩ>�3���+�S�s|k�Z/[�h��N�]�r��Z����!���zt�ixK<��n#eM�C�Ju��;�]��qeF��"B6C�+�d��%��+;�" �Y�v��˦��] ���\,�َ�px�+�C@�ݤ�=� �l
����n]\�%���+բ�#\L?_����ɍR��O����{������Z	�g��$<��#dƊ�,ROn����91X&bF�U����jsx���(�z+�f�ј�����w�5�5ƿ���sR�~����}HVs�.��b�z:��;5�'��KN�o鴙'ɞ��g�Y�M���.��/"'�A����ǘ3IcR3X��:�C�D~�:�������4kfj#��_�B�@�|x_(��o�s�`�N6A���w8'u5+^D$���e�����jXmȍN�qQ�f���.��>9��g�����bk��s�MAV)��h�藘�/����֙�]_��9��p��TQ�# �_�S37g��<�&�U7[���ւ(�Z�ݬekȀ і�:]L�7{�ެ\����S�s�Y���$����+X3�E�LQ���ߧ��2��e.P��=�����#����;�e����L�(p��55�?��/C����tTu�������E��)��_�۩\�Ϛ`�:,�x��/E2}c�N��:L��c��c��2�Ǘh�'�2y
}�:Z(e�����:�|�cBYܻqNa�M$��}c~R�P�uE[q�ۊ��.�� ?��[<w��X�֑�DK�/�Íg�Q�9�[;5�D����ĉ&�{t�Ѥ�T��.��f��-���d���( �f$�'��\^˭�����oA��k[��T��r�٣�cz�����T4:�C~;���YZ�c�l�GՌ���[���ET���b0C7^S��nSϯ��~q��H��ؿߑ�J�cM�r^���u�δ��	�`)�iЩ�S0��F����o��-(ؔ^�g�H�<JOoƦ~R@�X|`�J�
���,� >H�x*T}l��Y�%Ȟ�J��y8J�H���a1�JN��;\����퇶����l��\��VN�]�2!�A��PN>�!2)/�'�#lBL60dc�$Ӧd���C����J)K���)w�����Haݷc�9A�>0O��+�ogW�s���7ȱt�F��»��<�:�����0o'�5�n���7Hi�xMcU����KT[�� �P��Gꄹj]�����?v�N�����Ta�<|.�S�vE�X39i�F-�1@��C܈R���l������9���PͼAv��C��;�0�-�b�٥� ��|�HE<��F"O~���-����|{7e9ʇ�}�&K?���-̂X{����6��RiUq�۱��ƛ���E 1�*�+�ְ~Ǉ�կX�6)��?��l2����7{uӗ�U(�ۅ�DY����{�U�ޠ)t�+��y�m�������ؾH�����tU�a�9��=������m�� lF���l<�1nZ�w�f�P�o����#)$�hu��韩Lxf�i={̉�\��Z���W��B���J*�}.E2���$�G�D�I���AD|���:i�͆�S��Ԝ�1�[y�ذ�$N��L7��H��C�{��8õ�~�����5�������L�A>���*%l���Zl[d��n%�ɩ�rl�kv����g6�(`C��E=Z��5�*��D	l.��7���<]�8'��Q�t�
;E6�9��D�]'z�ޟ�!$��7�W�@܉��C�����݊I�90������[V����;w�i�d��k��� ��"��"�ϳ�('��eFp�Y%���P�%��Ckh+6���E�A9�O�7�Yੱ�v/�%PT5�k�Ý�ZS;D�����s?��\�и��a=�kii �x��U��';G���6~�>���<�s�<bdڊf �V��-�Ce�wUb?�W��d��l���i�p7Ϭ�*k:VOr���V�#��ΠVW��D��6b|Fl�r�4Y��cL��3Ʃo�8ާЃK�W��Ǹ����q��M�g�4�(+�,�*�^UƷ]A��O,�/����p�I圲�����=G<�����M�3D���g޻���<��f��W��ɿ�oɃB���L�,;��XXq��yA(Ad�⚽���6��c�4��8o�q��i��uEK�:�b���(�����!�+�xѥ�&���6�=M��<O1���k�D���X�G��fŊS�Y♤� �H�c�'�Ah}?
�;�W�0�qY�Qu�bO�#�3Oʢ�%k�~wP)�$�����%�i	a�O'XS�����ߠ��2P�5��#�_e��j�M��s�9���E"��]�F�xR2O?x� {B��~��_Č^��#���<�e�O6eA�,
�Dad��} #��J��G�	aT#�=��
�i&�ʤ5�'}�Ibq�I{n�y#rOZ��}^���-����R'�F&�B=�ۓ��Ok�2��j�lL�ےr����M�H�O�`%q�E~"$����T��J�A����i�ڂ�L�i2��zh�e��_����V��V��d�-`2��+}���=$����2�`����+�&Fj�5��z{��� iz�����I�����4��	\��%�j�.t�+;$iI&�x�/�V���F��u��6��@E�H�"`U��"*Y�1P��C��n�1�~_�j�+X���[�۽ime�ϭ�إ��в��u�#쒕���`x�O�*�y�?�4"��&������B���P�啋�Tz���s�8��o�5�'#�����7��Yk�Y����X݈���N#��]H���ٖ)�YD9`�gS{M��|
#|doЉ��\���G�R�b�dm^�����o\�����Qti���.m	>;Z㑅�;Nj#�ي��o�ˤ���@�>�j<��_��D(VL�V�(.�r��[��^^�?��tsH	�`d�=V�z
(�O7y�7f�4���7=���e�RFfH#���?+d0��(��2�-�gUZ��3�� ���`#"��k^�@{�5�3���$��V��<<��R�h��y���~.$�̈߰r�9؝x�j�p֐o^�0�`�����TT�#��toym���l3pܵ8�2^��X��9�Zؐ���d�D��ڥ��;�g��PX�R ��e5y�aN�f?;���� ��A���	tj�]ܝ���@r �AOH�	M���!;R�~���+$j����`������ɺm�fi�gr�;n�Vz����ё!��	�RT�,�z !�oka�l�$o~��W�s|B���[#L�m�B����ה�W�tt&k-7	�|}ۏk5���g�@Uw�Ҷwi�����Cc#���.�f	Cӎ��^b��k�*;%���M5������srY����|r`��ʘt�R�Ľ�+ӳN�k��PFŬ?�y�~ߵj�O{���3z����O�4��|��u���d9�r�!�H��{�`�t΁L.t�x~�7QW�Uu�Z��p��:s`���6@Aif�۷E�ڡ�󇁇.�?{a�i=�x�6ýEy��4�h��Y0bдyRj�{F^�p�,`�0m𺯭�y&������ˋP}�C -��͚|~#T���|QbX�,�l��n󻤛��r%iGKQ�'��꩓]�������P��%�SAZWN�]-�r ��1;4�U��o����y�2'V�:\�A�Ȃ���Pً��H �)m���x�:�����>k���,����!����~RyB^ݎ�)#�v�n��G��}���~$�T������b
n��Mi���E����v0����FF�Go�����
6(�¹!%47�%�&�y�,��LYo�Λ����G���<�������̀5�ţĞ��[�^���u�@8�*`�P�.���]�H�h�DD�^��Dv֣��0n���������r����GP��|�r'�li3����F#*�c�][����Ɉ��3_���g���>��.?fי7�k
�	`n����p�I?#G���L������� ��V�Sh	�5Z�=�}D=8'Z�=�~jc���-1?�`�r���D��Fж+Y�#)ۊ�2�]^�k�o��;�=�N�^��)\�� 2���8����$��-@�<���,�y�"�Nޯ7~�]A�5H�<�h��]fؗ��dQ�8�C��_���{�[��R��	l.�ǝ�qc$��g��i�>l^�q���r�e�6q�=�q���Dg���BZb���-�E9/�+Ή��k�1���2���F�X��`!�����E���Ԫ=�m�b\ �Hn��gf\�'�*Q��&��y���ɚ	L_\��Z5���T��奎5En��|A�T	+�~�7�ۜ5a�'�D�ƕB����-(K�6��Y��gv�� {�]��F\�U���B Ů��d�+3��$�U�W��$ޝD.T�r����Z�X1k�t�&���V�E x����9��M����- n�ScK���U5��u}!�wGR�65�'�0�d�L�:���Y�bB��Q�#l}Y�Z��F���I��T��ǚ�6�j��W衞�
���j�����[P�EF�o���K:y~Ӂ�N�0m�5��D�WPe}s�d[帻��)s�q�j.ҪN|)9�Q�喙�Rw���,~:��r�m���#�DFF�|Ƿ���^���R�Q���M`C~����q�r�2~ 3��ʒه�����te޿!�nCɜ��/�T�G����4��z��X<���!�
}��\�niq?N��Y��>�ʡN�� �l�y*��8����W�bqh�fF\��+V	�vx(BkL��]�CHj�b�l�E���5��[�y�X����1�e�oqxs!�ֶ;@�ۮ[��+���s�_?��<t�_� И�2�z�6�'PUBa^�<��gCuX �q\.?-�qox������|L|�ymԙGn�����ݼ�G&��)�Y%�1�:��|���������ţQ (��	s$��;rt�A�}��N	�(�Sy���d }ڠ�����k�ὂ���N��I"z�e-���/��l�w2�Q���[_0��@h��*WW���z�2׫ħ�z=Q�Pz,�����g�a�-��{�a�z���c���yۘ&� �#��m��:���ߍ�;�b�}c�0��U;|�K��\濛�5�SLD��� ���������Ƃ�Vk�J�d<¥Y3T��֒!_�)\Z��$]R�1l �u|A�:6n�Ƶ�
�Q���}?�r�Ta�r�(��3� �W��%�����`$=�A!�h�$^�LM��\�,知�v�����&����`�r�T�X�>Y�kd������T-��G������AW�B��aCq�m��PI�`}J	/~/�����@��;(��?�ViO�,�[��oB�(�x�@p���6%���T�1p���}�ˬ�� !���A��ʃv�~��������u��1���n�h���|�޲9U�S���).=i���	�d�%N�0h��A��A�v&��+�ܰ�-7��g�b!�O�? ����ӏt�楌�wU=�u'4��Qn Yy���v� ��C����6���џ�x���j{�dRC�Wo<s2�Op���|���xa�=+ңs���s|Z�6�L�KT����!mƶ��E�y%*���7k��c����5G��ňJ�}k�@�2	0?�ۗK���\_�d�Nh�O����8r�Tؖ.�)4��&���1�q��Z��T6�];�e,��*7���-�=-} p`���ZBd��]i���M/�7�`rp`�h�.,ݽ& ���ԚiݫH��e���2EEۣa4�k�'Owؤ��R�E�s�Ƚ�t� B\�W��FD4g�Ѥ�Idl=�m��'/��?@��/5���F��]�2�Q��+�fV9�J��*	����m�YoƔ]W���4O	���T	v���sb���&�����X��ݻ"P�Qt/R}(��0�����l�F1�@�禘b��]@9"ύ�,jH����_�HsZ�"lk��󸱇  ǣ��gGT���yL2�,-m�W�����!AgI�.������Ǜ�/m�Up ��T+�4�Af��|���\�9�::z�����
�Y#��:T�?�R�A S.%����QU�2���l�p�~�{V��d(�v#�0��m�4�?J��U�S6�I̭G���U_�O]8X�p��T6SuN����M	�+7�H
��pz�#&�smb��3%��Q��0�L�c՘�^�м�^����g���;{uJ�'���v�]i������8������o`ЇCX|����'7�� �&wS��gvf������wbc\�1�(8�(���{�T�17���=a�T�2	�e�PF �=�:�����^���5�i�����v�m&KS-�Z�dPU�A,n�j�V:��W\�N�T��� ����TˋFvf̘�*I����x3H����2���6��U_��ye��4@4�җ�ۈV@N�s�B2�g�ORW��<��u��/'H2G�~^�F�;S��P��wh��x6yQ�\�>p�-@������=
�Apgv�ZLpƵ�=b��w^���N"{��5�&����X]������ɑ���h�\'��K���Z�t��%D=�P*RG� ��%^��<�#Wz���*q��Nx�G�nO;�]Z��<q(/@;��ߗ��F�͡�۬���a ~6d�[�~ה���Q��,���s����Hg���GAZ���8��������/��{��'�$��C4K��c�P�o�\W/��Jc�����[�9l)l�*z�24��Y7��>���?I+wh�Y*��vc �����M]�xB���3Ug��I��c�7�(!M4����z �W~J��Aκlw�J� �)32Lo���Ru���;�5rH�~�8<U��/T%�O{�۟���VjP���dwʫ�)�⒪6�0x���9f���4�"��]@�H�=K��Y%�V���rfZ���o��T5�}:%1a�����?30'���zq��x�:��L�0%�W��IC&ɝi]Y�S�����*�j�^w,�O���$�����h+ ���GHK��T0�1����� tfl�����gV/>���pK�u��P�Q�rf�w��1�E��姺�'�m.1�Ƅ)呴$�[�x�My+pK��6�������$�9���Mf�/O?���G{몐ī�x���4��n_�ά�����h����"t�2-���;>W�K��~g���oj�6�e�ߜ=�ȑU�{�w���m��`����1����'�G�.)�Y�@���r���;�k�O��%���XL����}AH˨;"r`�P���T)d����7/��+Em���j�'�&����L)l�P����b�j*RQ�df���:5UF��H(�.L��~jU��Y��w��Ϲ��@6����j!��� ݰ|CnE]!�+�|�za� 𴶫5y0E��?G��H���}��45��N������A�z�a��6l�pp�>9���8��#f�nw9��6�$4
߉7!R��pK���">���v�ᙢ���h1a���kĻ�]צ��w:��Z�@�/{���Q�!��'Hf���Sq�o6�?|巰2�ju-�|���*S o63y�����X�J¢�%6F�b�J�xlHZt'�HR"�[��<�&����!�U�)�5)㴺�Fmw�b��G0>��$��)�b�v���X��t>�Av�M��OĵJ�*�.Ĉ���bd<Q1Դ����ԥ�d�履ԘW�;N0xH�ڭřY$��#|*�b//hvH�<E�1��$��g\����`�����Ƹr�0�%
N�n��d�����H#�g�Ɔ6��	�6��f�/:g��Z��
��QJ�fV�_�L"񋷸��-d�QG�����t�ӵ�o�	F> Z�|�����Y���5���o��CL�;��[���DYr���s�l\�)k�k�$y	���xW�EA�"zc�J��H���o�(M�g:�l�G���E�a(����A��I��T�$����]'ܐs�$��EB|]KS�ב�a����ңp��
P�)��ob�u�	�QS:���.ނ�h�l��}�����J��!�ȏ�mm�@|j9zaض"j��ɟea����'kǘ ��<�s�s�y�*̧TF�b��(uUK����������"j�z"!9�g���՝ �?�BX���� @0�@�3�j;�B[o���ŗ��@�@X~��E9�Lя���fMVŦ������ok8f[C;�Vi���x��\bU��-wNc��� 9ծ�_��]�/,�=�(����Q7����tl?SE:Z��@V���Mx�^M�n8 v�Œd=�pA���w��oͶ"�H��}�l-�C�,�G6F@f���Q�ʸ2	��*#��!�_�&݊���}anʮZɝ	�.U�k=�|���w�z}gʹ���YVGD1��dX���6,� oZ��rq�������+�*�������c��?W;��J♟���!%��O���vxU��Qf�:�W�| 	�x�E��)ke+��#z��M��DI>Z��k�k����b��\�%F��``���@mV���D��es��M,b���F�fs�E���9,�D��]9�-�$��h?{���!�������*d�U����xT9^��%^��ι���o[����>#�j��$�$�qDJ7��?���4��hwL�c�����Q�ec)��oL�(�����0@'فb�Y�W{�D�h��"x�7��-��!�T�riP�E�\)��ZZ��MU��5�:jҌ?�)^D�qӈ��)���3ҭ�
�* *p��k51	Y�݊C��-Yv}�
���+�XD�1Qۈ��)�o�0� �.1V)�i���%��5��Bp-o�2zs��Ί Q�X���l�쓳�g6��U��q���+����X�ٯ��jPxK���쒉�
����bS�^-��f#F�>G�5X�2�Sn�?\Ad�G%t�)~@�V��m��?��!�H�t���urSV�߿�~=���C��AZ`�h&�y��8]�$�3��@K�nQu���5�G���L�U���֮c|Y�۾Q���cd��C�T�����U�׽{#�6ɠCؠ`hn���G�/K�����x���a��f�"}Eo���Z#V(�=w�PY�.%c͈t��b�_䅒G7���,��}�s�@�&f�����&Pj�T���\�ǈtJ ��k�sL�����$C�7���p�2�m��n�����ȣ������{r����T��	��_$��9�����T��!�XDȰN.��N�J=�DlF�v�I��J��o�����Me����B�U��\xh�Rm���*�<2�%Z禿���G4�����l�ӣ: ����<���Z�C��z���G��>/��I+0|����L0	_�ˁ�F�$�nLGzKv�/Ϥ T+��Fk�O�%@"h��8�;Y��Ť�U%ǰ�g�ގ%R�9,��dK�F4��,=3K���4�`T{g��ʂ2J(��边E3P��γ�����D�x�4v��wRNw�R	yӹ+ʋ�]�4�}ז��&�0F�4P�s���[ӎ�~6*����4LY�h�������&�hmA�z�q��:�g���$�-*�.���&���Py��D�Z1���xH��Td�տ����Y���tlF��_��-�\�1�6	�Uiծ+�b����@}��1u�xD�J�����#J$E��%�&�Y�D'C=�!0�yґk�@	C04�ۙ��V.��wy�|��{9BM��8�)J#�)o�6�囫���#�����y\>�89�W1x�$���$���������>R�h"�8�A��V�G߈�(�¶�x�,Jw�0<@յq?`�H_ӆ��\��@��G$��7l�c[Oj	[��q�d� =`�@���7H�(�M����X����L��*徹z\��y�@��Ye��qQs>��_��lO�K����)��v�%��S0��&#9\��?dZ����ٛ����{M1w*��=�i��?�lG�z�"hp`{`l=���y,?�
�b��-a产�r�4B U��Δ:J���\��dt�w���N +�xj�_N,��t�P4�1U�6���J�6��^q�Q��P������1�?l.�Кb�7n7mQ�ɡ��D����2K��e4;��rީB ��?�R&ِB�P^�{��e�į�[�@�0��E�r1���u��8������ˢ�HƼ�O���fR�E|�����6Jvwo�&�=��6.��ڋQU)��Z���[{�>�'Ę�dj���Ŭr�r.$�h�}>D���o�(0oi�Y9��$v�ݼ��j�Ȱ��9����7��y�.M�*�˿�5
�:@K|{A��i����� �_�+4�n$���c��X	�����Ѥ���\�C��ʓ�~7rjP��T(�\ٻYt�>��Fj�$���?�;l��؅�P�?
wؒ{�6����G��G��ͩj�� �#��7N�\
Ǒ|�
L�d_��s��VX�b���`lB����.�l�hzլB�j�;��CYM�VU_�IM��TKx�D	��]�|@>'.�yv��U)��	��\\�֎R-2)�ވ�)�r r���rR��F�2=l1J����mUn��H�S�'#	_E����	ܷ#�9��t��3�'���/*_!V�?�w�����mu����CJ͔W�8�S�
��+�&o����� ��$n�Q\euA�R�d�]%A"-Ìܐa{�[��J@w@1^�f�k�S0|��p�ۺ]�&���{����YI�</�5��q�p�nwdm8����2�?,��C
�i��?�t�8 ���,��3��;��B�q��ʮ�^.#��9!Mٱ����t���F��$w󓮶��'�!�����*���Q���=S��p�39�6��W��o���;�9�9����J�o�sU�/���7�����H8;�U{�_5��)��f˿#};S�V����*�s-�#�)��]Z!��1P�!��V�'2��$�M�55�i�,�eu��"]y��]���xr3�V��<|˚ �d���@�O\�jT�(y�'��/0�#��]������1'�cZ���^��IMa�Dg�\�|,���w���s����)��$Iv���!�-�N�K��q�X���q{�be|�5�;����xC�Q5�l�y�IIc�S���Zw�=?���9&�֖055��T�y���U���o�y������U����;H��	����e�@����_qǧ�y�3Ńu������`�r,
Y���rf �6[ n(������֟X��)OB֬�og�&9�ht�[���.{�$�k�������D���hЁ��7<@��1DG��D<_֤=wȇc�ʥ����ż���I�]X��{�j�@�Xt��L�� �ꞅ9��� �_7������+�17�Z�K����s4�5
�q|,F{a�ŇJ�|�������S���\����[��&��t��,���
Y~���Dl�1:��RK�M������s	/�a����b`I�Xp�E^�^�Z�;�k�0���s34.���9���_��w�I�6��X6��ogq�**�*�ޯͩ.��	"�W���h���A��?������j�8Gq�6p�7|�S/�q�1GyY�:������XvkU`g�*�q>7�W��w�r0�Tg$o�E�N�>�cƽ
��-���oh>-����\-a�H�PR>�\�&J5/�mF2p�iGk����?��������\�݌��1��?�Pe�>Dg�%�i�Y@�p|��O�(��ୱ�#x����7�ۈF�/�/{,�.��.'�|�E%y������s%F�y =�����yi	�<����Ճ�G��wK����a����꫖pV�`U�`�H�c�T�����Տ$�*���wz���������i�B&ҧF�!�}��18��-��[n]�-\�G1G�����S�p����H�Md�8��y]���6�o�]�|��8$åT�O7���N�S�O�C%b_Dp�n�8�#�waSf�%�}�gY�6{g����c��JL�Piց����莭K�7�PM����BJv�W@o~6T����Ri����i��D��	rص����Z��P���nZ3��4�ڇ�Vl/ �����_�!Sw�4�g�X��� �x����P����֪tpk���r����Pb�[׼��~�{��n�ь.v@Ua�jnn���2 �}TN���&I�����H0n:̍$'Ž��C���)mt�:��/��ͪj\;���N��(S޸�/a��>'/�W#O�*6'��e�c^	/ۙ)���=d������"�{k�G��K�䉭�B!{} 2E�Ʀ�L ��@v{:Nb,_t3���}�}��*��|�Q9��N�0x��IJNr��iI���H �3z���}��w�@!vS*HX��%�H����I�Ű4-��e5��y��Ct�曍����-M�`�|G��k�H&�q12W ��&TɀK��^�P���<2M�A�<@ā6�S�HO�+/�Ɔ�ԝ���5Q��AI@��*���1�sو�х�5xI'�a%�Q^�.��!�y�4�����?�ꦞ���Tv�/8�UY� �馣��Y�D���n+6�gg]�����p����s�u8T4�����bMT�I堰*~h;����d���X;_�.*">B2����ᔫ~��8kq�{���6��� ���9���>��o%"_1����<��qi�e�ɠ�y�(���i�:���� ���� +���f�TJ�� A��?�"
*������j�	� �'�r �6�8�#�ܴ�V?��f��Z^�7�򧥇)�t"��`vN�� -G���?�u�c�.������iO,�@��@s����+7n�E��3]t�n�6x6@z�O�v(���P"������z)�dy.��Xij�@c�|���p���$v��M����ɉ��>�A�CU�:F�U�2a����ҩ�>�{�_��Y�f,�,�_��-eG��H&�u�~-q0�w# u�ap$�3�	�S��IoN2�'dDu����D�.�_F���y��".9�%x*�*�.����T����:D{���G~�sU07ft���r�����~�r.Sy���X��0,�d���?�a3��=�����0}�:J�s`䮄���C�Iy��.'u6�����Qv�+�ܢb�_m�W�0_�pK6�:�A9�K�����1���9�T�	Y���ɲ[�JFf@�_6浦7Oϼa��ѕ�����<Ez�ۮ�_��wG��&]���v��ift'w��`dI�̆��V��I��`��ikG�}�����Q�j�������G������vhWV�g�8���筹�ol5���O��Y���!�>4&�Yy���Jm,�y�ǳm��7��e�v��"����t�Nl�(���U��翽)�*�۹�ј�'.oH2��o�����J'E-�X���Z>]y|i����ٕ��1�v��a��#�2 � ��yrԒ�",���:��gƫ\ߍE
���1s�s�jq��zcA[��ē� 9X�[5���x���՗@�AX#}��z��Oچi��!�.u��Nq!�h���I�7�Nk��=kH4�u��' լch�E�W�F4{�W �fPΜ̕ >Xj#P��/C��C���:��Zߗ楑x����j�yr.��S�x�[��6��k�{~�I
�^����uO�}�{�M؊5J��&B0T�+�`��{�m��޷���w����iGm��bR<�A.�<Q�!R�.���˰$~R����OǾ]9N��nrm�����6Ǌpz2Q,�?���c��!凁��U-.�Rb��Ƽ=�&��gN�Y�5��kD��,Wd��8����-��l7��7�1\��1�wf��0����t6�x�e�R\�Ab���Fed�e�2?�D}D:8?L�6uơ�� v�g'�������;hu1�	���"�z@�%䠍0I��f�b=ekfx^nC����~7�LW�fV���Yv5�>���l�F�s�,̩?��yp��p�b�y�^��\e?��� v�(�$���97\cTY%k��1����"ޖ����ב:ڎ;�7憧A����q��Z�:��[#@A�a.�Ob�m����*�=�����#N�2z2����cX��z�����t��\�3j"^��r��W������ܚ<?���
L�sT��d�Eg���?�Yt'��^R�9%q���*�)��e�ѣ�6��������2�f��j��xC�~?m`�䤱=�#iֹ¼^2s�	/�W��Z��/6�i��L9h`ݰ�v9k�3�9w�9IE��T�Mij�h����G�D�x�<PP\�_�e��;l�)��3�7f�8x��ob*�G�gP�2��?z.�J�y���HW��t���}���Ļhuq�Gl��ע�=��������p�2/Q	S)`����)�1�B�g�;�ʡ�3�pг�@���u �TU�ۥ\Tujkn<!�\��j�x�,IId�*2U�hb�UYEvЋҽ����W}�$`.����`�DT�Q��.�v���	CfI����9�����`.{�c?�v��ud�Yt���\��0�.�
�1���3��$^�o1�=���nz�I�+�Mn�Q�ʰ��Ҏ�p�r�-9�<*�X�����hNø_%*�i��ޭ�1���#��>���	_�dɃ�|��rB�Fe��2Pf!��e�����{��R�:3YRJ���֊��%d�mm���Z��b�'��+��Ġ�	���Tf*<6I-��:�f6=:+�9�iw]:{�!������O��u��h���Cj���[�}u�y.<�dWX�r�p��F��3���#��c��Sh�cj���M_7��8k�Oc�k�F���qd�E��z�+��(=$��J��0�^����
�w�,y'�wG�c�Í��y���� 	�H������c�"S�w�^Z�\d��a����I#�S������jشq���R��'��n��z���;�˫<{�LB/���"Q�i%%��6&�V<|^r�������.�Щ���� N�0�� HkO�ɝ�a���o�L%�~}@��E76"Z':����Y�/S�m�6�1�kUQ��" ��릷I�7�zҕ��k��I���&����N#�hl�8H7��:��K0��x4�h"���1
�r`e���?66�'���lOW�L�R~����;[���S��:�ɕ�[&�N�W��F��b���m��T�>V�>��P����mO�r���c�/��)A�Ҽ��lz����Y��_c�Tߜ.e��'Q_Ô��53ٰ����u2�7-�w��"�QtR��5�,����z��,���A�;Y�z� V��I2��L�.�)!�OA5N�J���H���0�^m}��?'����k[a�_����#D�qr^W"�f"vj�b�'�Ic�] �۹8�[�t��_�'�M7��.�\r*�E0��D�ޟ��5j�t~��(�lR����f��u�㴋��n�7�,�R�p[�a�ت�q��h?���G�n8=����L��Mj~�0/P�B�Rz��-ےA)������E?s2#H�o���6��߬��5ơ����x� ,<��,�Νr�M��ԥH���w�h���ڃ �D��iF�@z��W?ϰ 7M�s
04�O#����~���x���b�����ڻ���j/���K*��i���p,s�)Y���U:�n�ٺ~x���\Ƿ�3c���Fi?�*#�=�.�^O*p+��z�9InP��D�]�;�F�V�4+��/���;�/ &b��5GMAX����}�U�b]�⥿l���,qG���$wKTCL[���>�b
�06��Z�G{H}��3n.p�t�	*cq!��x�t�j���xX�%��Ȃ�d�a����N��X��p�-�L�^�hW���Q�?w�.Z���?!{����ȇd�����X� wtFw��Lz��*=�Կ��Wz[?(Z���B��!��i�����k���Jl�9­����`	����K@�82����I��4���ա���t�0E!!�޼V.h.3��������h�����W�7nA̠ �t1�y�����d��8+���X�V`w[��t4J{�(��֒�췾��	� `#�3шA[r��'M��IIM�{dCϧV�y`����@*��(JL���Z��Y�����L�(00[:]��o��I��P}@_Q9��F����a?�{ːtSӵb������;P<u7�]S��$��@8"��U�j݃3E�Oy�L`.�ΦY���ϑdp[��l��/�MG�+�܊g�̇6t3�e�Oѧ�H[�U����z���m�8!��0��#]�z�f�>_%�z�
��ψ�#u���	�D�B=�wY��}'�6g:��BVbj��A�f1Q5�����u��V����	�@{.p��:Ii�\J�^}
�egF�e���g@����5X^�S�aRMK"��Mv*쩋fH�Y|��.zc@m�)�-D9jѲ^50܀�K����7���'��(�P�CD�=5�j-�䟐_�D��yv����p![�&&%M/�ގ卜���q6Z't��q�Tm��U�+�g|a�>�dߒn3#��(�F!��G�j\ϻOc���ڜ[<1b׫�8��*jG�Ⱦh���o�;rߎ�������ߗ����E�V��9�a�X�(4�1(���U���P�o.a�zJ����̍?��i�AD�+����M0&���,�5#������)>5�=7ez��9no0����}���Bd(yϒ��(�:�k8ToMcNz#��I�����07r�D�F��AD��4���n�V<'2&��Uf�cp�D��YD�cX�H}����/�n^W�b�?��}�mE�n=��	�7�aa�:�H?{s�@�`m6D�����µ"��z<�[�+`J�{E�2	�ViH���$���h���{�t[�������}1-�;!����O(����bt6�1��į����+����<?�s��>t�p�-��I�Eff4�����ܹ���ӑ�eoL^w��7�dSv�:T�0��b�Z'�|�|Yg��q8��Ď_1��ݨt�6y��wk4hwHY̿R-�%�;w�ǪF��ӧ����<��ĳ<�ҳ�*9Z��(����sCʯ��/�7=2S>⿊ڿ�_ͺå�#��YE,w�FAB["W,8�k�/Y��A��j�צ=2J�����?��М���^+w���x�y_�u�>s�6<q��/.���-�n�O���K��=t%.�^LH7};���&ٓú�)�dv���r��������]��)5VUń����3�c�b�W�P!���W����Y�t����.�Z����}.������8��.;6p�ɤ��._	��O�(��(�^���g�=�7�}����l������I�ߜ�|}"�1����$�#��om��#�A��vT��e�i0s�`�e�3|�i,�τ"8wg �y��Jze��̐�6�n�_�៮�f��Q���'r�j��!Z��Ò+�qF�lm�cm���SD\��e���A:���p��ڌ�O��Y�*�rv���s�ClA�Q�w)��n�&�6珡!�����*M��QR�`O;�8��~[֑C�S¨l�Ӻ�R[y���?�*�|8Zm�f^��/��ߘvQ ZL<�ܼ4����ض�p{��K���+99�1k]��}�N�{ݑ�uPsי��aj��_G[�o��g�@v�i��L���:���T-*ڒ��(.e�Q����{`z�q�D�H�&>�J;�"��uS�WF� 4�Ƀ�6�n��
�e�U{s��$ZO�������x������]m|4�H#���%�,���R�������V��K��b3���F1�F�ΗM�C��'M9���,��kʧC#ˆj&�#����
�1�3�� �O9��ı	~t�rJ���,�Q=8$9�k����$�uf�c��!��^�4h"ƒ���Go�jA��s�ٗʎZ���-GAі �7/�Ql��I�b��ǝea.?j����ݧ�g�����>���%'��l�ɡ���u����h�0)��
������������a�w�>%`|j��H0
Q!�pi/���
Ϡ�;�"G �1P��JA#/!]8k� ���y��X�=�H�%ު�;�h��蒞+�!]&f�NB>������79`g��=\�G*�IVpZ΃ ~JD�Ls�I��=5�@�$^P�J�hI��]�i�X�Ó�9��)HH���h��u���@y��<�(��
����r��Y� ���X���B���G*#�.մ��(�|���X�C̞#d����h�::2�O7���rk7�;cT����_�-���u�1Xy�Sv� ��D]�����u7r�F1A�-Mad���,M����>�|���=��k�h�G�h]2��,��Dj����Ύj	�u�W�ixf��'�j�{4(c9�N9B��e��S��nT!��۝�ΎډP������h�F�An��ܶo?q��=�}��T三���(�p� :M�5ؤV��!!��6��'�5e��֦¹5#�Zߡ�r���Z؊1�(XFN}^}sg �j	��4��-"�b2u�8�y�15q��כX3&=�#��>�=@��x��|k�v�,����实�#�>p�WO����mb-v���b���m&�ـ��ז�ņ�S������xa-Wyl�Oxª1�bt�2r����Q�Ɲ�Qy�싟<t���SI�� ���>��5�I���\�1U��^M����9F
�"2�����~כ��R�Y�O��B�&V^ܔQH&��؜�܇�4�MS�E4��%�|h��g�]O#�~�l��+.�DO��X��`�4����*�N��_�Ĉ!��Y^Y�{�cZT�l��|c����1��2��������ڡ0#RaނbsˁiϮ�&��D��9���r��ƒl/i����:K"A	��r��]�s�~�����m������6���Nt�?Z{���w� $P(
�	 �TϨ�����%��ic�c�dx���1ˬ����=3���ݫ+��hK�f,�4c�|�-�Y	�Lc��1�p<��?�D@��IpJ|Y��� ��h.��	�'QF)@�!�v���ź�@�xr����Ѕ�[� ^���t��ƛ%��T-Nhq�/ƧM���p���Q��F7޶�W1����8��ٹJ�w�E�83��T�����0k^^^��������|�V�'���	pX*�zPC9Ũ��&��ɫ����rz�Re���f�Dڹ����D3u�R� ���$�,�]0�ׇ5n��e��]Aٜ(اj��o�"�ѫ��J*.��$]{�+�$�?*x#���D�!hff0{��0{�BB8�E��TN�׹���>��<�\F(�'�ߐ?rM�m�9ν�$�o�\��̛���m�Z�2�<��z�_7_i ��Q����gWO�j�C��!^���f<��79:K���=9L�*N�F*�Ņ��Y��A�b��\Q%�L�|$�zA����'����b~�����Y���E�w(�*FŢ�h���mA��NA����ǯ�|�H�=N�Էt�.K��i��9�
Lm�����K\�-����e��1j�����6x����X��h�6A�A���j5m����}���
�S�(}>m���&\l1Z�߽�QK��x�k�®$�\~������ȝ�>�����mC$a!����}oK�,��甼��i�$L�G�0�ؠ�>���*��6/C�C��_g���J��$x�4Z.��'�ɦI�����v��*��rYa����C5 _0Ddt��u��a���ql�b}0�jdr��7�h�.�����MZ
B�n���ι'����u�g6�3������ il�)�HlkJ
�7�4��`��/�I�B�U�ݗ7����s�G#���w>�~��T
u���ӵx�l��F2�0�oT�=>����
J�䟨����QLr���W�<��Fmc�m��uLE:�HnQX�G:����b��m�'�.*I�'���s�"$�"f���*�0G�_baH0l�n��u4+f�N���E;��iYj��a؊���2���T� �k��Pͫ��b����������TTnӿ϶���׋=	~\��z����	�!�-G���B�ڡ�֧�F�����F*����7�͇�}u�<���8!�6�B-T��W/[U;pS�e�@�[؞4�0��s	���fM�v���D���J��g׉.D��Z�tgRW��"}�����N�������Q�`��V=�!�s��0m�R��?'��#��.�&��G}��O�;��(�uy�������+S��t�2����s��t�9W�I/TW�4G+�A��C
+ZKF�u86��Z�)+�������j*Yoo=/ x i���\8C]�|\A�f���M�ȋ�$5`�%���������[��G�S�ߥ5:ov*�p�C��i�`
Bg���[��@	��E�V!4^����x��f���%�X�61d
f���@.�]EU��*r���e��u��s�rq�?w�M�";���n�o���ӱoAJ���I��0�ǔVE �j8�k�n��I�8�����`Z =�8;���]&�#�ZZ�Y	��10gU��7t��,���V��!�G���p5ֶZȟm3�ڰ\߷�n�5��~�u�'�)�Nо��rx�l��<q�z����a�wq�ž_���7ˠ����8�9��4�I����/E��x��8Kk�K2;.u�O�7�S�7&�|��;s��6`���e�s�(���9�'��Sx�Fm-�f����#��W{V
��%�m��e_C��h�Q�"e�!��m1o+�R�@F2},�A�2Q�b/�N�{)��'��0��qc�`ٛ��gXP���d[`�=`fF�A �6��ctۚ�VM)ɱ�0A��A�<rtP�JdZ�ͣE�p?͕t�ȁ��u����k<�Ɉ�SS��8K`�`hQ�x.�.gN�&5ܺY�'����s���`|k�m��ry���X�����J�v��V`�M觿F#��	E�S�p��|�1M�Y{�ɈǷ�w�ѻ�{�v0%Q� �4�ʿx��;�<�=����]B�} ��6�V�*)W#���14�ġ"���B��AN�x���%��ث)�YM��F���@��R-��e�8n1A,����kh��q�G zj�����9W-A,�P�Ә°�'���v��&�ռ��y�.I���հ q��^�h�T�&�ʴ�� ��џ�>#J�Sd����WG�j�K#���}*^ٺ8��TI�C9�B�~3,/�u�\ShP�z�XT��T�~�����
�"N�	��/��k����]1Ϫ�Ő[X� �a�y�CȂ#.��2+�r豭u���q�bT�Ҝ^"j���ie<��QJ�f������k�1�gvA�Ǥ��ߎ|��=�_���4=[t��	�γ�	�"��R��x&�{Ԫ�b|�Ã�!j�r�z�l��mu��Ks�qO�Sd�<\���U΅,��/@�I�P(�Y�#�Xd��(��E]<��a����{!8��!8	R�m��3C��O c,釳P��谮>���l�����}.t �j�F��ޏ�V[#�q< ~)�G�3徸'�a�k���[�Hӌ7�St�1n�7F7;�͇��ah��\:V&��w��:b�!��.D��4�H,U�Y'��rҸ$ ��a.6iy����C�k�I�כ2L�	�%<�e�a[m�Jƥ�`)�8�O��E揝]���z�g�"ι��a;�r8��C�Dŵ\MY 2Ϥ�#���}�UJ���)Qnjv�o�k��F񉹣yǐp��V�ϋ�$��m��
F��m��Y�EfK�^
W�qa�.yM��tv@\wyٚ�c��{\����$Q��H����S����Ӆ՛B,���o�������rב��T��ӱ�wdJ�.�j�,�Tw�TcB��]�?+�o��<�(	�;��?�/�3��{���V�d�hL0�My����uf�V����dD��I� �e}$QbCD���y436���+v��%nt�$/Ϟ�^$�|���'���Ε]�k����D� ��6B=𞀦ǁV�CQ0���/��������/_�i.Q�q�Nt*=�o�`y06X�(_CY�����XУ�n�����dh�FR�\�Դ�+),�\���� �#?�њme�<�i���qK����Θ*puu����_V��joR��`5�:�D~n��Z���`��@U��?5�fF���V�e�lԶ�_���%�F.�ы~�A����"<u7�Ҭ3
_�_fx2���RL�o����,F��c&J�gǈ�ELk@:e�Gۭ���j�H��T��W(⨠'��/R׏�b6e�v��-
C�lꔌ�i"3ޢ72���V�w&O T�J8>����V �@W|����g��<���~Z����T����ʀ���j;�~�6Fg�,E��Jb/�O��	�X��x�Jӂ<���dfg�{�qW��~wR��	s������V����N��;���}Өm�5���j�+���ɯ��#��~���<T��&LKx,=k�G�E��F~n2�mn�%@��x��I�v�N�"���#��D��3~��;�t��� r�69�J�YꑒJ����,���e�Ֆ#��5HΟ�o�t��u�7�t������F�
}��#��:sV3���Kl�1��x��e2	$۽QӱHCL�w}�ʼ��� }(^4�෰�2ĝ|�0�oc����ew/]��	�}!�N|�H��ە�az1"��S�_3�5�< �lj=$����Y^� �k4���h1��z���#c�(>��ǭUJ].�&��r�9�0�)
N�x���cv띻OX�v��X��1��6+�[T�5S�|����k'�v��y��n]E�>��1+�X/�>-w�d|xM|
�����c@sl��������ށ�8����Ԯ0pK�����Yq�')R����V��[�/�� H{�1pC}(�Q���O)b������c*������F e��}��SkVYa�Z����ϟ�B��$qK��[G0zU��,���ο�[�WGi�Yҭy�L�B���ӆ)��4���D7eI)qx�C#�q<]�D.L����>��[�w��|$f7��K����:���C�� s~��Z*|2�.��n���P�G���V� �u��ى�V��3��3ھN�3�R��&�WZ�9�F�ǝ�Pڔ{8y�\5�#�Q�h���w��
=*9�GYp��S�s /���i����Ұ���d�I̟[���΁<<&5Aj�mv�ǹ�r�H�*�(a[�ˇ-��F���_�WXlxQ@�nb("p|J�S�r��yeN@��1�j�	�$�V|���w8����̓�=���D|DsPf��>ݜ	�H��j,������OV�=o]��� �8r����׳M�,�\���X�+�?�q��fkd��i���Pv��l�|���x��a`�Q�[v�^��e�3� ��cJ�t���s��=zs=r��ԭ����w�V۷�x��O�2��؞�����]��a�w&��k|���K�>�%�ke�j��QcU�'��C=φ��M ��J
�ReF�cT�cj����� ��$`D�A7A����?\=>�n[�6	��V��U�tޏ��K�M���w��W�N194� 1�l!��e�K���A�[�.w�n�n�sc;�����:V/��6xC/V��Xz�Z�'���f5���d|W�m9#��x.�תR����&�ng;䝕Ô ���HF+��Iӑ��;	N-J�F��T� �Ey��,]�Ld���o)O�5���ـ�c�����lۂ��Ȍ�N�E��
%�ezc���ຝ�j��*��w �Z��b)n$�c��])ȗ%�~Mg-�|��(�����Q[�bZ�T�ͣ��
�Z�H��2��}ƦQ�R��K�0��*�{�7c��U$�>MXl.qH�8���d�������!ٸ�>��A9�HSjW��\���-�Y���u��ޔ:�sP�T���7G?�Α�P���ީs�~��ΕG�|��Tŝ[c�;Ix|�7��TJ'����oS9Hn��ޢnk�|�77����h�M?���>�]��3x�r�����`z���(HL�釄��ł�:�Q���"�>�!�4L�.��VS��b:mU������,=�&��V!�(���wձ2�j%絵���nyԚ�,�?��8�0�N�Ot��c�M͊=�!#b��g�i���Ӳ�F��*8C`�k�F���Tdō�&1�=!5[������EX��Z�`AY�aT������V��Y�@G��3˹�������G�Y\4�:�5�D�g�{���ڕD˜q�7l;��ȯlB��a������%�9���O��4�*���DH�
��!D:�K�,���	�1�&���{��L
4�g^��.���A���4,�F�3���r9��K�m dسۧ�i��13�Us�m���0�H�+~&Tm��Mr6Á��m�X0$#Y�
��$�S�lʰ�Խ�Nb�x~2�H��/�x"��7ϰ�)5�O�����1�b�*��d������n�
�����Ľw�]u�0�]�b����·܏M�����^"'o\MU���
c"�g~{�֡3{�(������о;a�?�X�2���y%�.ٺ��� �k�{�}=��`�3�ƋZV{aq �W��90x��a�����4�:D
��Oҿ��qQ*�L Q�7>�D�=q���8x2��e%Va��D�<ˎE��(#����"=n|���m>���v�_lP�:z*M]�+����-
�#34x�E�^h�Co�T��NG9
��}���~��d��K��y��Hv��M	hJ��r|�Α��i���t��m�F����W������y~���HA~S��'RA��]�����������"n����Q4U,��	˰����z��������,����i�꿼��Y��[�վK<�20��/�)��������t[����5�/�d�����O���Kk�����L��3� �F!���r��5��r��Ug�?:=�gD]E�^{�%1�Us@��h<oQaӯ���ge*�C�'��ؿ�g� 2�̃��\
1!?n���`����4o2-�Lc����jU}.V�aA)�'���|?����:+�Ԟ��u�q�,2@+o�̠L�̽���_��lʩ��0T�¡;z�����	����]˅ [�}ѳQ_mP����`����;��0L�y�����w~���"�?�����T �,6���)����($o]eK��}�H�cP�v�b�U���c�E"RƓ�S]�'���T!oM��rVd�l`���G؏[K�]�,d��.=[��ھ���(��s�9��_/�bOd���L�0�2O��(� G��A���_� j¶d�A���w!�6�&z�� *Y����0!
��V�0&��8";� ���0��h�H(<k��}���g~�m:C4�MA�*����y��0X���\Ff������*��`�:Ȍ�)���
�F�3�y���>���}z�)�����?�p�5ې �YS}7fl��SR�����m5�9Gૐ��������G�����4���6lC��J/���ߣ(�z� ���5�X[��!?[M��F;ehF��{1+݆�q&P(�Cx��=�d]���h��!�w=�k�Y�Y�O�c����-1�H����Fo����Q�T�'�L�)C}^�E�ӫ�����[b�����9:EJ�6�-�w�̉{����rr�&��j�Li��	֏�@*�2z$$7P��X�>~�������d#�'�Adq�uk;�ΊRK�͸/�G&�r-?!i v�|���8�����Y���&ס�R{y
>g���qu���B6���v����#�(��7�%��|�*E/)_C�\���$�H>�O��Sk�y !�u�ul�A�'�Q�܀�>o�r�l�s#-���J��w���M��ƫa�TM�E.�mGF+,ڈT���Ă��0��������@��Ҹ�-$�=%�qP5��D��[/�{/�zO�Z5��s��ԩ�@hC��Q�C>lg9�x�aa����Om��lG'�Z�}T���U�U���7d�T����g�����SpQ��)��Z���C1K�J�(�ob�b�d�m	�U��w��͌�?�N�j� �T�+�Y
B�)J�Z���5
��#U�A�;�����
pt�6��	k�[�q6���|���|���*")���2��g2X�a<���c[�)�`�gj��±�Mv��'yiΏ��8�sfF���묛���)�݋P�o�}1���)q��'�g���4���*�d(v_
���F��h@�!ﱼu���Dv��G�k���-.��.	#��a5���
�'u�����&� D���ݛ lg�œ,�����j�."��Hm�!~�uݜG���y�����Y�1�/E^��H��We��&#Si��QH!v%t�Y�I�.��x�+��q�6P���Q�b˗,��A]�=���y�@�CIS#D�z���.�4A	�s'�i@�9���su)�$cp���D��:�\�[hj@�k���C$��r8�r��p jz$���$k��`Lߪ������?}�[ r�n(�H��JJ��&Igo����.�TLQ��_���M�GQ)���w�#=}�J���N�g���+�~�fF��u������Ӝ��_ND��<��(O&q����4��KP�*=�0��������[h��N4�a�2<ס�R;w}W]+����(�����A>�8.�1\T�G[F���������Z'7O%� <�
�C���2�d}MCl+(I�����\8�BD�� ���1�6���ݳ|�ei%�ٞ6-�?ɻR��'v�_�������)f�v��T��㷏ﳢ}w@�&�M�Ϋ��B|�do:A�������x�mC���gв������wQ����}�����
�:�A�����X9�*r.�݀�0Dg����apK"H�.R|�V�$.��L֧`����X;�� �����]�h���GX�'�u�6��x�@
qf�m9!�>w�^@�l���U\#�G��1�-Q�D�&򜢏�
e��'$6���t�"��esʱ~6�҃�p�����kqj�죸N�L�5�	����0U�XR�N5G���êJJ���LE�u��D��� S��D��6է%?o�Ms�N�	���1޷���w��v4J�|���-���YGs���l�`IK��<eozy=�CC��x��jGؒ��_L��{�۟�#&��r�"R?��	q��}$:B�o�!���^G� »��&�E�c0���U�~�<꘣Z�M�&�7�x.��YH*��9�I!���B%��w9�J���s�@����V�e��ሩJ���A��sb�,Ƒ���^D��t�s#�/�c�<�wt~�9nGK�	�����#�3�W5FjJ4��Vn����Ƿ(�ʑ�RPC�qH����L!���yY��Q_Ш�ö�¿;�a秅�E�̌� �ǅ�呹�
�\�f�h0��������Z��I�襾#k�]�5�.t�Qz��������l#��x�(n�4@�h֙�7�8���9}~���/KǇP��U�մy8�&Y�{�,`e����N��t'��2��졦���=����{��<b�uo"II�E����T
�դќ�)j?���Xل��^�4ޠAE���ck^��|j����NH̘���z���]�<T�ȈƑ�l�?w�Ԓr,L b�q���j�p�!���Rp	�`4Ē��}�8sy���a����5Oɻ��c��P(��sPaK���u�	m|�ȧk�����!�A�f	HY`�ħ\��ѲpP���<!�}s���.2\ J�C⾿��SB�.�^'h��I��(��+톗������-�E�+��7>^�3�DU���Etȉ�	C�O���n��;O��S�id�e��f��N%b�U�03{x� �:��)9�Ad/u�y�15��4FX2�Q&>�"��/����
C�h��i׉eG�ko{݋.�P޸p�Ț��\���t���ˊ�]AN��2^ ��s'�����l6�	F#h�����{N���`P#�Y�BK"����$�<?h*��-gY/B{�Ǒ6^	�A^�C��XF�q�@��ĺ{a�,��z�D�lV1u7�+355�T\�w�E����G��s甈[�>��K��+��\�X�*�BQ �?J�6�k��%wX�������tC��C�dJ��XxÆ$���:�YXSS�@��h��=+�R��#&	W��,�S�o&�) <vdV���;c��Ԝ���.����("����|���=���mYKӃq�h���Gzz6�ظpz�}�v�Aߚ��X�t�w����"��rI�J�Pu��	l��{�0I�D;�֬�:T�+�R�e>s��JX�,�1N���]ւ��?�c5�e>�ȍҭ� ?�P+~p�l��EW���s���������ݴ�APhU&NR�_�Y�]�ؖME}�6 �����f+���3�[Q�9�FX�h~���PM?�sQ��A�����I{k���F�� ����F�䛱��F���[�N��&,6�0G9I���]{E�Y鸫A];�|
��Z2|Ij-� ,[�]sE�?�����{��2I V�峜�F?��Q0��hN�������ZxiX��A���~G�C�&��Х�i݇��G�ʇ�<6�x�I���i�y7�����%KP�
����E�eg1�r�~T3�巌Ѧ�o\G�|�"�}��5�=�1�`���:k�՗8s-��v#��̜EJo���=�i��/�EW�F
�)�,��C�J.����U֘ :��D��"ã|���R�\˖-U��fz��a�&u��1	-|׵x�!�b����e���x�bٔC��%u���H�����H�k�>N�֖��,�N�����f6��Sۘ`�U�ۜv��6��ܷ"*q�>�F��$��ٮ��	��.�w���?�NV�<Q���]�_a�qs�[��0���H���*T �0c����mJ�	�P�PּPi�{_��A��ߋ ٥R	�_�{����_
�)��	�u_ʯ����򈚟�M�Qv��Х�@Z��x��=ޱ��ς���������0v��[o���+B&���g^P��sedc��^���A�<�i�����+���uK)����m �bXr�VU���]��Hy��i<�ys`���q��d���]���]����w�>s���٥Ǻx��^C���mI��|@:&�؄QG߮'0�z�5�Ɵ��4�=�ͰAǎ�W��eb�.���p%����,��$�����Y��X�a���������1e��e�߈�P�f7V���S�_1q��\1"��H1ܼ�"i+�бx���]u�dƉ�$�2�JW�5Y�ye�s��U�@%��s%���Q��o@5��_��e�|A�Y7�B}=�f�e���	G 1bpA����&�|L�^3�x� �n�;�J����'�1�����n��\C)���M��^�M;2��ѭg(x���؋�B���;��|��ݰ$Yu�X�i�`7������>�r�	K��K�Y7��0���B��ySf�R��B�13���nb�b*�����7���'�ě�lC;@X[(��_�?A{J���b��<JW�B\V�L�º0�0�H�������{9gop�%���O#�i8�Q�q�H���xD��뭍���'b�����î�.w���/,[�ِ.�s��57���6�����)�8��o�H��9Tx��� �ކ�eyA�as���Ϥ@�(J:;h@�1�����9�"몳�:�==]�T:[]�nW��C�l͸ï��C\GG��:�ډrR]Q�^�2p��t%FH�	��=a��,�R��ޮ��q�_ޏ�Ϩ!���m`��lG�!s����s��-BƆ3�NH�i/➭HN^;�'�����M��^,���e�����x^�`2�d�f��Ψ{D���϶���k���~�tT��q:�sE�V�o�T�B����|d�&�_���#hgδ����Ϩj�K�ˋ}m"vY� 귮XB�W!#	�rP^��_Ԏ�������^����cȚ�8��_����*��I�mZ'�# �}^�`[�E����Sק?Y�y2ʉY��#�a�͗t��ъ�UVZ��u�Y��rml����\��c����qe�+�EՁB0�L�2�,ɸ��C	��^%/��fw?[O��i��yb.�]Xl,$|����p�W�}����W��tQt8�y���ɒ3�1cei%M����Bؙ�6�h=H�gn&}���Ȟ�Z[��^�*�����S�nr�/�¿ㄮ����~͔�Z<�桖k�|n�yI���C<����J�4!9A���6"i�����:�4�]�9�Az0��V���� ���X�����>8^P����v+��� ��= {�����>�U$B���6JΊ6~��,�8�o�}��/_^C�pp!v8W"��0h$��wBh���x�nQ�^J{���WA��Ul:�$�o!�,��GQ��;�Y?���0��+�ո'
����^W��_.`��r�/�jӑ�ǵ�a}+��ךCzæ�H6�9�C0�qڻ�`!� E^2�v����D����*�rt���]��->1��V��h�=B����0�>aO�T��8���T�?�xW����$k�}j�h�;.r�uO�b�p�a��CL!�V�!<z�m�Oq2/x��Y�C���h������~�g=�_pES�J���O����?���5�v@HD�3fmnh=&~��V���O����Mp�Xj�Xa���/>��"�i���������oRAL��_mRɸ��23�_"�<0��r�㞘���bR��������aD�2%:5�x)�6�e�:��Ak�7&6ú �ĩ��ܤ@�k0~ ��t�׺�6S<sC �m�"F��%b�����2(X�����D����!:X�{�CLK�r�}C)�e�#L@��'��E.!� d�#�R5=��v��[�oN�(�^�"�P�&�~YC6�a�j�]0���%0QZ����)Z��.����*C׆wu� �w�m���M	�n�P�k#=w�#EP�>�����L��t`��s�g�:����%�d�b��G�C���A[ۃ�(�Ж�?���{SS�]��G�}01Qxddh]���e����%�X�3Y��8�TF���i(c�n�Mk,�'Ad>_�X�-E7"ʬH�>��d��o���vg�!�1ӱ;ް�)�7�������r�Hv�jcq�7�N�_��auN�B�rD"P@X��~qX��J��6sV�f���{���M} .@(K���~e���7E�����@��T�j�@K���-C�E��v}h
�8��9�=%��ں�u��g����I�����6�����o�~%�/P���r��3���,�aڀ�;$��тZ���$�[�O7%����Tt+��7'�	�
T�h���հH�Q��F��z��8�m�g��ؙ��~�>�M��`BצQ��6���@�q1�=�]�1��)�k��8}BN�tl%D&E��r�K �i�w���ٸ�f����r�&46%q&�2�Y7|
��/3��L���T��#ս�l�sOG&�q�:A����GO���(��s`5�!a�=����2H������bjg�̉r���w�:���Q_ΞB^g�r[�����.�z���șl����+%�8$$'[��=8c�*�EOI��B-��e&�{���-s��lPͭO����o�Y�f��3�Bc���u�	ʲB"5.���د��V��BY����kN]�u���Ζ�:���eun� yv `���]�i��ӠoM܏�m}B����^і_+�_��%�i4�I,��y���6�ݩLR(���-�(�2d�c%t�M����ۙ��ӌ�G�ݿ]�g��C��-����K�	kw�J����8zC�$m���])�N0��n��u����1	*eE��� {c���"P�|V���q�/�LCx���r5����1,���"�ʜ�9�<��:z���:�r�]���z��}�e�Ug�Ъ@��d�ܪ�t�yF<���'��0R����0���M���rė�*�Ń���*E:���5"��E����ì�dr�
&��~ǿ��X���o�[���o��� \�/�Vg ���;ҊruZX�rkă�J����+���7�5_�'\mӔ�:��h2/8���0�Z/��&���fa[�Kk�H��"� PZ"����X��yۅdşj�x��l	�K�t����'�$�H�� H��dy����R�0��=Jd>�(���Ŕ0�rD
!�\���1�o�iB)/�pQ]E��zm�Z�|'<D'O��2+o�F[]����F���f���"����ʘ��B�]D�\(:�mϓ��[�w���M�Ȋ��zxF�,��οZK@����>���6V{������������I�]�e���d�[n'�U"�����ic���1ѻ�c1P��8L� ��u:�<#��S�Wk�O������j�`e�/}/ԋ���jy�cȯ|�Q+*w����J�4;�-�j���f�VLϤg������b������-z�w�ܴ��5��15�Ҁ��2�ᯆl��VK��+&1}�v���ο�B����M���C���G)`�8�͉Y�	�V�|���D��u԰�_U�q�*Y���#�_�v���DcG]�a�����]HN1tlBIB,H�����z,�X5�'
���-±����џ�G����8��C=�I3��i��q�DM��\�mTu����٧R�U�.�X�:9�oEo�\�&�;�����쥩G���A�;c�=91��	���{�#|̵Qy��m�hk&�/Ä�.�qa�s�l�f*��b(b?�*�P��篳�9.����5�`\��3����G�
�)��X�7!s�ruF�&Z�`�bra�ο]�$\��u���.�E�2e�9�β�f�l�|�}~l�SU+`|~A4XNb<�S��ݚџ���p�������d��4����H:�|/��▇�C�v]����30#��ݜƅ����7�Mƿ�a��P@cǪ}�1W��uL���.�h��w����n�GF����;9���@���K�mYʽ�K56c�*���-rjƒ�����Lb�����|���Lrm�~s,~�.\�����fl{��Y�N�]��GN{��Ѫ��O��اu��5��)����/�1wW��[EME:_$���1���]�/����ޜ�=^jz�V�7��1��χ�!F(�8�i��AkCtb}�2���Xr�PLb�V}*�����q[>�l��۵���v+Gjex��J	E������r Xbb�G6����L�M���7�4��(�����X'�Y�w`�5_n<5�C��*R��(,��%#�ud9e��""0�ʓ6�#��]YF��S�Q��X+j�/?���'��~�וщ�@�Dp)�6��Q�����$�U�.�X��W�r�	:�IZ�|��L�<|���˃RL��kX ���(��B
|�b�r�N@� 4J�~�i�'��ra�x��g.$y�Q�H^�����E!��,m���˰�`g��(��ɧvr������!�lٲ.&b��k%��]�ܽ��A��'7���Ţ.�pr2![�&n�)i�?
],�5faa:�<���cɔ��%�u&��i�����|��>v&�5A�� >d�t������O�s�2�'HC�_1�½-�o��x��L-��x��>Ҿ1WJ?����p�嚖H����e��.@%�I�Y�D���Z��I`|��9'������ݫ~p��ud%�(�� �}��F�D�3L57����[Q$��|��Z#�}�\���G�����,��!��� r�Oz~�ߏ0�`�%s�}[����r�af��q�i�."��χ}:w��dii�������=(�+7�U���Œe�y�b�2Pz$�V7&`؈�9��b�L^o1�h�Ƿ2٘&U�!���X���+t�󚲞a$G�'����s��)��� ?�U� 8��S'vе��ؖ�į�B���oX�3�#Ѕ�(��(BJI;�H��6�JXc���;�qP�>>��M/2s ���c�p8�po����f�:Ha��� ϵlU(���Btq$��T����T�S_[���VV�WM�˴=�(@��2=T�@�Yı'�0�L(c48' k��4{�dFJ�J�
X��������ğ���k?����dBC�sG�������<^h<��-�<����Ck����h��GGYa�1[-%���2���\z��^?��'UIc*8&_�x2�~�-ΖiN	��)�N��4��Ro�R[c\REr���/`vH��b��.�M�SX���lR�Ϋmgr4����E��D#ܳ��0�|�V�_00�xq�VP��L���U|F+���J��bR��6�3E�0�+10��d#���������)�W�¤����IqIH.*��~f�	�k3���[GE�����%���y�����?���Wq�fD��=������k��Ն����E�$M����}��5���O=|t�����k8ˇ�fǬL�=Hp
�@�
��k���՟'�����a�"���a���I���z��f��;r��b�ߗ��v;f6<t��"�ϧ��{�G��jX��ֽr����ۗC�^ܬ$�	�]! ^t6~`(�T�?���3o��К�WgYƙ/�b�"H���Y.����
[��lʏ�5�W��f�R�E�4Ҋ��|���Ȗ��V��h���8�̃�(r�f�x'�X_+�,K* ���-{��(��_w�m$Eç5L�2�����iO��֢.^�m���xq������jL�nΣQPd)�F�YqH�p��??��Q��<���u��I���ϭ�/���WfoL�(!ܫ\[�ސc_��C|� B�pPf��.d��!�����=N��e�% ��8�uWN��L��H��+�����F��4�ߗ�!J3���%_[Mܝ��]6	Ӣ�]���.|���7F&�\[�����Փ�|���8D�������k�b�&&!��3�Q��hb��t��'�<L]ɔ$��S�=m��4�/���\������o"�e���@��^�薒Y��ix�W�J=M��j.W�y��H�g�]^����2��ʨ��'���| ~����;��O�9��cޡ�,����3�Q��V��S�z����O�4V��^[@�g��x�,N1���jN��# ���Z��ӂ<:��w�����8z/�+y6�q�a��VZERO���L2������i)_�,�5�y�ث@��o/�_ޤ��=�,xzzzmpO��0s'��n?g������4o"D�i:�]3�̓_[����=k9���������X5�<�%�:̞�h96���Ja����u��"h�E� ǁ�����bd�sx�(�#�d��)���� o`���]-ɺn�c��H��Ф��9.ӗ�S��������^�yU!&��j>�;s�O��Wa���KH e��S+>�j�%�nzS�#b���:������oS'A���T���5�pV%�/�y7�����>|mU3E\_(���(ړ7_��:|�=�yw�"8�>�ؗ)��g��	.Ȑ�ݝB� 'a�TY�P)Ҷ���\1dS�,�@P��gw!�b���p���&T:���k+9�Xw`��afʛz��0�Is`(P�=[@�|����`/��|��wo�������Q��JA͝�gޅ��=���l�sUW�/��[\�\9�5G�Yi I��M2�ö S��?p/̮����P�ѷ���<�r��4R�m��������D	��6����0����
�.�xu�L��N�o�O�i�?N]��5R���sg۹!n�i�sFH�˚s���y��*��?�k\�1�,4{5�Q4T�n�}=�)��� *����}څ�t���=$�fV�Ťy��o(H���Txr!��=�z�t�(�4Q^B�K@�p�qi����>[�h�j`4�����c9e�%��$V�0$"����d �� ]U}E��!�9�a�����C��u�Z��̄�1���]PBTSx�p�)�,��t?��Ǵo\M�2?V��� �c������uZ3�}�Л���Z��JX���x�L�Q>�+�s�0�<��fH�g�$�a권$����#���Ge����}��Ӷ�$�I�3�8�h0LW�1�9�|��M��r36�A�����{����g��z�H[t��X�6���40�ᫌk���*q�C.q���s��牉��[E�:t�@5,#���X~���m��^��Z�c�Gs%�Dcg��%"�ܚ��>Q�k5������t��f��I��ߒ�k ��7K�["����>H]��v۠��������=�LHK�*Gy]@����>~L��5LPb~��ˏ�1���x��٨bJ�B�����	��:
L?+�+����U;�-b-���H �j��Le�U�v�e%?�:�hC��8F�UV�\廗2ş��;	h��=VD�f���o�fݒ�#nV��)�S��}�3?sIdD�pj,4�{��7槂 ٛ��P^�H˚���jq��(�a0���x��X�0a�Ѫ�;��L�P�<?W1��<r��B�7�oqQDpb�84��
��}jhJ*���iK��(!�3�V?���H!���fAmr�Cq^ڑD���'S'8@[+n۝�7� ?������_f����k��K��U&�+#��{I2v8!�u���~L��Ͳ������H�㩚6��d�����cQ��m��e>A��c3������m�}Z$
��yc���6�ZL�n7 }�
,�����ݴ��o#*x��J�y�ʿ[�(m\LU�E��v!: �ζ�;}�u����I��ٙab���X�*���GL8���4ݾ8���\�w	��Ἰ��%�%ǌ�Ēa��=�9ِ�B	�d@�7��h�.ƫ�i׍kwP����bH���53'�Ru�m��Y`�_~�&�����>g���_?f�����z������ùx���Ce�E�5#>�Zz�~�<-��mc3�����˝�Ks��.-�Z���u�_�>F���u�}�DK�.c�/�{I�l���uT�d�W�.RǆԇM��|�����؆=�����'�`���-��k����N#}a�D�c�r�3'�S�͇�t�1���^�~��O9c�\�鎏�b� 8�u�ܸ%����|_ݻ�F �v�=f�}4�;�S~z��nn>v��Q�$$A@
+ q�L�Ӗ^d�"'Z*>bQ�P��64����Y2hd�Scm`�!�&�{���Z+�����)��	\���9����M�ѡ+�x� ���tE��!i��\%F/��#�!���܄ׁ��"d(0Eİi��"���Ӆ����k��g�S�ţ 5%��.��/0]��O���dQɡJ"�y�?-�n�o����'�M4���r
i�.���Q�S�q�w��2�Q�}TʿI�K%���$_�P�O�6U
0�Vc`P�О�G';�[o�r�I��� ��G�Um%`��J8����T��;�А��[4==`ʶ2�Ϧ\F�T��2(�J�6�\#��w��=��q�H���ʻЋ����ْ(cYF^٦62d��A��XԮ��y;ɂon��N8j�l ��+h�ulU*Y|�L�@���n�)��k�2��^��$w��?�iCA%����썣y����C����<=��N	U��Ǩ�E�r��u%ɢu�v,��ǒ�G*a-L-�׍�+�b��6�F���%}\7�6 L�����"ꏬ]��qxE��'�iLԡV�~KI�^
2�� si���v���P#�U�sds��Wr S}��*zN8n�nǼ+�� ,3�p�����	/k*�`�3���}y�a"e���(˷���W�N�"Km*e֖���xL�L\����P�)�zq�=<�A~_����V1�,��������vY�`�WW^da;�2< �,	�>�b�\�P�������?C@Z�RALI$�[[��@"}^�;�����X�2����s�t����������b���!��F�>¶;v_Ո>g������(��t���F��b�	��`9`��a��Ƴ�q� i�$/�$!zs��^�01�vy����\&���%E�r}��:�"|U�K�}�h!iXh/��"�jӪ� ��>�+�����a����p��)R)2�$m������͇��Z�s�/�����0���2�:;� z[�l?����Nt�[�_�W�.
�m=���l��J�CRn��� %J<�����Z�Wv��Ф���B
�U�ێ���E�F��s��[���-%�m]��WOƯ޺�K#�W�-�.��@ѣ�h��F�gI��w����dl�U����J��2���h�C�XI2�&wޢґ�&Y�����"ߟ����n|�w�u�������������U������%%�,'�e<��usÊ=���]��%�����Ug���·9�U� &\7k"�w�o�!������~(S@t۠���rLo����t��O�qm���(#j^�$\ہ�Z�O祼�w�ȋ����9t�ܶ�qU�u�Z��k^e_��c��zm�Rl8�����|���0S���ZLti��_�/Ph5FB�vA��3�Rq�Uy��J�L[��l0�x�a$^a���Â"kIoA9@�	�V�W^�V\~�$�Ǳ��L��	�qS=?�=
$��>�{����}���%��g��E�M��,���jz<Z~`#�O]R8��{�7&�%�N��+�(�+��US���ԛ��Uf��,:,*�'����A(����!�t�r�\C�>�	�L�Nڦƴ��h�M�0�O>n,�Q"�6�
�0�~kh:x�+x��P��qE�ʀ\����S�O�j�##Umr>i$r4T�!@šw|4r�+zi������%�K.�pK��kj�&N���[*K����~(}T�R�Afm���IRmDu�����3�ֱi]�:����P�w~*���b}��[�3�&m��]���~�*���40�xv��������$`���IPZ��
��W�/�����K��	7�.�/���xgZ܎���i(�r��x��靯6Y'�	��@7���(���圣��j~�WA׹9��e�1��i�ٍL8�7x�н�Ɇ���G�ܲY�@jq��V�A�zK!i�\H;Y3to\�-�uz���?�G�Z=f��wV"�.k����"TC"�~K���P�J0xg�#�`�\���`tﲀa�fH��X`�®�k\z�F�t����'g��A}�����-�������󐕰��,�]�[dtv:b�ԋc���K�}w��ڛ�!��O�����3�^p{ڰm��O���$����?���5����f��̥�8�*�v���=
�R�(D+ւs�������i+m�-ab��Ҹ������Q��JN��M���S�ɠ#t)&f�u����W�R���!���o�5����O-RV���~?[�J��S�X�=�����'l�ڨV^P�ե¥&F�4�]��
x���nmh���3���$ı�E ����ƾy�S>�"3�n�D�a���8Ʒ�Mzo5��u�^����aZ�54j ]�u��;�I��/�m �r��AL���>Jǖ�O�7��b?���pw�@��r���*��D#��'$�p�Q�S'������� �����O�6��̐�h��q���#I�z^��;�J�|<ٕ�OhQW��5��g�#��1�Zc�#�scT�9�����e�ad�k�n�Lʽ�|���v�M)hHk_F����j��I�b�$V)_�ڋ�.E�m5��]V��*�\��o[	���v�_��~��I/N��UΗ�9�z�rs|o�7t����n��>~T2��B�`_�p����<:Gs�X�^���Tv}_;���7��j\�G*'�yߴ���l_�y��ݐ��3�#=S��W�q4۴������Y�㛔�b}�M��}={a�[�A2��]L�;b��L��}��J '���FE�1�/��|�(���/@��{��޷�����1z��� \H:�5`���d���"
iM�Q�N.N�p*j�qs��Bt���o�����3�JE�~ɂ��u	���r��h���8���
����(dw{thU�Z�}�ý:�_�B-3H+��< �t*�����}_�*��xo~?�n���}ˤ܂�U��͛FΠB>�%m��޷M�u��H�``Ь���`����nw1����H���N�l�۾���P�/���pgm����$¼��#�_�5��r��Q2���f�)�Tg�gȇ��@�멸̣���1>k���E%Fx�������n��'��= >'f�xL#�%mݲz�Ғ�<��l�@��t���7��9f�|�/���5批H���_؈�L��})������)v0���m�d���}�D�x���_�?K�'��l��y	��.����f{��"�s�|��D��3�? �j��x9����l�N��S��.!+(,HQ���*fى.���2nŚ����^�.��i	1ͻ��\�l~"fn������KX��a�P����K!��&�����dq���*7��Qo��6mbi�,����F��qHy	��V^�}̧KI_��淑 k�=�/3���3�H<�Me�c��1�S����P�������i ��<H�Ѱ�C��k��V��?��y�R�����DrV�C�y�� �@N�鸌pm�5���(!Z�!�x��X+W�6��I;��Ƚ�MO��N�d����y*�	��u7��F�4Kol:��HQ�"��xPv�9f5��ַ�I��� k��=BѳD��?QX�R0īc}�=Q"�	��x��~�粠*���W�#LCۮ��6�䖵�>4����N�f)�%7�������� `". �h�1[��á����n?P/b�DPl�}�D�0�)}�$���S^�[��j��o>n��g��0��w]���e�_{���ܵ[϶<�ݢh���}��(.FiL����_�T��u �����=d%_��O#5�6*]�*Q�\r\��[��� h��
�?���k� �L���2��0���1�aw?�+�qd^:i�������G�N���8�S�T�Ƴ.X/��������1	�h�iuJ�˘�1�9�F�H�5�i�>-3�d١ �O��UK�0�������{p���6e��đ�6qo�q�z�Օ��Pǹ0�v٧ˠ�ڍɫ��et|j��>f:T�0� xm�����U�=:�4YNtxC�9��ޑ��nH\`�@�MFџ�~�G�|��7�N��Qi0;���hE���*2�iiٷ���c�����v��^�i a����[`�����"9�E�?�U��7՛���%h5
�R�5<�\L5���f>��n���1����n��d4Y������E?�����0�v|*�1�gB4T��[�m�W�^��uT8;i뉪����Y�,����U�ga���	��b���I�>�f��V��F��?��x���As��!�+��'��)�h���%���8Y��]0d����哃��z0���Xr������zyV�ˉ���/1��	�/+�4�b��/M ��I5��J�v�Tm�9ӷ���W1�&&Nv�߀ՉM����ͩ�W���4P0-��&�Şm������z#��+���*�v���S���`P��wp���N��11IT*͡}�rYt��o�3	t�o����9G���4���qP4���ew����[z	Yl��l��6��d��=J��6�~h/�&��;'c��8G�~O9����5��A�s�GKְ>7{�8M�m�X��:l���&`���O?�����2�v��*M?�6�+�yLvG\�iH�2/���nI�z� ��.^ߡ5xSx��5R��a֣�4����㡥?�|ʚ��N���*(.�P�RQ�hcaNh��e]H~i�S"�>7Z�+�vr��Q@��q�aH�����V/�+���٧ev
ٶ2�=�j���P����m�S�6W�252����YSDc�Z�Sҋ��4��63���-jt�(I�U����u�@�:3g���@1>9
�1�nz;D�#�=b�__wh�f^;�;%q��z*n�����ъ��c�Yk^>�x���&�* ֥_ܑ�<��ǒ�>�?�A:f2�;�}��֑��U7x���#7�>�z�^=C{㡢Fd :1�2�p���(�T�U'�)��3'SBt<��6�#Y�,�@+j�)��٧-���@:�c@�(}̜�1}��'Y�	��!I�vѨ���_L:|!R�mW3bIw/ nJ�zw�\X׸H:�Љ�xk������\������5bh��^��F�2-�Q}�o*��![�F~�,��;	��ߧ���>I�`�b��86,Sw�^+���QBs����E��|p_��u?D0�ޒq�c�|�����A�v��;�`���o��T�����<������g��ēxvj'�==Ċ�w���'�x#!r�����dK}P��9BsU�;�R��ћ,��e��78���/y%�C�:����}����&��G�s��=�g+���9Hx���B��[���VKfg���!�
KK� ;ԳT�?��;G�6�.C��F�ۏV�n*�=4�s~ y��ǟ��U��v�a�ة�h���B�y�.;�����:�ՆjT����h���-�j�h��_�����$¤ޔ8��ǋx���VK���%���f��|���?F[T����T�b��o��eL�r�,$�����1����a�T�Zz0TW2{�7αȘAx'�K���jH�Fh��t�yR�H4PT�����Ⱥ0����3�9�3ǖ��52��� ����`9Z8i��m+k=>CWN�	�˪Y@�WD�ڣ�L���
n���A%r��:��C��Sd~u//H���W�����|�
��_�p��Ev�����268��4m��[n�[�m��У���D�Bˣ�͢�u�\�=W}�jzs�R4e���w�`��.Cn��S�m�=��	�o�M˄T��������N�.���U�C��q��4���˾���o�F��b�sl9�:аoL�iW+X��S�hn_�&��:�cK�
�g�k�9��~�vA����������=̰x���<�栅��f�ߩ��=�c��3 j��+h�k�YFR�f�����]P��;�.M3��fA�����3-_�m~��ى�:; �8z���YR��OA�P=9L��`��G�m<Uy�N�34ǑdBq�R����`�ÄuH��&���r���QJ(�B��B�+�:ҭ7h�J�����%����v��U��:�����4* ĩAD5?����k������ocv�Y�!j���Z;�/+A�E����Z�F���$ڍ7��
l���j?���l��cd6�����%�Hz��W�}Je�K7�)ۻ��h��p���Q�7͌�:�=������+��˫d�b�;��P��bPl�^��~���LM҅f��B �B�#�
�{lݷ�@t@���I��Xж�1L���j�~�D�l[.�-c�n�y	��h��n��DW:;O��߬�6=�������5��*�k&I����1�:R@��fPB�6��5Q��u�&J��r�yA�j��M�A������ܰ�sZ�|)X�c�R$��(�\{Q���9���M��UM5J��u�t>��jk�.*���ikEh8l,���>h�� �����Ư��?��X\�'5'6�ɗ�k�fĤ(jM�9����I����~���u���eVnlK�i績2x�=��PǊ��]���P7��L��=P�̽����[�W^O�ȩI�K2��x����g�d�EQ����T��X-9��{/(z��Q����<
���J� FW�ˏlA����q"W�c �_����)�l���BJO\�-��^խH'-�d�'�JRk�T�2����K�SAx�YLQ���nD~{Iim��{b��+�S3	Dҍ�9`3�9�������.�ـ9r'��oX�� r��'S�b�#U_ �U�y?cp����Z�@�	4XDV�}��7��_ٺ�����6��r�:�B�9bj���x����M�u��	��V�*c����"�H�e���42����`�`�S�t2m]fߓh��&�i�V�>)�vw�Բ��x�$qV˜��bK���.�X`�d�Ľc�c��[|R���Fr4�ײ}L�Kk�@���6�g	�[a�0���-ٔ�������U}y	��_Q���%�j���	ʱ��"���DZy��Q:X�������E�3�#���^?���iU�6�⫃nh�=hL�{Z�b2��{
������(���;�{`��,ˊ�v�..���U�6��Ŀχ#�Hj�Ow�x��� ��e=ʱ�9�C�GJ��m�Z'�J���$�d�HW�Y�V� ך�֏�{�ڦTg2Fg�y�㎉�="���A4t{w�0�%���AW5�+ܤ���"�H�}}3󦴫W~�A�eɎ��P���܉Z���6{�r@����k稤��p��K	ͩ�#^,I˭1ş�Ơ�^��s�m�b����X��ʄ������zB)P�K/����6��~j���B�����]�zt�ͺSV8TA�5�!tJ\+�A�J�t�xU�C�)	d�wg�"{�7H-�s,g��m��m�o�>A�����3�t4�ɰv ��e�bg	e� V��6�^ΐ�#�
��&>�'�Y��C5�-�Z7�o����a��p�UMS�Gvm�B����vi�mt�3�>�},�ʣ ?��w(�?ۊ~^F�-x�5/G>	!�Nzࠅ�)'M*e��:��^�g��Vj+gXA*��cs�鸐����\Ӥk�$i�g��l� ��9�޳/�ԏ�䈶mg�#�՟A&�u�V�ɴ�:�e� �=���j�紪1)t���I�h�ٳ���� �*�'	c]���;��A�f�Ő��6Lcڛ�69�g��mI��� �ж�Ϡ���Tj�}H�o�Y�.XsUE�����'?�*�p�"��M#��yTsA�]g���dS�;^��1�l**�J�%�n��A?�ߋ&V3�<ܰNDi#Ó����Y$P4�f�F9���ܛ�;8�
|��T�Vpͣ�Lٕ[��?�o�ģB���^^��ۣ��+��߅��i7G��0���<_��<6����_��sԒ�W��ܑ��s�u;�a�)�m�HT���S�4$F��ע@	W.�O�Ԏ/m�ͨ����q������a��tGj�zv�U�z��eL�k�:�m��-Ff�b�"b-w"p4,���ٴJ���R���%����SÁT�AY}��c��>T��*��m�
¼�C�x�Ö����ۻ����/ψ��n�Km@`�4i3\ޓ�؟zq~O��s��2j-5�V����V�Vf�� �Fw������3
�^c�g-8s�fgJ�%BT���.Uk�c�)��nC��g�������=�j�m�ĐPƝ���H�@�����:YJ>7Px'DIW�>�n�J��ﭢ@���ky��k`���c%��=%��mL����H҅V-��	WB<��#m�:(Ɇ{�;\�	�"BFl�7�	z�s��Zc���:1T�<�����iE��"������u�bOW��e(V~خ�(�rm�s��%�Fl ��ޫ2���'3UțdeN|i�k��^#�.xߪs/u��=��br��-�h�o�%ҠI�8ܫ���B�"z��
n����fZ�&d����,�����`���YGFIl.M2�׉�����F[awK�N�L ������lm�	��}�c�7|b=k�y���Y�<��+��q��ϧ��	�T�"�Ƭm�k�<`mD�]�����z!���A�EL�d :}�<9�����\� ����b�H���·�E��n�V1�"�k����x��k���8b$�E�桾����P�D�Fs6����b�Ya�K�S$ݸ�5�p��3n�d��t9~��h�rISu���KS5�"R��������儽5!j�����:MbEȗ���H����qlˣZ���émAHmC	�dzW9cq�a�6���4���YٓhRj�X,T�bS �ㄋ?��!� 7��i�O�3G(���A��8�gF���U��5)���E&�|��g��O�:�ٗ�
���r튪��@)6���� {6�������UF�Ãu�Dn�ɼK����qų�G�#	��锥.N���[�ދ�S3՗R�H��|��<�jVl��wQK$q���Px��WLݪ6��3�<kK�Wo���_����\�k')��M��a�n��C��x��[C˨�)���w�R�q!��'%6,�ِ�ǖ�A�m����0��CqؕU�Jƕ�[���W���+=e��1Ꭵ��n��\:xX+���eR���ʠ�L�I���o-BY[b�#-��8y1��xH���A�m��ih3�H�� ����ܩPվ R.Ob�3����.Д#:ʣ����l��Ö���&	�D��{V��bٳ�5�R٥�����~!c�\	mM���r�q%	�$����C�)��T� �qTK��D�A�
%��QU̇a~��&��.�:�)����n�cX��Dd��@Qz"c�|ls �S�������e��[�w�`5�R&,�Ēq�5�B���E|2�Z�u���X���CH� gg>=�~J��FO_�"B�7*J7fy�x~�[7�Z2����6�H�7���s��v�����̒TF�M2���RU��*��;9B�P+��Y�C�|oS���q�D��7z7�hU;���3��-��(��]gmנ6���"?Z�=B�DňdJ������"H�i�ߗ�vb���h�@,S��D�(�]�ǣ������m
.�v�Ѩ����<�0L�d�K	�42 �t�a0�5h!�����F6e��!W�<2�&?�+�^����GθUI`����n� :W������y�M��^B ��]���x�{#���kV�&7Y�;I���	ގ�k��-* ּ��Y�D(�e6q���@�;e�V�Ti]�"�|S0|L��
�7g�K�2�:�$�=�E=�L+ '���K���A�ܕ�p2�
pI5��+��C�
�g؂N|zR����d|��4Y�W�B��8��5���Cy ʾA-�X߰	�M�	8$ ފ�����3�U�]�	d2H��\q���R��R�D�0�hq)ѧF����J`Y<���%d`��C��]o�K�@c��`´r�H˨1,P�W�~	��W6~���v.N�(s��9k����KR�_R�u9�\Ȉr�t��F&6>+��y�+7�D���
2߆���ϊĻ�����������T$��a�&BE漄�nz�J���3P�v	!��b ط��r��նs�1�#,�
n���"%�	k��9��@BC?C�*�x�gֺ�h��+H����t�p��-\X�"�Ś�B�M����H��R����������l���1*8rԔ\>9��3:�V�t���ݒ���fB�>ڥ'�!���'"�>�pG��n����h����K��-*��(��2����r��3g(�7p������{�Ŝ��O��3�k�'x,���"��lw�"Å2;ph/L���U-d�\�#�tJ ;~�(��f���b�o�	2:�m���#��$����xϳ0��4��rgcа�8`�D��&���ϋ��the�A��A��a�_I|x?;n�q��,Ҕ�^��.�g��h���\>!w�LH���Ȗ���a�mž�0�e>C(/<[���,Fx􈡜��4z�E�s��2@4�xj��}�&78R�^{j߾g"5r���׊��g�u6X���P�2����M�i�J��q �����yO)����p"�<wf&|�'$4i�����H<"H��; ��3)����>̃��(WUz��T�leKqN1z���.E w�}��um�gU������D�⮅���%`�ad�~����<fJ�*�	O�OfH�ٶסٷ�t��~i@U'+YS�Jьg�e�`��q��Iǀ>265�[m�>�X{u	�<�ʧm��y�Cz���s8�K#Y�>=%V-P���=+�����V��,�\�Хt�2�������|W~���Ж�,��M���AFt���)�(�����?h�b�?��ף��`��c��<-��h�Q�E@63�N�a�Gۨr�R%��Gm}���wGW�Q�e���-2��k L������)Y#@��eˣkm2�Ӣ<1�
Ɉ�:�X�e���ٕ���Q5�X��&�K��Λ�I���s��w����#���d�t�IG�(�J9�I���h�z�����IXU
.h��JM��}L�3n3I�:�+Ì�rB�_�	�ϓ��'���K�t���"RC]��V�I����%F%�����M��!͢�\}i���0h����/�#�a���������BFh�C6�z~�St��~u���F�w��E���	:�Oŏ�-��s�N#�}�����o&���"����r@�bq"9�KG�ϩ�j�b��[����������U�����m��=Ww|�M.��ڽ*a0�h�זۍHN�����o�Ʋ�N�Р"�B� =I��4��v�2Z]2g�|�y=�eE��P~k���4Qfi}� a�G�Pk�3�YvKQ�� �M�q.w�v"��� �l+#��N�����]�{���hg1� �a��|�=!9�۹b��r43�Q"�x^@��fa A
_��6;�~6��dʰ�Y��⍣a�7%�c����7�F��NE	y�?g��.X'wz��n�V8ښ�?�Kkh�LY������'��lB.Lέ��UAԯ�a�S_kܓ4�UD����Ű�KK1.ɢ{� �S�~i%oJ�� c|�!U���^�J���(�`��׊�}�w�p=͕�׳��C6:؀���C>�=�� 〶kr�����,O��X"ո����z0��ʦ���?`{g����Hf�i���o$��0�A2���
�#���	h�U�l�!�����
����.���EQgы���ͣ4�~���k�A��[�
���D_��EkYH��,Z�n��ޫj���L&� ��o��T"?�T��e1�.���t�n�b���g����
N�B�;�yk�)�x.�Nߞ�\��2��&�H[�U-�^�&3$kn�U� �?c��w�/M�]��uV\�<W$�E
Ä��Ղ!�5p(X�US�nYw���Z�G�>�ZR���n]@n��&j���d'�Z�`�<y�p{FW���y�b�Tͦq����mmz��e�kD!�U�O�s��vM��@��j��M��Џ���C%S���"��\���l��6�����LG|.yt�ۏܦ9�*�G�:��E����S��/}M��V���R�vh�nKS���#�)@jq���9{�O�J=�5�g�^{H�5�a�a�+�TU� .��L�Nr�w/���a���	֐�ڻF������"HT�Djk6��R"|��/��j�(��c�	C�oX����M�m����Qqq˼y
遏�w���|*�����(�H6\n��(}�"w���l��Y�K��M+̟r/�y�LŶ�R�c�������8�
S~=����/^^u�h���`�����{
��l8A���͵Z�
b L��ƫٹW��1��wuoYAW-����Ԥ��2b��;(nr����4�ϙBM��Yy�0�ᅟ,��p
qbė�_�;-U v�"��'_XtJ�;j��� ���H#�0P�v�E����X�����t�pX8�yf�9�pnħ���lرAšeU���h�xx���?@���\|����#����ʿ�0���y�ֵ��c�骛�c0�f��+�b�;y?_"b����#W�-	�Pg��He�<����E�8RQ�Ei=/�bg�jl�۱�0y�.l��D�d�������|'��zІp�F�N��侹gӐ�����3�,����r�I���I���� �O��pB��rT�� ����7�N�M)��p���@X���B�ĂOޒ\t�K�0'��	�b�=$�J����'�(3>����"I6�;�qd�nY�7��^�Y<T�ɂ��7@��"��l�**���,�Ef��b �[(K�)����Fm��5�a,��^?����m�Q8"��|��d��I�^&/�2S#I`�kɃI-��Pw/�5�,z�S>���<�%�L-���Y�S�?e���a {���t�D%�膎�Q�܁�w�Ɔ.��4<l��fK%�`�m��}�_�{^1%:YW:i��E��r]x�Z"�t�׹V�zn>sj�e��l��&EO��7ק�o�
�Y�p�w�������.s�.J�f�B{Mڴא�:�U�Z���@�a~��mZ�9FhO��_��G��iӦ5���f�#=y�;v;��'ep�}�J�%[��j�zbi�b�4����3�o�Auܶ�����5�~Sy�zq6�^/唵����*���_�.G�B��j����"���I7:�u��Ew�.�h���b�n��wc��&�[3K�T���my0�^Cő�I}��V���E���#�[I�^�8&ȱ%���\�3FC�%-���v�GPЕf��N?�ƫ����Jrݫ�Y4)+���BY/\b2@��c͉�&XV�@�>����'v���F���Ke<^f��֓��1�K�ޭ&�w~'\��r~9䋔߷��I���F��6�c)�TZ�C1�r j�2����Ө���b���UT!���q+��gG��ݔ��Z�rq�+ۉ{�5�f2^x$����ϊa	{�Y^�E@����V�B�_-���o��0�JWm�S8;�j��d_�-��ž���=��ND�h%C���w�#ɢ%��n@E�H��Ч��%(�������~[&`P��������&!�ڌ�l�G?�B�"ң���u�A{��ʗ7/�$�5�����D�V��;�궃�zg��L��=^P��g�+M�?��F4�G�V^<a1���ұ���oX�黻q
H�>���*���*lr���g�$r7���{3���fX�Z�II}xs���?W���`o/?t����C���~�İ�u��u��E���V.5Ԟ�j��b�v_ҵ6Q7k�=��5�D}��C��r�"]��p��A>w���!�W��\���U{aZe�ft�A��ѰD�s�7�����	�=<�l;ك2@�Z�
��fG�z�@ӱV�:��4�}��S3UW�� �]�!s-�ܚ���gՓ����@�����B����R���l|�̛�{�OO�31�3{����P2�1]q ���g�9:Bg�(
oW:�19!˽HB��|�7�/pB��я�)M��������|�A�%Vq|V�׽����*���Y:�e�^j����+��C½2췹R��H���k޿�],�-[%6k�|.Nh��8�-	��gms�r���[jr�Y�:�v�$AX���Abl���G,ӮMd��NHO�M6Z���+����V�>a?  }��%u�ү��ן�|+�DU�Icsj�ljI;"xA��z��w�&=oW�Ǆ��Z�A�9tk��X�q5�)�;�}7p�����v�Ċ��4l"ڸR>�-ݼZ�<�	=!�$(9U��D����e�&lVB���*4@�I����x�R�E�c�����;@tO=ōp<Ŀڴex���6�n�n�iw���	�nЅ��͉�!��  a�3����È�cԟZ楧�ce�=��veG�*)�&�L���+�J��z�j�3��N�J��i�����p���r��*obhP�V��5�c�Z8�4�%�#�P��A�KW�2(`[N���we�t��<��I/n���!�%�ɃFV=N!Y�E�b�0���DS5�P���k��a�c�d���إ@z���7n�����=�$�׳�-�@����2\����5r��k�:�s'�`�I�Sh�9�[]�?'��-X�!�;)��CW��P��G���1��oS�||"��w���%��i�
���,6X�^���NL�5��	��6w`��6���0	�=�aٰ��g��i�r�����}�N�.�̷j�1 �S���jdԡt����Y���ʢ��[:�a�t��1ԞJ��}�i96Gyrh>{B��p�X�Y���Cߠ��¾#Nr+�0z�X�$� �)�V���zv(����Y�;��tX�%
�I*;�Z���\���CB�8}C���,�-	�m>>��)�wkqq��o�W���wY�z)��H�11j�n�Bx���Z�%��d��.,Rh��$��	9�B��pd*M~O����JѱʊOL<x�+����t�F�Ջ���C��x�D�zR�:�7��r��k/�$�W-���Nu.�Зr�X���H}p���Nh	Y���x��P����e���`Ql��M(݄^>�n��}��u����[�@R�<�  #�:��}�G��b(圴���x�]7� Ƨ��!>�`D`�tfU�xO�����q��"n��������Y�AW��k�~"�t���bIdQ�
���>Lо��Tg���L W�)��%��
�!�UX�"�k�55O��I���c��h�E����V�<���B�l����_�,���unϫ�cU�J�!�-1�hO7���h,ty����e��6�JAU����W<�0��!N$�4��m
�T<s+3�A؉3�^Aё�i�j|��1�oH�(��JFv�U�|����ϗ�>z���#oQ�{�cE���G�E�$� �dSIѓ"��I.w��4��X��O$�cJ�g.��Ne�h��]�'.![�쎅�o܀^�-/��棙�T1%Yײ�K|[��j�D��)�f�N~~t�Ŧ�{��g8R߿X�b�Ϟe,W����M�nm�(��c6ͦ�=q���V�	,�wZ�&C
U�#\�{�9��>�Ԩ�!��l�˧d�꺜�.��Bՙ�2�]�?3�Qa\6L��~��T�	����֌{EH���n�R�16��@N�����u���6��mW�M5'���#�Y(�\�ܸ�K��`vj�#�� 0d<J�IF�p ���f=[!�K}K�E�c��{�|���f�~ď����G�R�V��-�H1hr/�D�|D����q{����NC�����e*�Mx9G^�0���0��wi�� *
	��F.�ڧ&�lIb6q.$X��J4h��ܠ����G=�d�:x��ī�e�S㊮���օ�s���vMi˹�6I��b��!��_�ڵ,�����������b��ӟc�I����MH8�� �v��m���ނ٧{��Y�v/�:hp��s�ĭ�$�J=G��U� o���5�4�R�R	G](|����$�cJd������6[�V���ƱU���r-0ݩ��r�6�T]�`F�ga^&��P!5�v!}�+KʠRQ�^����Ov�+qts�ʑ����b0�A��!t�&��v�@��^.��a*?�D����v��?O�z�jS��M5É#����j�ה�*��AH9?L��w~��鮙�,i��k`2�)A�]@϶^˒�7`JuQ� �=��� �N�)�^�>�hWQwu�)������9���2^O�����ۏ�0C�y��--<c��{Z��/-�_��J��U�P�|]C���.�g; 8��݄�����j:>�ɏVˢ�����0'fq!���x���~>���|����Ŕ�˥��`���A7|��z59�fQ��c��t���m�������A�j��~%󭹫����[������"HJ��	4����z�JIeo������a<�|�}�sǩ�{4�H%�\E��rcr�%��ۢ�5J�П�]9�wq:��3���3��6et���S���p�F8D�e����!ȧ��Q��	n�g_'�ȶy�rV�{jP[�v���@ے�51>�-���v��ͱ��nO9U�F wכ�.w9G��>[\H����4�㿶���p�=e���=�����ъ��xS�⧎&t��4�h{YҒ6}���V�{E�D�}�4�;h��Q%5���yR�F������1t�d����A���낥��IZT�ʟK�8����P���H:-���Q+/j�Y���D\�5� m)���}�*��AT��<�gkIW�vmT��&�=K��`3ȉJ��?��֊=��������y5;��zoSQ�j2� ��j��@�)E~c=t�d |���yY��Ϙ�s��T���ৢtX9*��j �}���eo�֣����5�w���5|�c�p�9���N�qo�[qy����$�Zpf�8���'�<n��	&�Zb�F��&�����0}RY���:U~q����o�A?X���rA�5���O����Yƿ�q�B5T�m���r;'ЗQ�T�I)��.C,�~?�i���:ڋ�-�ѯ����
%��|a�0S�Ϫpie/L��I����+�s����1y�G�Yʠ/�SlCB]�U�^7��U�n�a��C}Ȫ
Bƞ��R�j��@ʉ/�@dQ���t8������8g3�آuחjf�M�S_��z%� j��y����K��On
�^�菪!XM�~څ��p�	{}h�!�7gʳR#���_dW�u?�-F<&:���a@R�!!o��-�NKsX�l��p3�r�~k��m{�+)n3:D�J��
#����v-�kT��!�P�n�FW�I�a��9%�t��_::��mg�D{<'�o�v���a[=қ����
�S����44��u��fh�gypoF]������V��uu+�#���Ox�QJ��{L�6Q y� ��r�.靓Z�T����6�E`l�ܟ�}t����IQ�W��U�V��>�_Wo�V���r��w?����jd��H��3�Ԫ�%�8����]�ڃZ+u��
 ���,p��9"�'	��d���W��Y���Ӝ -;�s;�(����[�~���ܕ~���W����Hw��tb��������]��T�FӔ��ឲ����R�Bڶ,;��]�ҽ�vq^ӷMΨ����"��~t��O�}\(h~��M�)Ef#�[��mm�e׀��l5�{����v��o�'�u�Z!�8�H`�� M�O�Ѫ��~�,�wh��=�(`D��4���Dϡ�pS��68''�[�U)���FV����7�����rx�IiB���h�Uz}(l�R^�g��V�rlN}�(KFד� @��\z��h�`�8#���w#0����w
�c���I����uI�򊞃)4zį�X��Az��6F��Y��A^Ef����-�y�����\��w�S��ؾA�5�l1GR ^�%`\����e3�j��G�PH�+�
ū��z�Z���
�I3���7��N��F~�M������(��D7=9�(��Bț@�m �z��M�F���\�"��a������G�s5�
s�zǉ�^�޹�%u���e��U;�[�cڽ��Z���2Jփ��5��8y��o`*�[,�D�.�d�ub���Y��v�On%W�֛���mg�X��8�C���nXۨ��d������$�k�9�O�.v�uX� ��+q���C>:�F�!��������^���	g��H4>3������3%�z�CP]�-ҕ` ���S: N
E�����8�ěM�՞J�P�.um�<W��c���������y�㞻wK���� � G�9O8M�M�dN�@��C���׺NT{��f�f"�̱�N{�9t��mCʍ7u7���qX��ʿ����̮��3K��4��g��kWΚVn����+��9��,���t����R)~Al�2,j�1�-�>�0
`�d.����ǁyi:d���J�"�{�Dw�w�v���M�lز0X>�GS��^a�?Bn�N�e���{����R��	�o����Y�;��d�%�7���{��?�J�h��;;��zN-{8K��1.�*�	8\(� ̿�Qźo(g����pS�TJ٨Ѥ�-h Kd��Ͳ����S&:!���9�%G�?��W2
���,dq���;��{��cؿ��
*M�ͤN���׺��N���&QcN��=�+���4��E��eva0Sj>=�)�����$/3t�VCq��<F�1�h�/'}\�u�X�����?g���T���L�� �%��ق7���G{�s*���PL����_�C�R�$]΃�k���/��'�D'9���ٖW8��\a*���;{�
������6��^��t
�x�l�s��e���k&R��)��������
U����r��,Z&_�(x��y[�f���^�R͟ӽ�m�f�5l��>������!V�.��M*N��LPF��˴�t�jv��Fs�!
�{�����E�Ĳ���_0'Q���>� =Xx�� �T�L�����)�6��RM�i��4�a�vG�	 z�9F<X�>L����hn��S��`��L�ڠ��W'~nr �vRR�1�0H��,�����>�Ύ�]�`�C\/��,��*�@P0ۻ?��X����O�)���Y�ԏ@e��#8blh"�����4xeE�]�-����@Џ.˰%���bΣ�(Ǖy|����>�F���˾^�v����;�6&hsOH:N�Xg���_��BGR4=-�D3ׇXx!�<��8����}?�4����پO]���Gd)�.�s���&2Dcn�8!V�	K_2/�X/9�\��1cyN�B8AB�,$����c�fK1*�x��4!Ll�Q��;⠃M��Y��և|���:�X�����I3H�����*:_�=4=�t_Ɇ���/�W��|�b��68�U�sѰ���s�|��K� ��� Np�OpbaQ�9_��	\�8v���UB!������:�<|�H,�u��Qd_��W�T�Q�ު��?��^���`MWx`����ǜ�� w**��Ř~K��]��|�yA�N�P��wR(G�d���r����Z�< �}EfK�(h�b����G+�;QDc�ۆ�QmT׸	Y�4p��=@C?�|ٮ��b��q4�Eg	cH��ɫM�0�JnyH��n� ���� m9�G3R�V��z�zt���!沊��Ĵ?$�G��	���F5�N����,��zW���@~B�n'�� ��*7�ޑ�� V��J¦
`sc��Z�=~��ʜb���Q�ó�����~�g�^�;�5��*(OA���!o�h^A�va�Y���FIe�#׀�(f��0K� ��`���Z�&��Z�q�r^���@�~y�Ӣ�)���a�+`��8x
*�^�_`�2G��#}��DWw[mrGT�r���J�38�am�g���|�rD�=�$xfB�;�(U֐ �V���>tx��P��+��˥0R��&=ofs]DĚ^dEVhЊ?L�����ƾ��Vq2��vc���@���6���w�ѣ���Qt���*`H�rO�;1��hS�>�m��љ�J���p�Gq�3�D*�ϯ�k��Ϣ���
��1��?26nx�bTrKz�)*oZ/��������Z���-��/��{|�9���E��.R�,�7^��nJs��\s��S���s ����<81eqr�ډ�p����b�=Ժ76�y� "_�j#8�8tLE���r<��Fd�+Q�!ꪧ�ʇ��F�� be	����a��ہ��k��:�F�$�����&-ހZ��+�Y%������	�~��JQ�����1t� |�8��ݕ$��t�޻r/��/j����"��co��]3	�U(�,i��?БR0�"��2_����V))Q����w|�Y�����
F��[�b�VﴠWs1�~�/1Ⳗ�݀�\�����vR�/S��@Z��)�b_���AW�������|oB)�EtQg���f�e�X<�����IuJ+ K�U�P%e�;
�+	57����oA��om��Y��<�>m4�Hğ����B�y�Ke7t����=��㊞�)�}H;��4����v�f�{��G�E���Qz��斟�u�%Q(1&�qn�d�x������/����u%������Bm/d�(�����{�zadŋTI�papO�u؇غ��;N�$�wU�XTV+�0z��<���Sh�����G���U�Y֞�;�Z��n��B�#�
õ��",���3f�`���ǆ��g�`�M�&IaU/�����p3����0���_���V��9���/�nN�T��7!r1�^lL�RsˍonӢ20E�	/;�r#��Z��Xī|U
���?�[+³	ig`2{���K8��հ�3���:����=��W�ό��=@�RT��TBB!���H��	�t���Zf�3H��N,�0񇺎�m�	�LW�E}<�O���pD�\*��>��d�~�q�%[|fօB���CҴ09�!IL�+�	������a�9%� �S���>�?�|A������C�a+�t��C�[B e9(&!�P�e8������ڗ*2E����[�5�;e�Y��ɰ�@A�b�Z��G�ZSEQs�Q=��>����uѝ�QC���ϓ0V;���U�.�r�>
a�P־"'���N}"D������z��+c{�i���ʹ���1��d�=]�t�E ��YQ�2aa P���Z|?(��s�M|��:�2R+A�06Î��y�_���d�#�D��I�Q^�C#��,Dw�� ��,^j�6;�P�2���"\S�p���%�7E�A!�4י2̒pM`�O/5�7�}`+���.��)O|!���)"b����zD�E2A����J�Yu�fD�@LN�%kk�I�_,��SJy��q�gQ�Bÿ��FPHc���"Z�E%z�1�}q�9�"��϶0n�<N���e6���ѓܮ�o���=���]��NŬ_� /7v��c5����,�(�~2��J=Ӷc{�C�"@=�wm@�1� 7�W�㦮wzm�n^�!���+�ʰ�]���_�F����5RvK��{��Z�{���7��h$�h-�/׻���n����h�H,�D��V47�k�O^��x�h�3B����
�Q%��Xh��
�pZX���Ҳ���� ���(ۂ��7���P��:���0�m�-�Q�f��ڲ���$��/	,'�'��[ �&-�þ��o���v�TΛ����L���:���H�u@���Vp@�\�l,�C��C����%�/��m��\xN�S¬kI�{�Ř��3℻~@Y0$�w�@��Z^�U�Hx�s#�����?D��Yx1��)��i�]14�!'+�(IL+��Vsg�{g��f��������*,�97%	�>e�W=����M	�
JN�%�p���0\9���v��a|�q�v��L.`O.��Mլ̹��K�&�^��e��.�3M���\	�<u�����N�[O�O��m�e�L0D��M:l��,�:%Y{aS�� Bq=4�VO�W��	���CG���e�"�2�1Hq�2�����т6�c��&"�L��U�����}�<y�r5��t''`���\=\���k6��9p�>)��-�g�V�;�5�ϴ�	���,o���U��!6侟-m�)�$L���'������T�ר��þ.A�-��J|��q��c�.1ϲG����:��fLbss�W?�ȓ�.�җ�x\�$w0�	���ˢ�E.���$Ŧd��D��':Vk�����$�r���X�i�ʣ=+%=p:Y�A0u�������$f,{��T��?y�׫'��֕�Г����$����,���ÿn`i	�f�i�v��"�I�y�u�Is���Iݲ��Ć����zS�
��A@OF��)����i+O���m}?؛{euX%�����,�P��r����)���;�.	E�F�g�O_Fo�i�D��?�������b@)�&G���[+0(��z?"�����Š�X��zB��[�c硓G{�tD�xok�A�=b����,���$�V�`�Rb[��5�A���L��5AR�-V�(g0>x9�!��W'��Tt��RUs��)Шx�A�ꁠ��/�I;�rq��0�
j�]�zdů�k�����(W𲟅��R%��,���7'��lh���͒��(u����s��2�9ډ'V�����dS��Wh͇X�)��A2s�*���� ^;$�d�Rs���Nl�]"�oz�x��U�#�Q�hF�t�����ZXl��1?`��K��1{� '?A��V�"�B�ʒ,VD5����p!���F���8��ꬾ�@{+e%��q��n�����RФg�X-9��6$FkCr�a����R��x�EC���J�gHS)yZ ��s��G0T���Ϛ~%�z?��}���@�R��U��ԉ���;�g�+�T�V�o�L�,3T�D�a�I��& ��z����"�H𑍙Eg�HqM; ����gZ���Nʟ�5t���e\4�%HC1��?μ
��~�o_�55�NSp��q	��-i����e�	�q ������E/�A������䉭��|5��[x��	٤�����nF���c���؜2�K��)�4W�+�&E��U�\�
<��#@�J�v���d"ܡ\���7�
�U�`i6 � ^���a�h��4��k��O�;oc�N��kg�>�s��<)��{�B�TM�ee��+�����RdHHt�k� �%�[�`]�����a��1H=.�}��gR5�jr�~���E�q0ƾ���l`�>P"��E�.��o(�����V�����1~V� �jP�Cw��u ��IoRy�rK��a����|K�F�E�+�F~|�_� ��&�(y�<
����檒_�p	�.*'���ׇm�� ��=���l�L`̴�3�l�g�o&�Xw��ӵY[Et���rK6��(�x�K�|)H:��j@�-����Q-��b��v<�����Y�5�Ԃ��v/(����Q��S0?
���m@�α���%����Vs?�}b��q|�92ȕ@*'g����x$q��:{������)1,�z
���5��_���o\�mF�H��m�p�Kv�-�|q.و���3K7���{8>��eu.�D�$��?U��"Uٖ %
S����vi�&����eЖ<�T�)s߈0rڙ�u����t&,Gvr��O�e��V4J����$�)�x��0D�A���&�m�>"��І�?h�Fo�hF�C�2�W8�RL?DZ�{�n������V�������ȵ��kaZ2��x������BX<z'=Qz�y';�m�@��t��v0\! ��֢p��-��fqs90Y+�;�5�e���x`	T�w��I��b�r�j�5�!.���=_^.���F��r������������(��8v��m}���jȆ�_)\>����g����/����O��F��o��~���,��Hv���5]+/\�)T|��p6+-�mG��`��Hy�R�����as���\d[�9]�v��C~D��RPՂML�`�Y�;U��k��Q#���_�5�����<l)/�Ӊg8A�]|ۯ���t)U֞�55.�l�A�i\��e2Tw�F���!g�3V�N@8� �bd�tb�,��j�dl�D�H"0`�R�g�)K�~Q!��ҥ�r�0X¨JR�x�0�QU0���<*6�y<!�������/��o~�N�p��1��G���v�+̄�<��W�][��Q���	g���ۼ�b�S������'и��$��r��nU�O���1_n�>#F����7�`�:�T� ��E��q�D����;�gPx".�9Ƙ�f�+�c���?g+w]�v���J�h2h~!��mq�~A� �1|�$_.I���S&���u����w5�I��<s3�A������!X�6Yߡ�&�
GE�>�S�ۭ�-�Nr�{$��b"���E��b�-t�d�^�C���o&{&l�*�B�
�
z��m�ӊ����̔n���s�x��������q�����9n
���z�n����n��I�=6Þ��G����6�����8dy]@�7�h�	�ٛ�&g��#�g�p�`��3��"'����N���|�Fm?��RX6�h�b֘}T.	9��� �i@(U���읨�L4;'���~�E��3ݼ#�I��� l��]��^r]���o��#��	k�*���a����Ȳ��*¢$H�uG�d8�u�,�`������%�����s��x��ڏ�4�
�PՒ_p�f�t��7����F�,'S�J5}�6ڱ�Og��'����:���S.�6�j8��(n�o��ٛ�s<����)>��ʃ�'-���x^�Bh9�l%�"7�UU�x&]��/�2�Pע���%d��8ʹ$�U�n�Z������ݿ�eV�Fn�� KCUY`�Q|�;��������%��O�6L���P�{*�O���A�Ǣ�(����< ��1�.X����ߏˁ�.�Vv��|�&A-c4{�E!$�$�_�t�l˲U��uZb����iw~	�$u���|s�z�=��f�F�;�-���Lv\�r˨�մ�Ϫ�ɤ��V�I�e��(��F����L�4O-���Jd���@�v�|���K;����������߳げ���r�B�Z	�'�VVk�P�ܗ�iHɮ�&"�8؋��k+z�*~�z[��e����y�	��R��􌊴����o�?u#o'�@��x��G���#��xd�G���=ʯ��N+� S�v�c�G��?)�%� ��MsrZ	ꋥA��D�j����V���*|�E]� 6�^}�0F��l)rK�ο�쓑��N���g�z!�8�DD8K?�W`�j�����7��%��*zi�HA�o�Y�zh֫�t#�y����X��@�aO�5���ӟ��;|u�mtE�2x0p^���	LuR�S7��\z��b�aiiA��pt��W�Z>��L��#J�
Ό $)����MY*�>=��
g]ij��avȵO��F� "�;�:B���U/�3/$��R&��V���[��V�VY)������=hy_1b��NP�����r~4�a���Zi�y�2%(���2^������hd��L~����K�L�׾U'��V�� <��>Xf��f�~�72R�k�ZW�lT�^4�!2���(.Y�嫽��N�+�M��~ݡ:�d���T|�񝜻��u:�%C�[�]�{��y��}�qktD�ns�?=��fk̘���[�@���,C.�ر�su��1�72E�Ľ�a��⿂̋Œ�b�yY��f�� �VM�N����}q�I�d����u��L{Cա�m���U�Ό���D�ŮkA�u���A���#�jW������$c�M(�f��i��QĨT.B�I!B���x��@i6��~_�ebyw�����l����$$�e�(�pW�+`��l�t�`}<s/� %�T'u��wI�<�l^��([{8/�L�3D����# ���g:fZq���Ҿ5��f�ӦD_���6.��:7��"X�Jڟ��ݴi|��D[�94(��=		���[y����>����E�Q����mɁ�8�W�p�ո���յ��a��p�Ff�Dؤ��	�uX�e��V�n��{'O�d� Db�ё�80���q�d���*�����%͊Z�t��>b�"AQ�G���w��uCt���%ya|�;(o�3g�����65��h=@�.�tqM�%5���Gּ�Lt[%�}caz���Ӓ�{������#�UV��\�"E2����"���>n�@�Z ^
:!�n58F�*������[pÓ�z#ƜZo_0���Ie�*_5�ۛ��)$���+�h�bN��?<������Ou����3��m��<E���u�#����:��?f�G�6E�}r9w31��ᖘ������s+M�)��O� 쟤*m�>�{t�} �;5�������9�	���^��2���^!�4���X%+@N����s�4�%"��ک�_qʭ�LF�f�d>y��Z϶3W��6hf�~���i$>Pž����2����� �@�S��i�&M������
3���O>D�@���Wm�rc3�]��C`(��>����l��7�\�$��G�GT_�����6�\m�.Չ���7׃�-�ɵ�u|�`��D� ���ܸn�*���,�^*�0t0�+<[��q���ݎy!D�m!r��9k�?�AfE�O����nA���Ur������g� ����Qb��l̑!ؔH��4#�Z�[�bv#@��X^��9P�+~���x}��r�F���s������
��}�r�L.��~�;ֹ�a�)M"S�M2�X	�<ڋ�`��ͨ
w�Fdʿ�F������Q:A�Ӓ�ԟ��m��H?uQm�܇9χ�Ak�_y4sG�   z�7T6�O�T�HQ�R6۸v����g0դ�=��B���A愌�Rd��ϸ���`��������=X�h}����K���	2��HDt]S*�a�c;�=�S��-8�-u���k����v�;�9�	�I+%T�X��|"NI�ҰG9y�ݹV���"�À�e��"O��S�43��Ȓ�S�]�K�m��ږ�'�h���:�R�<���^7F�Cf�"&q�}V��C!�Y�z�����GswL�5���4�Ӗ �=WLо�k�/!��X��qb����\����)��`Z�o��D�{95��vD��+��|�2x��+V-�c�t]ͬ5X���w�z4L������d��8q��o�6�;��h�a��  �\MS�I�L��-�����Q|�s�`�PG��ȍ��|�������s���2s�5l�Y�&5��ftQ�/E�P�"��@����\��z$EŞ�'%E�E3���F���<�c�j}���O� !��F�[�]�$������]�F����z_���(Ǖ�{�9��1�٫��+��G��r�*-��U�쫚
i�3T�0��X��ε>)��#'r����t��*���I����3��.�����Z�s�%�o0$���kuJK�w��|g�c��W��|ʏ�~�Ɂ�A��Y�δ2�������@KJ�����5<nIk�LJ!bԆv�h�`����a�f�_�~���=���yi�ğ/y̜/Y��Vb@ju�N$nQ�h︘��qZ���1����Iu����QB��#��ѕ����7�l��[#z}�zF���II��b-@HHWS�Cwg�G�8Q�x�w%8�<��A�0�̠���qHu�|��/{��*r��:/����'�_ᴯ�)���N�ҎT����^x )�,V�8��Q��x����� Ї��P������#��q�_H3�5�mKZ�m�@�T�*���l�k���b���9  y���;�6Y����`�ų,m�����pn��5��`�W$++��#�f��B�6�v�`�:�����P�ԟ�gy��hЎ�C�MR���Ϗ���9�UEhw�
 �me}��<+�PM�U�~���+-@Xp�z��� ���Q����hd�l�"�
ޔ��2�������kp>n��e�2��f��)f9�T��Ūz1�b�ymP*A{�d��݁N���
�Ȅu���
~Fe���3=>�M`����Ծ��=`\ͯN�Oǫ�������V��Y״�ˁiu�GcF�9�-����sC�;KZ������� r��X�k��'}� RIE�l�".$ߣ��Ss�������.�?{a�>�.8;�`�IV/q��ҭ.���˙�����Q}�%&�����n�=��w�\���SF�j���}7����F�P5��`�B�g�P����Į�AY�<��y�?���NN�}�]�Ny�g��V�NB�n�d���G��h�a��9p�U�l:���	``@��ԏ��uo:qN�Z&}��'\;��YG�<t�Em�,��4t��{�\q7n�tf�"KR��!� �0U,u�v,(�&�h7g�t�Ď�߳�%���A ��n���&��I�e��* ���tA+hZl���>nPyyP�tj�<j�i5Zq7�l�ޠ�*\��T����x�n%��p���-�����D�nw��Ƶ�t~��\L)�k��"�=V�pk��*�F��Y�(���ͤ3f;J�5e`�8`�d@葶�O�.X>�H�8�~��~ȧ\#�w7�Q0L�i=$�&�	�
���-�J�`�15j�ʿ��L�k���u�ϛu4���>�����ӌ?)/q�.��� e�o,m9$���v�C��r�[�,d�zT#��0Ł���6&�䴤Tn����X�����;�q��^�taֶ��=����X4zw>?�����D���4՗�����8Z�ĥI��u ���\���0���p�g�PǸbb�ݫ��vb��G�8��{,��;�4��;m�q��u���4��k�*�HݧX�(��:�G ;��~��`V���o]k��^�5�	����P@!c?6Y,�W�G�ŋ��W�����1&��0����Þ���#���k��ƪ�.<``�> �KԳ�f-���d�U`g����P��#ZPꀟ��k�
�,"Dj!�d�������� J��.�6Y>��#���]�ɄN(mzDh�P��?M��O���=&!��c����h�.+Vg���{!8��TvQ��ȝ��Y-2(Yl:#Z�����ʀ.*x����Nô�+�<�=u����9�� ~G�~3jQ�*sh�Pdf�Ϛ;e�����A �����Gl^}���5�#��B���%���/^��VRQ�Bۇ��	�--��|ƚ��<`�:!7�0����������*�AY0��\���.Ze)��K�L�0��L��E�$��-�	�
�H*�$��gZ{p�����Y&C���F*O��_�@� 
�C�p?Ha�qO��_|+$��z����� 00��P�{+
��OtU���>��m�f��O�R�Ġꕴrt��_�"&��Z1���Bǘ����m �Y/[��^嘛4k{چ�����-,P�}|��e[�S�ʮ�ȑq6Q�0zրvNK����E�5��|�I)6o�����'�nb�'o�v�`/����$�]ҜoX$]*�3�ظ3D����IJ�[ݵG���KB@{$*:h4 n�����㓑,���� �"ݼZ©r�@��7�C۹�%�NB���j9����K:6��xeN�RG���D�zÍ�IS)2p��}n��e	[��!Ssd?�Oq�Lm�$:��ho�ln�x�+ȆD��뤼nu������P0�*� T��T	���Q��]7T��!�ѥ��`�gP��Ζ�%a��*:�Wc�z1���[�6�)�v���,M��6TL͡H) 2�hr�y�GK)�O��Ƈ�׳1m� ����bu{P�QĀ�m���|���qǃ�j�j�iG!����"�x5f�^R����%W �A2�� ~!�x�R�v��L��"��*���j�%�IO��a�aI�c�>�i#b�9���26�����ސ���oZ�l5b�Wg�C1]S�s@�J��)Mw;F�Y��nwp�]x��>���߯��L:�#��0;��44�B`��H�����׵?�ן���LB��׌��p�a�Rl�7����.48��JsgA��.�������[���hQ�,^  0��S��2���6c��ֆ��B���5G�;���HB)�5慷�{+�c��<�P"0���G c ���\w;x�ŵ��h�k⇔�
CG��e���a� 7A����򔄁�j�V~���yuF������D�]�s���R�P�ڤoII��u�T, A[�a6���O�yL
�v2YA#Q�{X�^6�FubB��ǔ$Bx{Y6��\�O3�_����3����$r�#-E�z��-?�++�r���{_�0õ�!~6���d�"����>��bK�Y2�Z�r%o�y��7�
Ϳ	+��Ծ�Y����:1����U8q�]�DCw��s�vȿB⎚-�C�=�������đ9��&b������i����YD.s�~�BC��=�O_�H5�HK^���HnFA�I(PFwz�n������wr�_
㗶zF�[��W�=FF v�o07"�z!&�� )��\P�dl��r5�R)g����8�'�(M�:y���������[+�U��g�:ee�s�,��B�}�qP�ʹ-, �巿pɂ��*�G9J*VǢZ��wu�����@,Q�*��ɐ4�s��W�����9�'5u?��Q6B�m��~�8��$��2�%�G�e��5s(c2O����
�Й�tT��Q�S�4��-M���6
�>c��"Cl n/[R@h��#0xb�z�D�o���$��8,-���ɹQ#d ���1��O������Ǖ��$<Y�D.��ǢMev�Vf�c�ӟ�vD) �W�w�2X����b`ײ���$ɖ�u���S�X0?��^�Ro�Ä��	��G��Ֆ�%Ykd�u����X\���@=ZO�K�#u�(�͢S�|����	�pU��kv�Qꞿ�<?M�q�������"7�,{���Tk,Y���Zp?�զ��H�E=�B@��I|d�qg�(Jb��`�5��D�s%f�DT��7�x��l�����ԉ�2:���^~?x}&	1��M�,�D}���b���xv�p�z�֩�\M������S�ﮰ<���F�:,z�B�/��{����"��8�� �"^#r%dff
��y<*{��t�9Ã;�=$߳���[���N�'�Hѧ�N;G�%w8�@>Z^��W�=.�쭥�/�ì��.S�H,�%�ZoB{Q�E͂��i�Əf�d_�20�Cb	�N���-���z�m�F^���Z�:(_�w��:Q�혫?���ͅ0YC��~霯�r�� ���	���t�m�+�$��dF�S8"p�~J��?vz���V���lc)f�7���}A�S5
Q�	��� 8���i��5sU�N��Ѩf}8�B���w�xN�աfl"A8,�	l�`\�0�Y&\)nx5�J��1#��f�";d��S���l]��g�f-B��$�bA]��
#Q�d@����U��w(�S705�|���~6��`Sb�Z�F�P>�٣�� 1|����^�z�;�4�~I�,tb�.���}�^�,nEG0���;���F�0�?�e�x[,wn�5;m����`EAᨊ�$0#B4,��S2��8+�i� �e�F�H�Ŏ��I�K�����lٕ�q:\���F+��0��#9>�16�$�i�1�1"���k$�f8�t��!�b8�P��:.k�/G�i�y���Ħų�z\툷�U�|ͧ�����D��㉒K�X�´}�Y`K1.?�]���W�z
�ȓ2;���*�zeεE�ރ��r�d��z��Ad���ڽ�.��PЕ(���G�Ɇ��T����w��d���"0��Ʌ�G�K26���$�V����6�c�����dO�YΈs���-�ըrn�,�y��C��N�/�4#GT�"}g�$ا�TT9>?2	�h��Р�\sKRJ��Ha��R������F��t/���d
��_���H+B�3{�i�FX4���N_OH'�H��8���&�u)n$���Z����ذ�#�;�����v���-bR|r���P�}��f�@�`��ϥ�����V�~G�����sD�u��V��c�t�������/���	u��і'n�{/K(t��t>6}T��pJ�����@��o��s����ɔ���������׽�{#��P���a�:o�\�AY�����RZSn5�)������2�(��w�Kʦ���lU"og���_��?�,�f7���.3�7Ø���A�0�n ��mVDF��3�֪�&=���]ė+�K��
�A���V.�e�70��r�%�M��;\��e6|�[n')v�kE�ʉ��'���|��夠�n��o"�N[�L�.��>��c���"�����?�O~�z���1ZK��;K(l�\�9�n=H�f7O9�j;�j5�<)m��fr�4���Yg�pR���`���߅ ��i����y������q-l�Ia�d����orF�\Np�����%b��ٚ�%P���8;�n�Mٌ�lk��U��$�������J��:Ƚt��#2F���ء�E��>�-�e���Jx��Y�	��Ѹ�8%�5�%Ŷ{y���;؝\��Κ��2ӓ�	9�2��{Pj4V}������_ł`!��L��P��t�Z�P'*��c0 =���~���S�ͺ�C�؝������X6YD�_�*Q�/�Đ^���)��ND�[�r"H�q�����Q9��F�<���}@��[@)kn�˜���xc�62�|����hB�e�.G�	7Q�Iț!*�u#B L(n�r���,��@�C3}�t�d��Gx�4"H���Q��Y9�'�?��n<mu������<;� ���=d�c�:(�����"{gQK݄�IzE`��cۄ5ߺ���"X�"���Ќ?�f��P"�,�-wh~|���_9P���������"�K��ϭ�U� ��\.167�F�Kkh}<Vw-��������L�F�;�w�t{P�m`�Oi�W<�x�n��nk��i�9�:�+��żw���yA��%ଽ�Œ|��)�q	��,։:֘���G��ʤ�G��k� ��XԲ��s��MqY�pa-+3d, f����˯)B¡I�IC7y�:a7pF�0��z!�_܀��N��{�|%S==��jchfT�'Q%���y�"��j�� �~'>n�.J
�|�@���	˳"�}E�	d�-��ia�ڥR����`�a~�C����`F<ƀ4d^C8�:6`���� ��XG>��p��UV��H6W \���7�h�S�.�lY�E��_�r�x�T��txN�7�3����jTc���L,��~f6�Ѽ����9�;�y�/?���0|P�s#kӪ��*{ ��8]�Q�a��������L�X?�Q�!�x�I�`ݫ[x֝ȿ{�M�_�?S1�w��!��G���_.��uy��xsٕq	�_�ڿ�� #�.���Ní� haa��c�],��`���%9|�Px��6�F7�����h g	
�å�_�ь�d��V��uTC�ƃ�_�
�g�:{�P�oz���*5_Wۦ�!`(t� ���/���=#�	B�����d̀�&�p��_}����SCc<	�9���[�i����7�%�˂ԟ�8ts"�b�?�w�y��F����Ȟ�#b�C����&k�vC�z���"�H�|�����2�y~����[�g�3�fSZI�G�����v��j����Y%���Y���YW�{�����('O�Zo�Jr�,/ sL_F��]w����� ���̧r�l����9=��Q��h틐6�^��x>�[@�9S��1�W(b��h(�A����3H�dH`�h�`,p����$�|^��	�Kd��\"uv-*y�v*�Ŋ!6�8Pbb�e�%��6�7�<�j�̜0">z�z�i[6d�L�֓0��Ϫ�c-��b5?�G�:�#!/����2����jh<t��[Q �M_���j�Ҿ��@bn��*�_0� ��j7K�ɸ\˪Z�������%��8 �@�౛�j?G<h~�b��^��]d��>��_N��qX�|S9�o|��}�q��7�ۈ*�!	�l'���}Z�N�j�py���W�WpFL@.�O}����L/t�ϔ��s6��P�`XA�a'sEJb�u��\��5���H�.G�Ic�&���6����~���IF\ݜ[�ߧ�[`\�23�b[kq�*���D� ���=%4R�M@�^�z���Â��sS�H�����yLbA� ��� n�oЏ�1pfP�|�'�{-R � ��|�B��N����^��<W�e
F�2���7�c��u�m}�-"}�SS�N]���V�[��fc+T�J�H*��!�n�In'����y��uX8�S%{��HDߍ���{���H]���\��&�B�&�M���� ��M����;��2�O��CW;LD�5j�u���
��N���I��o������8������������,*|SN�ۂ��C\_M[���
L��N"s�Ӗ�j���ͥ�	b��0&��뛍�k�֟���'���̫ ����u�H� 4��5�4���y�k�@��Z
�l,.�PiԳ^`h�I+�ԟa�E���J��{���x�_,��j<I���"6�A=�,ꯜ]���d�'�ؘ��DU��	�^�N�0wa��u�s�[����VQ`�?��x�BCF����0�R�.�w���7�i/������� ������@��F�E-��<o�UH��P�Vq&7�$q������;�]sA@"�?؁3���_�U0�	��4��&��֏�������b�A�ңii\o�;5�x"*��_(���O����'�C�9���6�G�<�1y:�)x��պ�h��|K���?o[���Vڃ��{���k���]��bL
��f�q;���0�v�PU��'�����=B�!�����6��:���瘓 үuwԑ��M���k;m�f��"��O1��*���<�����T�:����P��r#��w͋ϝ�-�F*���X�x1�Dj���0@�8��Ej�+�AJ��w6�+���Z ��% �6smL�K6��Kf�C��k�m�I^p������U'�(wLƄ�Mkk'���s��9������`�I:�ߟ,�b
�,�ݎ˟��>��K�CT7^��t3�ќW,B�J�����/B����c��槛j!��ڟ��a��U=w�=�5��l�G��U������W�d?���?c�#-M�k��Q�BX���*up =	�I<b�%�lsDſ���Lek!:N�s+��Ԏ�T�E�W"\)$ �[&�rG�խ8��Bs�^D�{DjX�8+��p؏���6ՂN帷��N'Q'�(���{~�o(�9lh��=/̒s��&��qz~uo�)���شr��a���Y�I1N����V��x�wܵ��@	e"��ww���v<	�i�8�?i39��t�0��v,���w�S�0bL�+A�Y�_Ƚ ����J@����ڋ߰$�x�&_/(�xr�G���d�������H%)��)����(!��^�H��$�?0��C�����R�Q��8oi ����l�,�ִ�	�Jʐ�.�͹;����-ڮ� f}\x����x��(q;i�i�2�l�t #�%�%BsR+N^��eB����H�H�Cْ�g��c-Ѩ�
����|��E�ĳ:�܋-&QM�Gn�N��n�o�W��Q����t|��.y�~I�{&���O?��%��L�=P��}���3��9�G�09b�i䛢Ii���b��|��/t��XGF���cT�n�)k�����4�t��F#�4U�m���Vu���p`����(��S!��p�F���fÎY��8r�7?%�RӏS�^"����/4$i�Z�C��p k�"�v�(��_���3|�1��2FO#3+Dɇ
��^wAG&�`�iKY�ھ�pi��l�Ή7,��]$ޮI_���<[ͽ��X��%�T�w��]H~P7�1��5^����k���4'�ڎ��6n�E�#�e�ڳn`�#�ê��2�{^{j�C��S$�ݩ�T5�i��KR�57I�G$HWr4���|E;;]s�O�1p�E
�n<m��D{��ޣ��1D����/4*���#�J2����e�4���-�K��ڽ�����F��JR/��}���F�X*G��(ĝc�pP$Yz����[x���^�t7j����Id#�(�#�cue����2Ĕ&�^����a HE���}��,�j[uth�:̖G��P~N�p������f�?�B��f�^~�p�;Y��X�V�4�.�}е��؏���Mw��@c6L#LϨ�R
�K�q��8�mC�y8|r� �n�����̵_U��g�l����+1Pt�����-=���A�>~����!�V�0�_b�n��C��}{��	s�Fy#��5<�S]R'V?%S��BW^������F�d[0�K�n��*{��U]}���������=���dw=�Qt�]�B�=��Ǽ��}ߵ&ťD�L��u����+�;8�o���v:����[�U�AJ�إ1m�E��jE�6o���e�=�@뚺���������A�V��{�7��]䮈����W���|3��l�k2��S��R��{��mh���6����EDj½�I�Ǿ�@���p��G����Y�A�D��z�'jp6Yk@<��x���G�1' >Nȡ	�:�l���Vk�	%���$1pJXͪ� o���Ʊ�5�*�5�R#�<I��>r�!�9}oK�E0mo�9I� "|]a�U�YE������Ga�u�ׄU��2T�m�~g�y��w&!bV�y�]o����RB�`;�{3�s�\go����hB����1���j��&���,��聟L5Q�J�"��K|��
U�pAˣ��֎����2ON�8�5�
O�>n�/p2�3k��2�ܸ~ڳ.w��[��+��@���G�xwTF�2�����Bň�n�<��ﾈ�f4��p�%	�`�b�,�6�j�A�G������`?ʡ:��{��)�4��2+�I�O�Ӕ��Eζ���s���J����/Xq�!�@�l�>a1-ό�&�::�߇yJ*]y7�� 	^b,Nߋ��!Em������OK����(�R����{~�F�aU��ƨ	��,���b#���J�]m)��>�6����C�
&�4�Ȭ������B&��}��施�*��+۰��I�晨�j�͙V"  IF]ϳ������;&$Pg�*1�1�xO\fi�>~����-��}���-ˁ���F��X��ܽO�ѳ���rr��a�'fO�_��70��?���/KvV-Pz�������r6���#ʱ�]�(F��~����N�
׎Pǔ >�������Ұ�P���g�{�6f:�b��%S�k���J3����|k�SlF~3�N+�F6�P��9�7�5�� ��>cJ��O�o�XӸ�[k����P��}�f��!ى�*��y��
�M�({�ڧ{���^u�ڃ�O{�Df��Z���qҦ�XZY��y�t'���G�p���*Q�B����#��I�2��i�.����ݰ���7YC�b�P�p���\�ўJ�A��S�g^��x.��Կ��""��zyZ�*.!ۈ'C ��*�E9�bNӟ�t����o$5�N�t6�|�H	����T�����<\��.3�%q[wz�>��h��d������#�Ϣ5��˃$�i��B:v��^d?��H8�V�.:��'�Pԡ.�4��{�������v��U����om����慓�-�,�I-�����|���'r��8=n�Ym�%w��	o�$��u��+-��6�|���ų�h�#���_l�ޝ�'�Ba��i��}�D����UJ����ͨ U����,؂'�� ��93h[��*b�#��l�<<A�\�k�����1�̔���Q��ߏ/�~��3:�B/nt����1*�Xg+@xw�	߇�s'��iP3�lS��5�#:M��N�������Ąa~8�������BD���*���0���]�������YRpx\����	ǝ�ț�ؐ�e2�w��0���XO���*-��}�n��]'�1��Jb)��b|m{� �����Y��Js/1�&�N����f��Q�Ǘ�o˺��g�C��g����ʩD�5zD%� �KmN�{�͹�6J�Ɵ�?��Ӊv��.P�!ME^�.!^H���m09T�P��,;�@�-[H��Fj�5���V��-�S�cO܎�P���j���.ץ"�t���SG�e<��^��"��]��]*�)7��B<�o]��s^�u:��BLh�ñ�+f
6��_�{X\����y0a�KW��Z����N%���ЧO{���n�m�@�����yj�ZX�����ꙗ�+nD
%$���/�^۸yj9�3m���"Ed9�N��v�m����f��C(�;h�W�|�����4�R=����W��-I�\�<n��&�<�Lj��3J�CH����ŪF۞�;�d~���ʪ[��T3d�w]�@XY �6�m'��5�ԆƓ�P�FWjQ�?	�L�M��L��sQ��Pe�g:Cځ�x}SM�hd���q���+��~�M8��2��af�V%ɟ��+R�:i�p�"�3n2;`F_�g���Zp�Ę# �-(���9Z�<)��`5�s��jL:��e�/,��Q1Ϭ;���ؿ# 
�F��N�G�L�5�d]�k��GL��}�@�qA����Z!����E���!G�|TQD5�����x%�w����)�@�{��K��4WU{D
Z�yDƝZ�ŕV���s��I[��]C��.�������2�U00�����Z٦��S�m%��s$B��`'p�,oU\�4�3m�rkW�]�淲g��e������Mh��v��y�����Yl{�o[.�\g��s[imu��q�)�9'	m��|�����)5J�VAk=I�԰��IEu��6(�i����3$lm��\���x+��;�ޝ��|�#��t0�BgN��F�X��m�A�I���o�l�+�(����i㆗<��!d��v�*=��W�B�w�Ϲ�l����</����Q�ü��(g�i�p$(\��;p�EP΅!�%#������졠���t>�r�W{���&u���.f�>��E�	����?ޥ�� *���kQF�_�(%�
V;w������1"�7��l�g�[6.��,ő�����@��Hd��#dO!W6��:;,��['�����Ӏ����	�$�_>�%v��`���.Go�ϋ;������
�IC���Է{H������Cx���o<_p%������v+����gA׫�MU�k@����'D�Ҡ�Oi�ԝ�_�4=y �t�Ag���*��H;8M����+.ׂ�@���ĺ�2�I��N��8�:��v�N�M/�Ƣ%�+�6���R����ֿ��ؒ�����l�*��g/�S��e�!�^;*��׀��z"'&�X�`��z[h���5�l���J�����2В.d�u���MW�xEy�f�rkz��H!A|0�x�CE�Xi�A�r���N�0��I$�_�W��#����m���"�j��:[��ߍkk�d�ze���XS��G�Gf����xQMm~�j3�5n>��@P�G0z/��PvI8�s�������}H�Q�Syّ����$��Ew�յ�w6a��D|��wG&(�jda�4���$/jV�k����kWm�$�
km��W�[�-��f�z}�N.-w�//�"�m�x 1#@�[]������	���""�(h�-�ۻt�)�R=wqC��ӻ�� /���֔$�<o���˰%�U�׈)�p��9�*�.�YTC����m\�A�1dF"SE���5���ݝ��9I�E���Y��3�:�����!���m�)��但��3i�1M:��ª���$Ң<#v�T\s%��W��LS�Ł�2{>w@�g������#-���w�/$���[T�u7��]����.׾�X��vz�tY�-qA�\G���8���.��E2�4�,��A���A
Q�5�ף+���� �D��̓u����Ȥ:�����Q�PO/�V������~�����#;�K��-<"&�7K�b�@����Kr.��q�JE?��E��mi8E5�-�}-O`<�'O�#��r����8[91��mG[���m�I�>M5� �n��v�+����f��xJ��*�6Ķ`��������Gۨ��!�� ���Y$�����]��2w[eR����V#�����c���t�� �>3:{��Yڪ}c��-�1#�3������@ɲ.��t]�)%hb�[�~�#12�V�ň���7��@��U�T��k�i{�l����g��~�n�5�e���s�;��}�ym�@��R����ŭ�~��E�.��8A�2ԡ�W�u�5(�sxhT�3����
|���ZĊ�i�6U@�ه1m�t>���_�܌=+�3Q�O����syaޚ�O6AR��\"cߺ;�{�z�ᔶu?���dw_��O >�XB',ʃb��/�5�i�߷����<���x�J��i.1A�nJ��9ē��*8�"?I��0RL$)M)���J��&�x����+ׂ��w$�t�א�U�ie%��c\�G�7_*����$�Z����hV�����'�!閕ٙ�4�I.���Li�F��ho�紱@�a�����4=	n� �w@�=�vHx�#�)|�؎�d
��|#�X�5@(
�f���
����W�`��{�ɷK�����*��ĥ=�T�?|Z�����������n�bϻ����	�����wb�=2֗�n�']�R�!�BN�x]����0Ab<�:�ɂ��e���}���� �������&f�[YL�K�ҳHdip qdf�"���0���@�4�� K�Կ{5)�)C�3�Q�wI�^Q�T�T_^M�@c1^����]��ֻg����=��^O��v���.F�.g����׌�+h����:�e�b�a�WZT��"����G���t~����f�ӧCLp!��J���d&u�oC!K��r�t,Z���5efD�\��c�#���cT?-��y"��ݰ}�k���N�SC~<I��:{�'��a������7y$%h��N'���C���l��g�摂���\XO��xJĥ֐�Ʉҷ�K�,|��ɾ�݌
����Ǆ)��r��O��e��j�T3�}7�	 WF]ǻ��`�-����P'8҃��mՐ��%�Kaxփ
���br}��Z�F�g�*�Վ(S�<�&�n9� m�"��/: �Vp^a>��حl�s��Z�
K2ffk.1��>�r�������#��sy]�� ��0�3�U=�k�F��s)	d���w)�@��4 	2O^O��Q���K��L^JUc~�d����#ϵeE&	��K�^�9�_�����&��l9|*�Pk��J�H�3�_t��T��L8�d�r��pY0�}�V��1�ޤ'��>�md�L��#̰8�)�g��YT!��Uw1<.�+���S�p̟8�ʕ�Hg!�����<Oٛ���ߒT Ύ�#u��oT���:V0m�֚d2�q}����am�%g!�i�~�����lj��.db��?o�@�(��E��sE�(`RIi:����o��o�o�PC~�H���$_0O�M���Z�mN2���(G�ڽ���Cb;��߻����p�{l)�Ad��#7�q��䂡'�`}#����j���6o�ũ������m=�jߪɰ�*X�}~V��I�X���F��=-Y�5���ai7��a�;zO�+O��c�&�F��G�n� ����R�MGʕ���$���Wձ㫈�W�Nt1r�EF�JVAM���I�����R���n�������=h�)�k_�i'�ORѶFS�P@��XWy4��	=I������~P��@����ֱ�
����c��~U�8#<Ud��p�� X�&]�$>JK=a��\+�,7Iv�&[��P'�����_�ҿEY-����n�������t�ŭ�oc)+{��Z3|Φ��#���t��ԓW��{�s����$��xf��8/��l��yV'�J\ζR�$��0\����*{��_�����ؘ���#���D�ۛ*��9_����?��5&0)� �t�@���B�|{NTe;�(��6�TR��0�1������[�z})�𣆥0WN6*;���L���rER��|��A�j�0҅&̜�ِ�UGSy��e)��j���:���=��1���AayT�j��osʩE��]v�g;��(&�qH�����5��a2���/Ɓ�)��?��%���0'ۈؓ(J^���&�c�OB�!�mBSh�U8�	�	�2�}�Z�B{��~~Ps�Kd��a/<���@9���j������׹rg����.?�T�W�����1 ������r����Z�}Q�02�@ߦ�X%jD�aU��f6{vC�Y"���ҩ�>2��
!K��L ����++\z)�Ǌa
:�g��'m_�N<�d��4��
����l�9�H��T|�Qٷ�
n}��$e��"�J���w�)~��K�=d%4_5�D����N���t9X�F
U���Hd˅�Q�~\�"���V+<uY֘+�?<E>�Q7hn����/���Ջ�f߀�{#��;�`G��� ��B3���?M�̥/�Sɔo�����q�hMr�6�l�|�!@�=�	�a2V`5((��7�_��1S���@[/��dS�ǌlū�h=��A��]�R٨�]v'���׽��G�[�xR�7��Ƣ�ׁ��m=B��#�Jۜ�� /1��:���L�f�t m��b���]һ�2��X�5�q��8Hn���M�#��)�|0/P��^`q�5af:���d�$�d�#�|�$/�¤bd��ʮ�OV@4�/�tq���xaĄ^%���%)�����s}�B/mc��#Z7����؞���U�/��t170q��O���2��pz��*�%�/�,��2��٭
�9y���[?� �P�4ߖ�x3�Y� �ЀJ���	}&/�T�r�J(Ӝ
e��P-�%o�q��uah��j�/����2��7[�6���m8�מ���]	DxOq(8-ΧQ��+��6�Hֲp�/%m�Mi����ڠ&�N�+�'_��?��~l �m�u�{�]�̌�R��%0��d�L�ޟ�OAw,��'a 2݆ �Y�b���x��	�;�@��4-~@>��g�^��r���]��A4�/'��e_�r��$h)��zR�Eg
@C��h�{���*
�����()h,P`4S�����2�@�b�ї�a��)��e��F|�V�w��6�6.�d����k����[��n����`㿬��op<=+#B��3j�-�᳷��Rn�y9I����'j���Pm��q<(�R�Q�+�,�یX�fV����i�떐�g ۈ6�U��v���� B�p�9�LbP�H+��[qn�� c���;��y��mM��?��Ġ�}U@���0h��g�L��I'C�`_������ě*oI%����׳T�������?�v�ޭˊG��/) ��0��Y�;xjܫՎ4 1i�Ƅ� КX�M���F����9( U9�*�D"I}"�R����;0C�F�:\j�d�� �
�5_h��>��@�g���;V�YV�g���jE�!��!z��Vw�K�j&�8���@�/�u���#mp��5DS�
KTa��&��4�ִ�Z2ĕr	�"K��W�
�VAo}i�HO	y3� �(~㻑����zᳬg�:8N���{ޞ͎�T�6;�z{�\����t���*�������O�S�b�#�Y��4�x̪U�M��]�"��֍�dM��$(z*�N�������,��h�~o[�:*s�JJ��:k���r�Z�Cpn{ׄ�W��eoi,l�'夃.���:������"y
#�l��P_@������2jD��(����z��mJ���\��'E9��ڃ�u��Q��@���s�2�/l�Y��?��+?��<r�����'���렗X��p!D�Y����t�S~�=�V��Oi�X/�!\(U�cŉ
�ܝ�,�ߩQ��T�>5O���3Ǜ���@5Ou���?��l�t��B�N7/1������Q�!�hJ��!:1X��:�o�;��iF�<n�Q2�7߿���q�%"&]�G��W��m�@~�Slh�|\�Ԙ���l�(��A�{b�A)��E��h���|��{: Q�J��W�@B�o{�^NJ7[�Z�)H�'U�Zz+��A\KqE��$]�vZC��f$����bR'=+&� �2�&ם�}�S�jU�7NT�$Ы�����y�<Ć���x��ZDl��qktnʪ" ���S��?�݃�/�0hΑ�_�D��HK��1����;��4_�WBRj=��s� ����**�9Eq�5t���
�F��s���jA2������D�gn�:�(����+f����5����S	@��>r;#Nw��eq��Qq�7�s
V�&u������G&Mj�Z���K0����g�K ���%�O%tQmD����$���KH4�;���
05���4�W#�(�%��!���"�|�h�/�f�˺ӊ����>]0/��^Xx���V΀:�eL�$�I�(��0��0���N���Ir9)��6�2�exx���j��\�@�',�p�,k���t���;�0u��"n��v�V1Ŗ���$�*K=��-��q�$2�����}��)�x�K]o��\�{*�"Pd�"�ݵ�cRp&VJ��1
N��dϠՐ}[=l�w��W�5���*�X���r5�����*��?W�0A��EL�����D�����Oz�X�u��8#�5kta�mS�*7�y�i�D�B�QD� �ҽpN�A�N���45���A�̱,UZ�J��[�ͤ7F��ꖁ��޶2n�������,]e�p�)�a��{ɟ�o�� �\I1��:'�m�,��"�Z����d�]���fAʅ0�hV����uE��A�@uO�fPCT� ʉ���Q�z�����L�*��j�e��A������i�B{Z<�<�`����q3f6�����44�Q���#�+|�	bnKQ�z_��~��U�s[��S���*�E����>�������3�!�oڎo$�+�\�K��@�����D0^����uחI�%�u&ne�r_V޾E�����e�K�{�MI׆���r���u(�3�W��.�&#���	L���C� �G�r��0��7e�B-��t�z���\���@2��C +�'�9'�r��Ѣs��2o��kE�Ю����M�^�s�!.46I��>��K���ͬ��Ý4��v髬�7O�F6�I���MA!�����ސ'%����X�y�~:d��)��}
����.Dz$���a�9S��ݒT�@��?$I��?K��V1�[�N)`���$��uJSl2������hc���K�h�*�{nܗ��h��ޟ�7�`�K��
M�>g�Q.��}��B6T��Цu�}�����bʘ���2��OufJ*�Zs����g����Ek�'4ړ�� ;t]z�d`y0����}$h�v���5���{�z	���!�i��d��<8Ӈ���ύ����J�76Ni>�RBa�F?�Ql�q�N"�
��D�6�UH+)1�r�k\���g�]h���^KFlIE��l�Ԣ���)L^��G�5�u��I�-��%��>̞"��|Br�ڻC��F�W=O�?8��S��&�����Na.����_T���]�f�K��,_��G���8��� L�U��j�O��Ϻ�g]|�X�,�f��|��z��7�xD4���9�W���{Q�<G�*�>��7��X�ϽK/����Lϖ�4HF�	�� / �l�@�1�@
��6�m�����yg��'��O���=GUC\�Y��Q����E3�s~��� ���^� �����c�yY�s�;潓�X�@�}՘�q���/a5���[�=7���3?t�sDm#���j�����5s�@DRg\$o-����5�n��ܦ�z�8X�
;s�K`���V����5M��ҹN�)�A�Ż��}���VV�	<Is�c��ٺ�� 
���*1Y;��l�j���p���"�6���ε�D�Sc��yf���9�
sǌ����6��Z�/�~jo�O
�-�?��g���f�� �W��0�AS<���1���rrK�����KP��q'�3����=���s��P!'���8;~l�}�Ą�s��tdG�_g��m��ݜM�ĄE^��t��v��GX*��#�8P���n0��D Q7.&nO;w�(^�'s�œ�G�N� 	���ui�,�hN�������߾��EF�m V��x�v�RU�#�*E��aK� ľ�^y����̇S_y�J�Ox�7�g�@44<�N9S��@�n0�n�C�㑺�Mp 5�8�� �L5*N��'i��g�L<h��n�s�^bp6')�筌��A]��U&m��x�[��R�O�`�����2�޲4���lK�mU���bfK�sy)�B��D�Db��z��WS�CֽՋ�bw��`��E	�NO)�5L��9`��鋐T㌅�7Z|��.~9d'�f�̱�T�P����@��G������rS<+n;)���ߌ�I�����0ݿ�SKpP�fb�"���6�Hk���s�@�@���KdD�mv�"���Vf��QZ�I���tRp4b��)���e|�L�3���2�q����'��u{2V�1'�T���a�߆+S#�#[L��v�
�ɵL�~���F�iY;�4�W:��~R۶��o8?Nt��b��5u�KZE*�_�EC��2)Sؕ���`>ޗڭQ�(�Xg�Fo?������sC׮1{�/T>ה������xF̌u�:v��*�����l��XtF�]T��Y��D���qp(���������׋g�:��]v���e`RFEN�x-O�?2,0�V�a��K,�����*"�0"�k���%(c�����Y�}�O݂��P=*; rD'��H��)g�6�Yt�+ٌNiL�m�?���m��rmDf�$
��CҌdM��o���ě�i���j�α+f�w6i [6<�<P�4���P�h�p5�P@˅�.$V���H-oՎ�\7dkOu��d��S�_L���(��WH��5��r;���-�`ҝ����MC�IaI�#�{�w��I�b��=k�rz�i��<�i�� �!�®)r����*7w�^��2>_}�^j�*}��G��  ��+@Yg$5�yB�����������c|䪪�|Q�MUQ���d����א'�C��ihz��3�Q"x���W!b��XF!�P��S���-$ҳ&�sR/_�Η?�L{�$L
�J�:���&rP���$*�L�VV��_$V�`K�p�6���0�zI��/*��%`��x ��_C���Vd��P�o�6���o�ս�g
Vxj��~X�������	t437�yj3^�i�F�����/�^f���U����V���P;�_�uP�Ŭ:�F�����r�՜Q�����-��kUhhsd�`�Q��%#���-�3�����s`��0��[Z	��8m�$P:�(����+α��k�������=�:ԿT�e�Zd���bO��(���N>��v՞�!��)�Sǌ��bj5�8�w�¿�0M���0�u�����`ܰބ��h�v�=Ғ~��I�>�?�G��<��L@� �7�d0QS�|��}sro8Y�!�W��Xs�����Q��N�:nٴj�Oo��_���Һ���,z��#'"o#"��^�CWLӵ��Y��Y� ݦ�?������3�M�Ɣ��M�g��
1Z)�H��C�m)~4�Oݰ#���StBD���׉1__�B��/�_�������_���NEiH��G�w[�����.Ku�`w��.��>_Q�@#o�M��v8�6B�k?Тx^\K�<��aF	ŒMk���DX����� 0(���h���Ug��=B���]+�:a���A�)P_�0�C�M`@��� w�Ԝ��N$,B���+��š�6ϝ���!⯴&��C��hPF�	�,�r7��5�۷���R,��f�t����HB��f�'��R\$ ���O�IJ��z��@^��4d"5.�?����u�?�P+�������ﱤ} �(��O8�m�r�R/]^��W�#@<�Ju��І3:��;���#���L��z�|��r-2�;�v���ПY�e��)�-�7J��(��a���ɋ�y�7�;��;~��o_�e�i|��ϊ��О����O�(;6���Z��6���-��h1~��n�Kh_j"�������k�a��d(R�0D��C�BV�\�!���H������6�S����Ka<��f��R��$É��XO*��mVQ�f��n��#��n��m�N�M��1�M���'�a�0�.�Kn�k�^_k� �#4U�:���M|Uek@�YLc�O��qD���3^<OQ�����#j:N���r���v�0���n�\xV��E�Vk�D�ޑC�5�;� 
IYk��ů�$�1^�#��D�j����0n(:���1�������`*l=�+�\�4��U���1�6�|���W�e���3����)�<+�9��Iʕ����I�DCXÊ$������5�e#��ڃ$���;��^�n,�MY�+�3�l%��ey;Õ�&��<���þk80r4`MtIMw��ݚ�h��u�����*��*����sG׬b$����T�q ��* ",IvLLA��� ���ǽ
g,n��χ!�!�Ӝ �!Ϭ��P��r6�rC��y�i���'�����&�������U�F��v��9��g�v9[DB�����J"]����lY�<���^�p�ͦ�	͘@��m`���9������������<��ݱvË���\[��(��ø�Z�Y�ߏӒ���� �z�Q�N�����@�7��;m��r��䖏�3��㲘��dI�����u�=�Ҥ��ȩT�W8��;<U4o��Q0>>�]O�����鰒7&�|���t�_$�os{���l�8Q� � ��]�eO� r*�d�5̄��z���x�Y�+<����"-��5,?�J�b#f�ud�G?Q���~����$.���4�����A�������x1lҳ*�l;3��'8䇌�6��N�+	W몏Ve���2��rֶ�D-Sc����qlP�Ԗ�d�%�B��Y�Iq�(~C�J��A;Ɩ�����k/�/�ʯ��I�I�ǶmO���:��y!bQ��2ށ�\�҈�%F�ĩ��f�*�E�!Uo���8� �J��0L��1jC�
��>넺������糛h������s���.4wN����O5W~{5��y1���fl��a����p����L�;= �O�0��-�5���b�>.�.ʛ�V�a÷U��2����E]Ҧ����8�-�L8��`��(${ʀ�Q�d�]�"J֯�oW%����)G���?�����e�[C�����Y�u@�������O�(��Ϣ����rDL�>�U��`����D�B�
bE]^�F-�ڏ�
��P�Q�n��V�!YT�	򋦠�k#Rb|��@���9�j��Ǐ�c~nR]nKܡDU���V�qM+XE��O/�'�@`��L���Z�(�j�t��C3	�ߖ�$�"�1[~������d�S?������3w��ܕn���=G@_|v̡^	�{�'1�y��k��I���5�����6�
`IMT���T}J�-�V���ST�x��z#��~���;�yōlq�s�Wo�R!�E����>t��~������#�Bqb��nte�#��-�#�$��N���ݡ{M~6�]a�RJp��f��� �+���W���4!���<�G�G�g{�ʠ��\@��lu��-U���U�0_��k��$6M�rcC�w����6��xMi�{q_�.#���
x�%W۳�u��h�J	;2K�xlT>J�7�W���a��Ϭϳ0;�F`�LXҿҗ�$�2�:ŵ6v{�Ec��7��
�����5����L@��f�k��-�s{��C�Tl���sx���ɡ�Lh�,?��n��m�ݿM�h���2���"$D��O�,�w�7����ʬ�7�K�ܡ�R��i�nM&�=�⫆i�\�#G���(y��� =�;Dzb,��p�'�u��Vx�s����W�Jyk���?�K	@���4@��o�o������)lHkd���ד9�-�z���f4]6+�#�x��od��)�q;��-�m�,��]�1����:��#��$�0�1����R79B­G�;l<"SpF�>�@���U�&���f~*t)��'=Ez^���<�A)�3jb7x��3~�{�X|�<�@����(�rJ�0�W0����UfhYr煈�]\�7����hx�����׶����K<���9���ђt�\^��iT褆�f�_�C0�I$1�/%`���_��:a������������E}?(0�_D "m��{TH�F?�ɉ�����ɜ�����<�� =Ŧ=1�Z�ޯ�_(?��t4S��C�>CM�]�vn��è@���\�U!���bT�ԓO�y����S��=�q>���P���� �ue�w�4�Y�h�������1q�������A���Y:G��Bm���d�;��[MhD�:C��Iu�2(�.��ĵpe^����lI�ǀ���X�X"s;?�x�˺C/2������g̱�i�<���L�mB��8�����$�ֲ�6do�
d��fIsR'�8�%��b���n�+�]!��1mH���.6M� $�U�Y���%�d�~[Y&m^c~��w��[Fip
���o��QT� l]�fs�
T���g�Ů���!ד+�>�:�>�l�9h��)ߣ�[^\&PxA��QR��f>�� ��,uj{����O�N�ڏ�I��28�(T�����Z������%��Z��41{I��mU�c�$��za2��p��t� ��w�4wi��������T���~벲
�/�xu1��[S�3A�!�_+�^����
-S�t���2&��0g&�� ��q��J�OO(�r�e�R�-���Y�R���I�) P\X�!��K�O��b�h�}�2�S�Ai$]֡5D�{])N���oJ?T�`�n2$kY�ژ����Z�.�r����vi�`~��x 5cI���	< &�3h<<����6��},�ض��I1�ٽp]Ɂ��pv1�p�n;��kK`}���P�:��� �S�J3�8����!��}�湋3Z*�Ԣ�$j�C9#����b��>'���Ո2Of�h�ʃ�[���[R�����-�һq%�G���J�Ai��d�������l`��O��*��6��G�
|���w�{$�ca?���~<ug��m����;����'q�O��!��NǓ��t^��-�Z��N����j-՘��� }��i@O
'���m!Y�r�=�[{<-f2���ߕ��L���//B����&O��"��E]��Ы����e؁�2��-�G���x�j���h�P2�GY�C�x=\q�Z����Kx�U��[s�M��|�~�����F1gRKpbkIku"��&��<dId3��Q]�R�s/[J����HY���
�a��^77f�~ TX��&P1�4F8֊FT��g�S���t�(ː=J�IR�Y-��^ؐ=����Ɇz!b�7�p�{,�%�v+թ2�h��H=Bc�)pBU7���Ʈ|{o���`K4�m�Cܗb_B�T��%��#������V>� ��]�w��d�� �i���g��΅��v��]�=����0?����4������W�OV�<�=.��l	���xx���q^(� �����/*�q� �?�n�WS��\��*i�Uϒ�͂�%�E{�7��F| ]�#�m,b���B�6ܶ�[��X��ά�=���d@_WP������|����k|�M̏8�3K���֢��fۻ�S�����x���>�E�r80͍O�����`OE�E�T������r$m��4�hx�v488?h���]��<�`T�wU� ���d�g��S��b���k��**�����y��n����!Y���FY�6u�˿\! Q���q�?�@��;i���zf�0 X�z���b��ǃ=��M�N�}�]���*��$=���s���w.B`�0h����jU��h1��,˻�^MIm2wb|[�	��c˕#�
���$�~�CGa�ca(�mU���#�>j:Z�Υyg^=�+Oi��]3�5�����"�i$�
�������4�_�:;B=��V��!�_��}���w�g���*a�M��hX��4,���ET΢@�DΥ�x��!e��=�d��p�rQBh��>{��S�y��{V@__��oA�YK;6ٹ��2D� 6�E[������l��ܴsd����������Oڋ� jce�yU�gp���l�=�C��r: ��%4�G{_}�M��7Y\P��5	D߬����~�
l-"!l���Q����ٶ`�P�#�/�_���A%�Rp�]���d��>����޷���<�`���}��R��x�����"��gr����o�P?��Ԗ��*�r?���<��Po��973��f���ى����/�g���e���,����l�Z%sW����q��2��P��ϕ���hb_ڳ���
�.Mc�+�}O���g������~$$b�
�1���l/<�T��R�B��87=q���3-��CJȾ����
T�Xp#�w_���+�����[Z��s�Y��1u��FYv�pl�/J�b)��_~����AD����?�Ul��4"M�J�_�UdA{��5nu@U%��*�ֵgfP&��w	���\L
�Kɏ�rn¶���^��i�,@��tH��9^b�����mF`�x��k�C{�j~�]�LwY�sg�u�(j�6v"�hKw;�r�\���|1�LƭĢ:4��x	)n�eftXڱ����s2v���[F&�TE�-���j�;�jҌ�/�j^�}��;�����W�;R[eG������?�IP�M1��X��TS+t�r��|� C��<�1賋SD���A�;�Ƃ�2�Y���[`\JP}���)2��@�9��!��$q=��g�����",��q�S�z>,W��G����N������[Aũ�t���&G��9W{(�ڜ�;��.�)�B�I	��Uj�\A@f��/��_o3}k��3� ��~z�)Й<�n�]`�淋5=)���:u��B+�,�ˏj�|_v��d���2�J���pcgƈ��-z��X�(%�=0�VB���mγ�& �qB`����֎զ��ob�,�Si_�%\1d�ځ�5�5խH���� TA�F�l:�������59��F����HG��:��ݜ/t·@���w�O$����J=:��@��e��]E5eVKG�M�o�`����c�ɞ�y��r���h�3LEh�H�8�aݓ�;ǩ�V|7�~����9�|+��6@I�ͧgI�8)���2�=��a�܄�"�X��{L?ro|G�����D!M�� l�F��r�Zd��7M�&�_���W�c0�pǑ�"��S�zR/�����Վ�f@��>����6f�Jq�)�]�)���n����04fX��.�ܕ�j=:���B<�u����m������P�s�Ȋa��E�1���Z�D���?�����M�c���N���!�Zs%�eٍ��,8v�\�/���}\ư^�z�a��g����Ah��Bl00ZoX�O�>����?huq{(����ӟSĨt��>����t̤�o����ogk��w�u�#��戀�R�T�����68SĳwJ�m��l� Ml��smcχ�0�������i~ӟa|���DϺ0W��%cb�6J�5f5���-,��95�Jd�"���+0^}�F����]��݀P�"/��$d�n��L)o�NI��_�r���j�ת���V:*��%j��1y-�*�)�A����|�g^|(��s\��]$u��ms:[՘���fx�Y���"FsX��.�PU�(��,��Q�k�{��i��_yG U��J�� W���1jM,�X��`x�W.���P�iO�v�8��}l�$�d, x*H�6G�f��rT��Fg
�������X>��HJ4ξ8�Zd�}�Β�@M��f�ŋ�A<WiA<=�io��P�b�'�%H���B�.�`Y����뽗��.��u1i3c�9iX���!�6�9�$z�d���v�=�{�Zp���Z����v�{@�r�9X�J8�Q�j�\���t}��~��A�od�3
ʦ�:���b3��<�xqف�'���O�a�oc�A�C��#�h@����^&0o*ߎS����v`ɄֱĬٯh���u���!�-��j�˒�Q�#&�򰄤h�����doiƲ�8�����������v�H�K:g�X�z��S�����������3����v"�v�b9�c�҉���u1��c����ӣ���s��r�Bj!��j�;�2�!$���;��*ugK�$�������>�ZhrZ&BUO�E*]�ƀ�;卖=�oH��ZT���x
�e��}2S����aNe�5 uR���ʟw��w��ݜ@9����k���;Aej��������徆�W0�k���"s�]\0���ȿ��[MP]��$�b>�cc��ܺ�����4�d� ��f�S�"`ZQc�0 �5���+q�Jmx�5OB4`����2�j���(v�G�k �+�l$���@FY���r3��z��Ӯ	�'�1P�z��=!bB5���{(Eup��k��ˣ���	CL����Kj~��v�V��^����s�$�Y���W��}�U,޺Fq� �ν |R'+��"/��-��Q��}��@�i�.ƻ�ޙ �f�f�!b�Og�̀8�ݭfy;:�\�P�ţFOS�ka#�n�]��c2�p<i�zz;0�H��R���[�����Y��	׀xnG�-C_ůʾ��%���fas�ll9�~�';��x�}�a����!
�l�1|��&�;՗|�E�!}��������T��ҥS���h��H�����W
�K����0>Ws�*�7�p��yk�"ԥ7�J�X٦��cq��3�e��<�M�%Q�Q4�]K	7+��1�/���P�n�
=��rn�ħ`��n���[`6��G̝H��k3�0)����4�;9�M|E�*P��j8�:���
"QM�{ӾK�Ȯ^���P�+�o�P�p���tI�ρ|�߾��ү��M���'qu��d��':��T_�� ��6?�Jݪ����& z�$<�5ˀ_F�x�0��<[Y���bj
1�P���8K��d`C����\,~����d��<F�}
�σU�/���]�*Gٓ�N>�$in%�eй��HJ���T��~��҅��jI�J9�޴F]ڹs�2_!�#%�T�%����g4�������F�x�Y�ą1�K������rE�;�3�Y�˲r�?�J��3M�AŻ
*N~plӡG�sȾS�A+����v� ��m���u�!�qL����ؾA�υ54�:d��>r�[���}��^�3%�"�3b�b*�6��c������2�]���d��c�"3�Si�-�X�~KB�w���F����N&��[����n/�9B��L<��̆��y{�J�Q�t�fY��3hH�.�H��k�����l�%�$E=~�B��ZM"Y$�9G�qP�[���z�䍫
Fw�#J+��u�9Van�MC���(�b.�z;p�1M��;����}���w�5k�K��`���]~N��P��p5�֣���<cfr�0^�������R�D�^�讼u���Y�+��`��mI_�ۙ�z~::��.Fϴ�?��~���dw�N����m�������V�b���^�xԎi��r)yh������پ�IU���P70OI��l��JT�|At�t�l���Y*d����Q�F��!K�� �Fn�;`KOѱ��A�̫Y�3)��M�鈾�RZ��i�L~�$���/l��]��)T �p�[FP�]*����4�u���L�o-�5�A�5�!~yWΐ�pw�����Fi�L{�x!�bw�R^������֦�]i(�*��u�5G��K);-w�Ce�Tu�-����~>jBxۅ�!����'�����{�⊛FL�$i�qL.Xk&�Et�����վ��T�g�e��-�5k@+��0!�Q��=�>�FeEs�v���jC��Uʽ{*=��t�l�4���l���� *�	�N�M����7�7m-`�O��vN�����{�2��6���W^$���v��ƁD��(��σ����-��E�ta@������.ev�Eѕ�/�,엓L����5�T�G@�7G��G�q�.��"��B��h���^��2f�6��m[n|
����h.���sNT��*�sTα����m������J�wZ�\���;����uD��HT9v��X/R7�g�ޛ�Ȭ:�b�*zb�kڭM+z�)�I�gG%���)��"�k�!L��'CV���ށ���Z������Ѳ�t`0�m�]����gzxk���(s�#���RG=�� ����YҜ��y�@KQ;w���mp�ӄSPyޙ�$W��x�����,/�*��솠�u���'���1[m��t�b�ѧse�*!�KD�UE�>{ى�!P3\���)�^�1/��O��'�Z: ӳ}����n������pZ��z����E���� ����"�ɾ�B�/�G�j�0yh��'B���T�op�-C33��)��E�w�����C֌#r��z��Cڟ�گJ��V�T�=�U�|S��+�=�e����s��k3yd�˨�We�$��m�oy)Z��K��2R=���g���v�Y�r�AgMq��x�BS�~�.t>��}/����z����%�V�e������'ch
O��	��jdL��5p4.���r�7D��L��E0�4�����4}���I���u,�M7����Z���l<c��0��;ϝd��8a�Qx9ߘ橵��ݣ���(WKT�]�>�<�y}�u�]��(n�|��+�;sL�)���Z��j�S��0�����q�͋����f�{���>fjM*��SdN2������*�1~h���~ʔ���.N��S�O����K�VS�'���"��1�x��!���Z��:k�)�Od$G��ڍ�e�n�"� rW',0 ���}��b+��֤�3�c�Ul��2��t���JT�	�(N���!������x������鄃�����l�/���an�Zz��eDx*�Eo"M�ZLxT��O��&WO7e_L1�4.��ΰ3Ўys���z�9� Xͅ��Y�@���u"�}���vx֨�(bP�	%��^�j0�������q?�*�ݺ[!�z#�n��_�،�tU���5�W�P�b.�"^je/&cπ\��� �ߞs<��-�p��9)���#��x�\�!��5Q��0|�Hj�
��@&��p��/��m|�ϲ��`���6H�ح�d�&�ĉp�E�'W玻��<S	��	b��%8՟�����uL@7�����w�T�A"j �z,=t"Y���Hs1YϾKڙx�&Oo��|��˲2����KqJ4&�UluF�-Q�M���k���皪����ㅳ�Ҩ�V!J��'R�U��uӵ�a�ݐ�i5��bYݘ&������x>���@}
�����������j���z�Y�1��x
)�܎�[���Q��e��R]�ج��Q��kz�~�YC�^�5�O�tPi���p�ʃ���c�QFFl���1��X���1�u
�*��:����:���/\v	_�}�Mћˤ�i��E%�H�NO�m_���tx�*��`�����
�5��	���؁�'��Ǵ�٠�0��c��5���7�xp!k�ݠvW�F ��P�0���4�
,�L=Q���`l��߄�r��O�f�#�,�òVO��&�!l<h�ނB���k���q!���L	u=�&�DG��݌F���c�7-͐> ��1�ct|b��]4��a���:��,�r@F�:�^�X4�ӊ���̪�K"~&7���u�,�>N�J�b�~s
������ cQ=�?�K�x��Y·�� ��-�Z!��-5L�` �G��w=^��;����=H�Re�Vj�w+��BN���F�cR�0a��KN��m:��4	�ً� v�%v>��e�m=�%c�6��ގ�4F�}��rRo�.3��.���G���0-gu򩻑]����|���ae���\�F]!���>7��d��%ek�RH��AI<��N/+�4��W+Fz8�Z�R��C���t���h�(�e�=aA�y9�x����zǽ�M��V���	��6;Q��FP�H��ٍ���M��6R�D��9��ͨ�eb�'�(#��%�P�fX�ès��鿙��Xp�AW��٥	�Ql!ef��-2����)S��A=P���7㛈-	Nfg�9X����6�$N����w\��� �j`�댇q(�j�F0����d@�n-ʯ���s1���f� �?�5V�	���6����L�]�`P�s�<�%V*8k��Os�c򳣲>M$�Y�?o��I�+W��X9�D�:�3�'}ɇ�k���ҞG��xV7+�;9B�9�GUF>����"LG�OSd�z�~0>%,������j��R*��ow��Y�MA�n���_��ϊdͷu)�/����(5�-"���ařu�雝�n�a��h���0P�_����`�Z]B�5��oe
��@���VjZ�j����2�U���j��>��K�<��$6�'�*����,�s�
��b���jo�N��hJ1��U���v2�E�d.�����A&�<�w1�>�Z�V5J6��|<h@������ȴ5R����(M�n`�% �$@��Т���f�@���9�@�V
���e!ʬ�߫�휆�9w杭��G{�HjU�,(��,m@�U�XA��!n(�_/�y0 �7�@�)l�����^�U��a��9G`?R��uOT`ǹ?�P���.=��MC�IX���~�.H"�24�@rA��@fޟ�2�>d�{����I���5�:�ުi��b.fzņ\'6M���J}�a]�ep��i���+�9B�����؏�hst�"�2BI0�(=�3�r�nu^�*��5r��ݮ�5U]Xf�i=�����e��A�戶������+YM��/�]�v����N��5�_T�dQn75�33���J����nc�f䄹�}4���9Ӭ�kr.x�Ǫ���� �D��T��^�Ҫ���(�_�JmY~%0��z���z "�㏨a����149J�UK4}��+?�pubA o���Qhq	�o�&�II����d4%n4�K�B�ǒ}����5 i4z����BS �Q_�T�>�1�NS����;�Z�ַ�q������t~Qi1d��h�j/� cёc�cٯ�D(��	�[�R���Jr�_�&�⹿�
}2y9�#y0V?�Edb��F�Is�g�V#��{I��e7Ў�8r`d�
��5r/��[?O�I呏�4;V�PG���r|BP���!)�|�|�=��zЏ��#���"A|�Z_�Ȳ��p���:�jK�2�6.Ҋ�s=�x�"`�����( �d�DH�]'{�q 5�/
[%�ڏ"��������kҮ�1C�g)w��V���
0�T� �Cl	Cu�+���^����R�ۏ�vD��Y�-+i���@�CI���sрzÜ�ǖK������߯�VA����{ѫ�+.)N�U(���H�g�����If��'�F��u�������F��GL�F����_��R�4�*��>v��X� ���s�H�T {�OŬ{������y��˛�:�pWݘ�c��A|UHB����ga���a3�Wq�tHI�,��Vp�6���g9r�4�E٤-�������` HC��Ҁ𲡽;���߹g��ި_U!� x,Z�Ƈ�^:���}L��{@�c�.�Bv���)dw����VC{t5klYX��P�tg�10��Cz�����B �����ߗ1	yUn?V�/+?���j�m�����Ǽ���OM˙�f�fcߌ\�.�ܭ1�*�J��W[a�Q��w7>��z�K�7�%������e��K��|����-�-kS4&m�4��D��Kp�0�.Tfna$����U�[WW�$�� �e��� �4W���8*�y*u�C��>@ޣ�7�|R߽Ga��G����}����m��ħ�`�)S�LL�<�Iڔ�+ �WEh2�������Ȭh1$�y�S|�M��H��?f��{��,�º0���J�,E��&������.� C���
|�Q��r���������=��	n�ki�yc:����u�ܫ����p?7�:��\���;!�#�<��:�	��/���
�`z� ���o��1��uC��j���;E�s)�SWs,�@��X���$�n	���ÿ��(3� +���x:�ϯ�E}�}���sV冭��(E��Ұr@���G�^>�X���'�_���iBy�
<�v����0�(� ��
��h�f� 3�}i�1)1�a���85'Ƌq�WC�{��V��J�M[��Dp�jah��rY{T����ԧ����4 w��j��M��;©�{�)�;� ;}޳K�[A6�DK��#�%���^�%��ׄ�sM�]�U�Qߒ���EՀsظA>:�1.�G'�.��`� �)<���C��#a( ��}�u�Ay�g�+�9mᗣ�`�US��P+kr�� K	���� T{� ���G�YP��Â�f�v�1<wue��9b�-��o5�p�Zo�榰��d*�A��M�q}0��N��D��U7^�,�	�4����Ë4�D�f�cK�@�^Ak�-���@���W{�V�(��������o�D�s��,�-@�����c�����3�K�y�I7�\�	j��t/�/���C�}�J�%�7��u~�2�r���A> q����;�J�U2�f�y��٨�~c�=x��}�G�K�	՜�4B��l܌?Xhɶ�wX1��k�}Sy��!�#�xܥ����gۃ\?Pk��$���4@,�w����K_�QS+�{�l7 m=p+Dn&/�w�5|�U���Ʊ�V@[����O�J:���w�)�+�t�0��#u��⽀�����L��s�I**��+�C�f�PBT�s���[T���V ����d�!�����]Ƒ���{7�����D�s�B	�F��Ѭ��qS�0�E��]�ދ���5Mr��	߫�ǁ��kpW�sQWCt
)���!lI��,��1� ��4<���r!�H��#S�L�r����(�2��0�gdH���S����}��M���%�_���5H����@ ������ܵ����L�>�I��c��6�!�S��SbVtS �*BG��{�bփ���.�X�v�aP+�*�$u���F����f�0@q<hw/�:"3ʇ�|B��7��Й?�<2Y���q{��p��Fȫ#qW4'����]�X1��-x��(�,g��Oˮ=c��G������z]7���M��\��C��������9��Ђ�rR7�� MV v���hRx����q|&p��̹�������E��"W3�c�N���]�nꕗ�����W'[a��k�7mw��=�;�6�cӟ��m��� �Wc��犪YyT����{�*���NeUM(>�f��dWх,K^%g��:C2sc@�o2ޤ��u�X���n�.�E�tK[�wL�>í�:�p~��	��\z��yc�1�HI�������=g[��C���guU����H9;�M��b1Q�0��#�iVr�Z�;А~�?����3����",|�t�w���6���x�y���� W�`��_���3�M`��3���)yq�	q{����T�?�c�vp�D<��/��f/`�g]�m�7q�s��Y�B��8<GO�x#oq1�X�Ms�$E�C)޵Ь��ĭ-�Ea~`�@�w�Xf8�I>�sbߍ)\�z���lc�H���e2�i����G�C������H�ؔ��.����L1�O�Lqw�^�ݛ�%g�b�n�:{v%f�bJK~נ_�痠��u�����_��z$�;�}�v��[L�Q(��	�-&���r���q����5���
�F	�9PA<��3l��:�Otì��1��e�NY�]�4���}g�t�Z�U �to������8�]��C�����pJ��3"�Y6Y%�s�w�)~�ç0��s ��^�r$�Hy4{~��뜵�����sBP̲��q��g?�(�.�D�S~
m|.��go&���O{�	'�o�G��)W<���_]�k���mnw�������RQ<�����0��A��y�l�K��#�oǧ��hs^{q?v(�tЕ��������z@�F��I�-��' Q�w-��D{���9���E��+��}${"}�M0�i���F�0!��g�,/m��K���Hs������6���A�(�KCǆ�����	�Kާ~�@C�vR	���C��}M���{�7Ԕ>�o�f���W�s���v��_�F� ��Q��S���C���ѿ�Vl�$C��x�WS�k�a�&�wʴ!a�L��T�R�}?H��Q�MUh
`��h�V1z�>���)��O��H�i�!�p���(I+�Ls��f�F&�C���u���i�Qb�{ ��2�6t14N?�S�y�}ڌ$����.2K��S��;�7�q�#1s	T�׹ٙW��X�fT(k�|����gZ��&r��o�8����,��.�)j�/"xp"DFl�K������Iv�d�#�{v1����#e%�`j�K�N}��;-V����L���I�E�\L}4 ��SHwf�YQ�����70k��+LB�8{ݳ�868���Ssn��ATm��(�7c[U��NH%�Y��9^"�i����U"x�j�����{����B;��eR�\.�Ux���N=����ד���M�]7�'sY����fz�eAM9b�����J����ϊ�Z&nK�' �BRp��܁�x���̷aG-�.�8t�9���I��+� n�c����ȽW?l��榿��W��z�ΒR��\מ"�G�Tt݁�t��_1z�F��"����,��-�(��S,� �B�U���0L�c�ګg�v1Zx�����I%�\<y.9Ŝ� ���[��2N�̖2�>w�}2�B����!	!�96/�D��kQ�P.-�Z:`�]���7
��O�k�i�{��w�_ʑ�p��1�C�`���[Z�Z����iCv� ʠ�R��zj�}9�R�r�E�cd�.�
�0�0n~�
+�:F�^q�Q��d-��0ƨo�Ѥ6�D��EMz(y+>zq��٥��H����<���Б`�>�X���0���g`ߒ\�I�g��߻=s!ճW��V8)i�7�G(>5��f.�XdcI5\!,,*�����(���D�Tt�$�o-�'����O0Tx�����I��,��[|��a׋��"�MB�aJ�G�����)-�n?�$�ןX%������q�)>����T��W��XH+�~i6"r1�*��Q���#�7�Y�K����i,F�mڂ�-6̴bNQ��������*R �E�}6/1,�����&��@Z��F3�B]bǅ�1&��oPT:�I
&�l��K$[�R����hJ��<��߷v�ٳ�i�R�XE�ě�k�W����-���'^tp��{x����2!��U_ڈ /�*��i�5��=d���ߐީ��A�̫6����Q�v�X���*����������u��%��\�k98��O��	������y�sþ&�Q����$}ҕ�3��i�
�ah�J�_���;�_浼:b�����3K�d+�x��$=v6�W���Ӊ� � �R���p��㩮Y�"����'���WR�}}{�{Q�9��������QwE�����
l�^\OI���L��)P_�`׈�����z���e�Uf/%V���oߥ�c�J�k�~�H8G>�t�)ʲ���B�ٗU���)��P���Y?{���-i�&����~��iR�K����?���� DЀ�4�%:苢qޣ���c���J��W}�6�'gK��ie:^&��X�����J�h���vWe���:U��vP�*�X��� �b<�[n
jE���	�4e��Z�2ʠ6�@�|��z��q�f(�����i�臺�\�������mw#f{XF���p���P�c�t�:ɘҝ�<(7)zf�G��W� i���#�b�L��$��}����#D�.�����zq�&7���j�X�}i �
��+���}G~n&Z��.���Cv�Mdj���/ͧG���r�K�����!���v�6P@�Uq��%.��������\���]<o&T(����	�`qTrL*�� 1x
?{l����=^�;'����K�7�����
^�s���� J{��(�}	[��	�Bk�^z
�;r�6-�t.)�X���f��q�9*�s��38�'��l\-��xvvWһ�%�����E�;���jffylRwM����t:P�Ȁ'�V,�9	<�����o�,�� \1�0��س�m�X���rW�2�A-�4j%<��� �P�t5fD�������Qم��)�e/C��F�<~#��r�l�A�*�Mo��S$u��z��
Ӟ�ea�aE:�1Ů���P�M�Je/�!RҀ���_���_���6�٩�!9��2R���N�����+.INnMؓ������dk�r�<>�&��-�RO��!(�>�{��
w^˖�ή��ܽ�9/nJ��y�_�G���'/�G����c��I;\o��|Lmj��Q� 7�UE��a���2�AnՐ��ήN7Т��FG��t��pi�b��c��<dHe
�����|4�(t�P딴�T	���߭�S�\��8(q����ғ�*��>J��l�MI+3z$8�C��s6��nII93��%�12���k�Tw-�y���Ңv�	W&
��Z��	�!K�V���-{-�~�w[yf8��*�z���p�Y�8��$F��2~�)�*�eC������~p�������i��#�W9�
h�V��$j���P�s4�}���c��D�P����n���/�X�f'��fu+�*{r�vs�q&�vF�孕��%�-p���[�+���d
k����ɪ�>:����7��c�7�)��ճ�$}/	ö}�����(�"�չ�*<������PC�#\�ki\}�+r��x�Qd�nF~)vk��\Lo��@�"ͱ�=yk�Cn[�˴��]��㶓 ^�s��7��`Q�w"p�=*imK���6ᜉ��6�{֡J}2�lzX1fv�ۋt#2��Tl17B-b�X[�/�N�K���\O��*�:;�2P���g����~��b��o5T�=��&�%]�v��߭yr���nP����%���yl����I���H��s#����a���5�S����bx�;���ǒch��tٵ5?Q���	&��=�0懏z���s3�nװ�S�#�5{!�F�Xv��t�vT��	�s�g��KY�$��~j�e�a�8�xf/+���{������B�~\����a��S&�;�K1$�%�ic ��� ����W�%���:+��k���U���n�8�9���EdI�f��伔F��$pst��9��|�AЂd���C�ZUJ"VUT���W�Agx,�_^n�1�S��#�q�b�|�5�hk��(������B��>���<�'�$��a}��ʸ;��\Db���@�;!I®�$E��9K.��#�yHĤ��T�Tm�.m�6{c;ۿh�|_�^5H�,�RB�kG�ͦ��5�4��{(�G������an�ͪ&N 2�/n���d��<77��\����S#?�e��
#����(]|��][�"�H]�P���mŨ��J�zD,�n�~��~>�h�(S�(���L=k�[0�Ht���ڦlᶥ��NO�}�G4�V�7t1W)�J�T���qv�cFí��m���r�gsNcݐ�5Sb�S��X��rkⰔ��_;]ɝ��y���5�3�+^s��>
,���r����}��<0�̀[kr����UK1�N\IT26��]FHN�_�2�"�!`d�HX�����nGox�z��9���Z��c�-�+ؔC��ǔ�?B�]ʊ��A���|ӊ���=�̏���ɝ�7�2��D��q�"d�5+3��Y��>��[�਴��U�Ϡ��#�6Ty�lF\/�����IV^�K3}jD��X�ݛnC�e=M_��UvIn�%
��)�V�����{�s���	��DE�]��^�?��<� ��7u�Ў�b/�-k-(V~}!�0�oW�#��	��u�DUx?_IE�OzUz�h� �g��3n�� ���..w�" :�4#�۰/�Z�L5�UQ�;H*)1�)K��Ud��-7���Ԟ�
�j�tB6l�wܾU:q���r�
-�h���W��QM�F� �3��zu����В�xy�
�>���J�I���Csݔ��]k�E.j�(�]a���:u�}V�z���S�o̞���[�jY�m<.��� >�I!�u��A`�+������MWT������åq+`Zw
�hA������#)@h�������"�������Pb1b�ߔ��>������9�qݣL�(H�9L4�g�pC�$d|܌d����zP�������G3�:��������Ҳ�/��y��|_�}�<|�ە����9�_���zʭ��'�Ja�-ٺ��#Q�H/�Y���P�	Z�^�\�hP��>vX{Q߉[�SJ��ʆ!�$T����&C`����K-*c�ړe:�6LI�����g�f@/�?e��������;+�S���i¾��qZ�Ƶ�;��	�u��ǖJ��^P7�WӀ� 7mbUˎ��l�;e��i��H��\7�o `@��j�:(vzm��f(�~���F7B;���ma����]���XI�UG8��*rj~�����c�A��8H�tO	�[ �C�
�7[!C�4eq��D����qm��2h$і斕>Q,]X1�p�y�3�`�gs9�)[�Z[A�D�Q�_ބ�!^s���N ���Z^��w_o:<�v_܄�!��x�vBK�S�}6b/��i��X�y�wmI�{TZj`9(Z�O�^#8�P��R��H9؟�+-U��+�%g���~�����}&.*j��;�y��_J3�d�eL�u|�*�O7���Y��>�+��G�K'�.9���7�,8��W����t��9��-�i� �H�OϾm\8"UٯD���N�#h-���U1A����u��8&�:n��Yo{�൵����-$�}�p��2�u�w��Xi��ǎ�B���ZK�k����Z]X|`:P�� M>Q	�%d�0']��vcjޚ�"h�ھg'���MZ�P[9#�zK�P
\��@��F��T�^ҡ|Č:�5�}�(�g���mz7�� ��.�3�k�~E�����i@��Y�7�M��G�9��D[LG��KS%ѣzGY�V����?t�Ք���s�a	>�o;m��ۖu�W��S'���*�b�����{P+�Ծ?+Z��]@��*xUJ)��3@��D��+@�4���h/|��l׏Y�)p�z���;#��L��|d���R�9�-	IO�KDg	�\��
��]\%��λ)�c>R���IɮQ�4�ڧ&�e�lE�$.� �S���(�9@��$� W�T)uH�*����4��39yn�#�h��ح�n�/Q^ n�����'0�u0m��HAiawd�?�.A	tJL�_�%E�\dF���Oy�Q�ެi`mͮMۭ-Q�O�9��ep�@�i�`�J�{M������:���b/������/?��`ך��0���y��SKg��B;��H{�1	ΦgC0"�DA^ˮ�p�F����X
m����f��4��E���y�\�v�J�-�M[���	јJ�%��)%6M����|��P�!AU�+�x���0c+�ގ�I;DU?��w��Ў��=�?z�>����]�7�j�n����/k��@3��L�˳��qv�zM�2����x�<�'���.�;�ψ+qS�'[��ꢧ���ê	{�͇d ����٦v��f!s`�����oƼ��u�a��1���|�I<��d��9��s��.z=��z��4E�����&_h���������+Wx�Pl	��'r�������j�?�F;d��o�jd�G-��:P4���'��tI�G��E�(Aq{r=�#�Vzc��4ء�]�+d�s\�J��R]ċ������{�}]�0]����r�[�@8��)᷑�Wq�Y��t�o~��F3��|����P?e��	�d��E.��m�����@�u��u���aE�"J�CTs��~>��R��{�U�(@+��`�ё��\���b{����z$��z��koǧ����	{A��t�/��6�,����w@���0n!�A�
Q�p($�`̄;�.�S|r�l�M���7��q�9�OS�@���������a�����G�P��K+?!ymy�A�-�p���1)a��q%�	�l�M��ĭE��8���Į:w8�t�������!B���6�qV�剞EY�����6�/����&1�� ��^{�sTS���DH�x�W�Kds=���G)�
MHH�\�����=~bz:{��؏�P*X�G�@��a&�"��Ըu�"v&�rn0u(d�����>���2�>�|���3P�]^z��M�/��f����|J�!&��_��Xr��:�u5@�z���|(�wug�~�7�`��;�C�.hvw!&��\k��n�wY��m��g��ɦ3ɴi��\?�4ѫ1�؝UAQ��#�`D�5�LS�k���w�B�A(��`�SJD����0"x� j`g�F́�+5�(�����0ɒ�7�I�tt����_ti,�/���y�xXq[�j�3��BH�����n�
��?,J�6�8篫����ܪ��$8��1!��5��7K�͜A�ЎվosI����ؠM��NX~����"d�fF�˭�hg/��o?�̈v�9�	{����ވ��Ю*���{�k�0Qk ���|��#f]�>,|��%�s��C�F��,�$P� S���6a���TZ
�3�������>D0�f���P�p$j�/�޹��\��Q�TTV���Wd�ƨ�A+�I����l���^�a��l��@��?��bL:\+�ܶj�a��s��e�B�옔B������Pږ{�IQd,yP�Ӄ���AF�_CCz\o\l��r����u�m�\y���I=�
|���:�t߭����o^ʻ7O��ߕ�5�|�F�R%0��7���٭G�gjW���ᔣ�:;)iJe����h�`sF���S�ɐzk}BD��C��E1��UR��k�ނ�|H�߻ɢϻF��2
[�C��#j^�:cD��ҶU�-3���AZJ,Ƣ	�)i���4&��P]�I�̸>���.D��bq �e'7��bK��J�H�fxM�@�C �Š`�Q�t�?s�#�R�?��zX����(6Zʝ���x��"���)S�Z�i���5�;!UV�ԍŉ`��?U����Y����G���-2��an&��;f0�i�w���iS�u����p�e6F���p�]�gX��:r�|k{ɠ��}>M�x�!��MŤ��JqI�=!l~ 59)6K�BXy;�se��$hԫ(�r2�����A#�`�k�y� ���C12�y���G�~)��xJw\"D\��Zx�)��E��+���:r�c��\�<���3K#�3z%�\\R�ȑ�����N�p�V�yBlX]�>U�����K���|����vc�����q����1eA��{ڔF�X����9%�v��Jbeu!�|[��7i��7��M��$� ��;����:|n��G�ӛw)Z�Wp��+'�-��C��{um�9����װH��S��~]b��[�s��8\1T�p��yG��B/n	�S6�*XkAKP����P�.�j��ٱ��K��q$��"U|~Ȃ�rf�"�Or��W
�᫋Y�%ae=��3z.�.1^c�U(9B�;�N��&����W������BE;o!�X=%SJ�g&�N�{A�ƹ��.��2�+��>]W��$GS��t��>��L{�5�2�Tq���C�̅�!����])įIKP(��|�E�q"�3�]x��~o@Q�F�21������y�.3O4H����>hD���<��g%��Gt�A�0[��#���ٹ��w�v��٩�H�e��qO�Y'(���P��n5N����
q�.���Z���g)!u���L|5Y��T�~]	�8*T�=��9��G�����	��-�oj��N8��0����y@���hц��J�W�]NvL��/���>���zR�[���t�i"��l����v���>vk�!3��[�����qV���M0-�=�Ni��˦�8L��!)����K{���v��+fb�q�5�b�J���"�I��fz'<M��ߑ8O�|�TU�7Gy��JR=�5�4�G�8�S�X��p�z/���t��$��Ľ4�����B���@?���������PU�咆�CR����rcPm| 5|�nM�{Ɇh
���u\��9%�����ײ$�8��m{O	UES�T�m�eI��! ��5��W)�������Й�t1�D�R���,�y}g{�������G��p���gF!h������^P��5'1{M^�(�`{�!�8����|S��ao��u�!��(�{�_�y�r0"�^7\%�,q����na��'�mk�2#d���N���3�>w ��9z�� �lq���O���|��bQ�]����w�^�pD�m���wAT���l�?�ڶIw#*��rc'��	���K5��
�����Nþ&���wi�n�z.��� �d��c;,0���tI���0�O�Ha7�0lf�����4R�>���6�UDOR+O	�ʸ���*��qѶ3kѐ�`ZD��I_��/0�K����Xsz�t�ˀ�,m~��c�|1�;,?�����9
;Ac,!\��&�/M�.h�da�͢�������_�x1*� �R:.M�F^���������RxWg#�Q-�����=��bM���e�N܈��yTC?�IY�����ɂ��;�Wh�7����#���/���&e��ש�/%e	���?<������e��;jZ�k!��E��`@�2Bn��m���w!�� l��C7���������� Q"��ڝ�Q�%�=M�ǭP�X�Z��N|��4�q�w?=:�?�n�0w��/Mxby�O�=�B��9�����^��%}�����W� 
���߳��k���4�zAޔ>?;?v1�Z���ѷ���v��V?�,��!߹DD���n��ʨ��ԗ���}��ʫ������z>��ݴ���] \��EnE�=9���J^V�7��%������F�	H���0)�0�wM��� M^����v�9��ER�zh���;E̵Cb��[�� N�Q o��7U���j�t�>IX��d����I6J���{C�� ��ȧ�h��T)�KQ��~]ɥ<���°�FКa�%q2ZFy�J�Ȱ��U�y���M��50Z��Q�P��_v���ȸN�c�A�C�K�{���?�x�fyR����R����Ѥ��[	|���q���W�\F�b=A�Z1Z�ѯ?+�$�ae��'�{�q�whAYR>�{�����8�3"���iQ��4v z\bbD �@���-��=�3R���ٙI��w����z���98A%������lA
|(��6�5�J��2�9.�%@q�@I�ѕ��$I��up4��׻��L�����uX��-�h3q�
y�v�GC1:<]�f��#�����ܱ�STM�m�3���6}mV��l��1���z�=u�X�N�yEbı[hW�~~��Y��,��v��̸�x�&]�����X�!�UA�/���Y�[!X����V�~'�gHHo2Sz���2�M����e^��Tڏ$����j)���YX�wp��E#�嚄�o�05?&7�s��3�A8j�{Ɋ��þ%BK�*���m�pE3:^�s�k�q��vj��>	q�S(KZ0�@����&�U���~%��:��pP�Qs�fn񊑓$������'SXBi�qO�~��;�z�X\�Nw���@5b����#�zd��(���7���*�OA@i�b��ЌQS>�|��*�����&�� ���&n�R�&����R��O�X=��𳒀  �����zWp�o��7!!`󎞱͐B\"E�(� ��o�%oGJ�-13�z��-�8B����R+�QN/��&o`c�U��!Q�DIC`!��I���Z>Um�xo(�Oe����wf��`�b �ݜ���xē���u���URá���ԭ�^r*Dd�	��̸�~�>=�����<�����V�����Fv%���n�G#v�f���B�gj&
d=���zQ1RM	���Nk�[�`I��>T��ִݶ:u�Vƽ�9�x��.�SHܩ����+*���# �s���������\f��fr��*������_K��+C"�I�	�gd�1V�A@^~�����NJD�&�f';�?B�qk�}[#+�	V`f�h���.�ma O$��A��F��*���0��]�1'2�I�>�|�\F2���E<q<-��0q�ro�p���zظG�D�BZ��R��ȵ�?	��ǫ���jV�N�����DEM�J�Z`��i�:���$(��i�LVx��g�{�_�h����$�5+�L�%�����U�'ِ%6oZV2��<2��j��d���w1�~_I�j��� h�d)G�����:���>��KP��J�M��ɶ�F�R=E^�� HT�i��I���m�V�_[-*��nJhJ���;a�� �p��mȔ�t��_LI)tJR��ӻ�(,�k�b�s�I�B���}�d��f����C��WrIk!���&� �O���.FD�=�Fo�����C��+3�c� ��UH��A�h1Ë*'E��c��Kus@k���f� �����HLЃo0��b��g�l)�!�d�;]����<�;��ꈕ|#����>�п�"$j�H��	{KA_.�w�|����\�[��!2/����?_ZƑtT�,*���)�af+�2�A��J�Q/��Yf'��bę���DC�z�r�uJ�>�Y��09��h�6UE8��Xщ�e\.$�P�&YI������C'� �%�ԧ��9%�&:�LN��Ī��ȕE��0���ĕ#�[�am]p_~�A�i��3�sO?�y}��s�\hϊYX}��/�q|	�O���辇�H*g-8�6b��"�i4�b�<ʪ}��@2��=�ټ1�e����1�����?}��_`���{"�H��P�"D�gf�{:��v0,4#��7�0�����*R~mm	�l�|�D^v=И����t��}+V߳���R�5]���xOda���jl,P��e$��OI
��kxA�;��9Z�C/�p]=㠗�I����{
�8�[�e�~��hP��΂���2��G;zKq�T5��F���'���~��@2����`C
�!jUmIԐ�iT_�G֍�J��	�����q5Ԯ�-aʼC���&���ij�۞�8�bhW0yg�Z��f����Cܱ����ڬ�X��֭:X��6�q�v/�*���k��Mž��]���Gx��3���b�y��8�륈�q�N��f��ǚ����-2t�XSms��H��nj?"H	e�b�9��(4JR�&}X�4�;������� �ͦ�O�3��
��^�;�E6ɧ�Z�τv&�k�g��Y��H�(�\�N�8�`R߼�;z���W�=EU4�2\vNeƻ���nA�	D�`m54̟ �4�WB_�N�ʆƆ�BU�+�O���C��cpOHb^Fp�����հ:��s�l=8'B���2(K��`c;ʝ�u���A����CTjmnu[���H�s4�pR�ĝK��04��m���i�2��𑋈aH�O��i:'�#^8�`��5v�Ր`�[HxfO�qƥ�K�4�+ �~Yʅ>����f��)����2���Ɯ�RM�]>��źo[XSf*�F*�r9_C�1�7��J{�뇵i����>E�]�ZM�C9�9�rI�=��b��o�	�B��A�m�bXyA\�8��M<�M������Z,{7w��d�#�Z������|�����"�Dc� �D��`��]r�-) ��@0�Ot�?ϕSĨr��
/F(�&��)��L��J��f�T!�QT���.iI��a[N���ЇOI��?\�D���,�)h轲v���4yd����.fU�|K�/܉�AY)u����l�fP�
=(�qz���Ӎ`�K��qiE|�&�J5���x;D��f!iu��W���Λ�x�c&�E��������3s�
����c.Vd�pp~�,��N���q��8*�Qgp~�
^;���T���m���重֐1d�
�*�vV�B(��`�U`�^�����R9�d������"�A	����OX�e-<�ە�Q��^��^�B�,�Vǒ���(R�S�$m�9 ���̞�<; �\1���1X����{r��_��a{�o�8����Kh����@�1��]�f�ۀ��G���₽@!8"�gQ��BH^�i+NA�}9E�\�8��#?���/���r�=p�A���k���&�O: �M�����0�SW����������,�O���\&��%�T�	�������6^_�S����$�������G1��i�z	ջғ�t����H���T�2u2�A�A�}cp�።c�J�yG�G��S�*�O�����~���t����[�b�^p��o8	�R������5~�_���ۖ&��� ���fɎ���`�(V��
��z*�F�\]�8 F���0?�8F��1�ל�6?d��N��E��9,�w�V����0�\Y6u}�E��1�6N#�6kY����zW\��j�u[{�0>bs�j��VE�*���4�*�������+�Y�ĿU��^�fS�y��� ���,���9�����;�g������+ۍ��6���\��9�>���|�1�D��(�5N��C ��A����eO��ӓ�|U=��x�\F��� 5���q�7�u�^������*�#��E��Eχ��S�#@
*�i:���d�igo�tȔxd���j�!'_�o��ZSZ�`E�-��sF9������U�T�%���ԥ���x�������V�J�w��$�)�IY�䎝�1�,�����M��mP��Uj�PO��62k��h��DO.㧐^�VY?�&D*�w�kg�f�n���{�܇%�p~җq��Qz~í�r���.�4���cV��%�m�f)��A���&I����\N��/�� L��H㝔�4��G�Z�!�qK3;���� ��l��r1޷�?��絠��.R(SC;3�kWUE�"M�[;���:X�Zg�hk��A��a�q֪ءX�ΪZ(i7�-�P��Q�8g�+9Ya�n�	7�������2Zq2��1���ҭ�Z�=A	{��gs�v��Ʊ�Z�J*yD�����Ui�?>�,��#���'x���}śrG�5���2¸Aй�F$*���a��v#D��#	p��V)7���o�J�(ؿ�#I���C癿H�-�{]�l��_`�L����<��&׊b=���I{F��}��F���_�c�7�]�x��RpN��*K�Cs5t��J��JBi�$�{����jb}0*��Y9���\������O�S!:��RA�E��0����S��Z��C"��s~� ��#A�3<�~�s���ȝk
hd-�����;��OGr�Ӡbe��Β9��X����������Z���<���)~g�3�`�.��Pڋ��獛(�*��E�}py9Kۉ��I4q�`�e������sEi�
�h��$Ͼ�Y��7�E��7��M'�n<�M�]5�Be�ܥ���Ý�b��ᾬ�XI�ШaӒ��־�X�Y@��3V*
�++�%eX���
>��5�Y���6�᝘c���^	�32��MJ��`���=��~*�f_����,#XgH_t*�,�p��ɣK'C��ZG�U���Pn>Z�A5LnGf�)ɦuS��~˺�?n&�0�5�yhO�-���"���. �o��)�"�	��,'/� v� Qui�	@���Z����r�+73�E2�{�spik�f~Ǿ��|V2/!?��H'�,[����X��@�5�bE���FIk�ce6�,���'�7:��m�[c"]�	_>���zs=��1A{9<�ٜru�� ���=����{�br��ƍ�D���o/Yf*)3�A_߭�	��v4�$r
�$��F>���� [`+t{�Bn��]�	�:w��6�ݦ������A�0l^J`Q-V9Z߇���Q��eY��y�?�l�(�$%:�%�����a�$�AnOE[=B��\J:��C4�lI��af L�u�A�;?��	x]J���g>�Eʮ]�1#���p�J\ࣺi�P�͍�>����/����/�U���QA��E9�1�}�F�r��c3�:YW��?����\I��4[��%*7���w.��2������m�3�XxB
��X���9�܋P9�������P/��O�D�=D���@	\ T�v��-\a��q"	+�n�_���;m0�1�Dh��v��7�=�̡�<^:_��U�W�{����>�K�߀���iJ4�|����/N4I���<&a��b�=�����[.}q\���(zQ�����@\�`m�-�h���g`�,��팖��%�:�gG�N%˪,n���I�$���uѹ�.\��b��|l�t�"�hl�j��ɯ�%������Jӧ�
�I�q�+P�h������/x��+/��G�$k_�/�sG.�7�a�F�Ki
]ش��cB�� =,��Atu�#&$���/�9��چK!�j;V�-!���%PWܬ�T�&�3e�K}�)!1?�*���
[�.����+y?��3kd��*!3�����3$o��OP4�}�wl�-�#��ޫ?}[x��cݎ�)�N/4@-n�U�LewH--�����N��Q�Hy$mP�ǘY/���W� �.Z���!܁b��^([�������/:�t��&?����b�3<ȦftW��$�3�F��Cm�ѲҙW@�P���C����5ѡ�ļA�j�
�S8	���z�U�L<���u���kRE<x�m�=�7�P���g���8h܆R���V]��j���?*:��ɯ���� ���j{�����󘻵U7�0�R
�U��ʈ��D`�"���D��L��t$��#�y'�'�0*����d��xU�@8s5��v��T��h������$�<�ּUj}���F�+"�r�E��q[Uws}�bk��t_�
��SK��g�
֘;�ݮ����(5Y�`�m�|_3i�G:;�Y x�s�1�~�xk26��	�s5rw�b2��5��dF?�q�jIn@�R6����Y)�U���k���pZ2a���PFynh��?�o���eW�,v�V�B�v��4�
�	�t���k�g����$�׶&/�K�ЄI�-cpW�q��]��*�8�t_qtl���1%(!�؄��i�6~�����E$-��t��)?kn���#�
͚��7S_%�R����>瞠#G�j��5��@��b�iu|δ�t�i�D'�m�9ӫ��
�,������K��Qb2�z:$������̎g+ #Z������J�O�Ɔ�-0���k5T���.��y��I�^�^>�I����C@']�Ra�c�:�jS�S�sK(����`���6I��2g����q?��|wr����R�8b���
=ׅ�+%��]St|:*@_�[��7hU٣�����8�k�����e��ע��5�\��-�r�<m#y�P�s�~�q^�}��`v�wLjْ�/�)�7�*�lK�v�~m��ٱ!{�7uP 0,(�N4W=W#?��S��(����2�L8
��Ŧ�ʂ��/���iٛwE�q%����ْ1$���K����F^���I�놄�w�6�/םs�"�k$6n#y��܀�ԛfw�s�%�=���i�3���u��i7n�v��~>lG���p��2���4�*���]����ɩ�X�h��KM�VB�TLQ���a����E�&��5i��VCh^:"�޳�2,���Vݣ�({`�B���G���!7��:_M���WF���Z<8��O��(��'��jZ{=e�:��K��h��:�?6��^��on ��������sq�NݼR����Uz��*S��u��n��r�2Y����ra.����L�·�P`�$��r�P��-���U�Q��x�`D��q����:�������t�y�C7߷ QY���͋hS�k�P#�4�T�g��� ��QD����X�{Uy:�/�j�6/F��1�vф�Y:a(\���yL�8H������㜺U�b����.�]�\���P=+�O�[�i�o��}nh��d��_a�$|��UH��؂��W}i)�9�%��U�r~�� 2Ʊ�a��04���ZÏ�4g���"R0�MF�$��ȴ:K^(2����R�nd.�1��덑9�&������d��zCW��y*�|ӱ�{~����1��C�פ�@�������uG3�#���t�n�wRB�C$���q]	�r�ή �5� [�9�H23�|�|����<;)�ߚd��e �:B�6@��j��|�w�&� ��b�E�����:k+�ب<e����P5����������D�4�p��S�|Wݰ@h��c斱lqJt���#�]�L�V����,�M��gj�S/��(�g�)��D@�FbЃ��п�qq܆Y[�
*� OxV�.��FI���8&쑸X��P� PK��ܥ09��Z�x�A����������l�_e��R�%���m{Vsb�e4�o�[\D%j�5�)3e\{��}��k��:f6�CD(>	~:;�	8��A��4B>:����Ρ����;;�m�q�/A�OE���\VU���u��K�6U�����7��.^�LZ��ץ��l����	�9w�L3̶H����-��74]���������y #�H���&�J�6n�3;��XUȒ_AC�!��-��|���m��ϔB���yޗ�8�ßԹN� HQZ^m��|�tB��z��V��[�tZ���i���+@�	�#l<�W�%!.E?qE9eZrM�|��V�Il��w}j7j�Z��Q�9�)3��l�4��Jp_h���?��H�޶�Q2�#0�m{jS��c�~�g�`�&���2���v���8řeD�<����(�2FK�P�5�ŋ�qD��~j�Y2�:�'�f:�mX�S��1��@�q7EvK�@Ó����I��rw��a���u��҄H6�v��r�b�JM�\�L�]D�4�Y�^�v�I��P�%��tU���Y��T��[;��s�g�6���t���"����7���4�ޗ���n��4
�]�`�ֆ����O��ǎ�;�V�\%��E�N3�03�<�!�Zw�Z�^6��un������
S*Ǐ�N=�`9*aX\�{���;��F;D8݃�2�=�voek��A{�$�8�.ݤk�YB|���3�0�+��Q'��#p�|�"%H]#;LV9�z��_U��g�n���D��+B�~�P䣬;O���T\�U��Ǣ�<m3�(FK�_LuE��h���vP�����M��|N�h�l1d�Cl?��.;��	�n�qW�s��24�� �E���m��H��l���;�%��S�Ձ������3f滕5��/u��R��ê�X��ebf��_^Z��7�g	��LX�N]�v���@�u�p��%7ċ�$�h�����J��+���-V4M~�X�XNAbp�E�w�N0_*@,ՠ _]�<�L=���_���٪O��=�E�e�.!��>(s׳�.��H}��e�ߗJ[����t��M�R�4��.�A���'���2����qɅ���,zp������cfq��n|�V���gmR��{�t�0߃+O��Bj]q"때D��H} H��PWI��e�Po�F�ѵ+��@��:�	'/v�%d~`�`���s��?�������FimW>	��}H#v;��q����<�f���,Q�Lr����6���0�۵CU��暥w�E�)�긾@4���
�S��MO��T�)��ؠП���Q3�p��j�D�b���CH���1v�_�lD����:s\W(�۩�̆+�l�11	g�h*}�f�/����Uja���^�f����8�K�dx�g�9�5�l�"4+����%���Bs:��ɶy��~@7� ����o�ߜN�����	Ś�Wm£�8슛
�)-8���¼��g@�H��Z7�lT[]�iL�oSs $I�A~.	���Ӟ��۞�H�%*o5��ݬ]�T,G������ K?j�Mp����{�s�l��B) ����X��~A�)3l0���%�	 K���G��fW?���ޒ�:��OOv���S ϘÌ�^6�>D�2�U��'�����8ȶ��$/�F,��n�mQ�6	7E����c�/!kp�Hө�B��t>�1��b:�w��ڀKܞ�����z���W����^7��t��aDy�ic�M%<#�DW�g�s�����BV�Ѩ/�����g�S���a�����|$�G?�r����P@J�����D��Al��z��7�u/mݻh�S]9b4�m�;SYp#��ɦ�0�m��3k�:+�5P���)pD
Om�ͽ�̙�^��l�`��}�X$_�&[&�kOT�ߐ`������vѠ���'�Y�Uì�>�q�k��uS�#� +8����/��Z����t��V���6Q@T��QE�64�S&�کk�4����)v��4�����k���`��<Op˭������V��>�{$^EC"#$��d��zE���)��=f�yI�U7((��կ��#e��[o��t�5iͷ8��W��&8��hV&��&�;�_d{�?l��p�'�A2Z��$�Ɵ���W�"
�+p�K!�@�^�ˤ.�*�=D�1�R	�r"=�Y,���s��xfTp(�/�N')�vj�%t����)Kڸ�������S6�s�Y���$#����X��ڝ���'��Ԟ@��o7�<C���ь~�Z���v��q�EXǇ�D���G�r�#o,8��BNh�Ѫ~��6�XH�x�'�4�Q���}9x>[�cⷘC�1�����\А����ֲ��6�-f�e�{�1U�6����5e�ǃ+f)�e*O�E�~�m�����YOQ$:��o�V���#�I����gbT֮ˈ��2}�I�u�2`m��+��<�����G��N��&���7����_ъq�,�,#re�t��ʘg��/�-��]$\�#�)����Q<Jh��'V��\K{g�v�hH(��	F}p}�)���"Xʻ�L�>U�a"[��Q�P��܎���ȻД�x� ����RQ��.�Keb�����l�,�Y KP-��ѽ�[����v��_����y��~�~��:�Y:�<p0��xmۜ��)/�}���0��~-�He4����2�?���V|~A�E��er?�������3�*�0���n*�F�%����{J���Bi����r���gv�*qbz0�V�r��lW=J�B�kkΔ��C������7�z�ȶ8�Pj|L��L�\\�Xܶ�j��M��9�*$�iI;������7Mm�u�E��L���NQ�'E/���uw]���8<0T��nB�L��*y��[	���A�y6�޳^��޳Ӆ��Ƨo�
�}�zV�|����d�o��Zݴ�!a�G��8+&�q��%{N�J��t�ȥR,s���*\�;ƴ&,��N��N`�Ա�e������N�".p�!GL�� �n��U&��!��ۖ�WH��Rt���6h�g"�XC|7-�Nu�ô�Y#y����[�9�����Z�2�' �,u��^��&|)��"�5jY[Ff�\S�����`Ξ��4�&r;=OF���߫[��
�P�H�� Q�d��|vYI9T'0Nҗ.S)�O�YV&�a����A��c9UT�y�u�*�'G͠C�
5��M������$�V?�J�)a�	F�;���EȨ��|a�T�g��.�p9>�_�A��C����^O����a�~>!���U�=0R����>�`8ٿ�褴���,-�8��R��ڐѰE�����9�k��>�ڴ�~�����d�a.��ao�"4M!�@�,�z�� ���/���������`��̔�s�f`e=�z��-�v���̓7����;K��$Fj)!*
Y��SZ?��u�&��[��UDE�d���H��ບ��۝&0"�[$GK	*N�`�m=���NM��_�}un�0R���>蛯�ʸÒ���!�ė
�n���R��٬��E�� ?0��`)���_�Z�Q�7
���j�cAj�Z��M8-pS���D�x�=k����x���>�ɐ�0���mNp6�7j���f��c���,�栶�9��X�:�-t	.|�(�Aey���?�J����	��Df ����g��֢e�T��9�V���[�a��U��e}����*����4y���]��D�m'��S� �6�r>��ZHK5m:� �f�"w�,E��d�P���x�LM�#P�mm$�|�3�]�J3���!�.������1�Rjw�+��y�C�;{|[�Z��Kݝu���U���aA���'�kCW�ӈ?�,n.~z�����.w�p2��}��ҫG�=��t��ɏF�ymLaj4��,�ţ1��娧Æ��i��}��}��m��!�lno�Yp>hƋ9ͷ(�h�7"Y�w�Ct��&��>��.���j���H�s�lل��I�(��c}��K�#����Cl�c��U��U��E&V��W�I|jщ{��)�M6��3�N���l;���/�W�>�h&d��K�������z��l� '�n�r�yӥEO,},+@S�h����وG�E�R���/��<w8=@���.t�p�DV�����L�l�ꊶ����;���Vm��'E����G���'/y� ����1�-jK:�CwZ�z�t�@��e���T�l����/�~DR˙�x��k�m%�0��>՜A��/��
��6$����VPS�s�⿏C��|6O�s�,��]����q��I���\H����8��
��ob~������gXd�Jh���$!����^��d����,�`��fU����Kd�k2���M|\2��J̣
��Z�;n�p¹�t/�=���yu)5���WBT{�g5TD_Y��#�@豯@��4=-��,�(�.ア�B��8���(�[n�E�UaJߪ�<�Nh��ڱ�.�ˠA��k"]���B�`��(`���Le������>�@2p����CC�yF�F�?X���EVX��m��@:T����Y���U�Vy�����l��"L?՛ј�d�o��֒=��8$��}�G U��$�mrF$,�@у��#�E�$�s���m���TպK�6����5Mm6���P��K�h�	�*l�`���!���l�[�TYW�4x���,V�x���r. �����E�9���[�7��U�N�K�����xd@����廴G���" ݿ�I�Jq�:��z[���#f���ʒ�$������b�H`�;�ٵ�~)3>T+D#���ye�w,��a���4l �'E	/�}"�N���F����-+�?�#�*�RJ
�k�ST��Bv�X�;�*������6 ��'����gFk��Ouë&��"ү�,S	����KO�uc�̊u ǃ˒��&�kw'��� U�:�ʱxk�O�C۞(0%b������Q_A��r��/4s�^�����	��h7��r�q2C0&qdPPb*�2�[���##�L�i�
q�h`�#)/��qB����ҳ��	�������h'#�/�X�:�Ϭ�6�}eʞ0"N�#۷�E����1������z�d@4�c��'�ͭA{�j>Ga�0�	�~��4RT̽
��1��ķ�2�ǅ(J�2�J�M���	�r�f�4�>j��j�j�G�.�s9GL��'O�RsU����U9���9���9:��6�ˣ{e�E�0_~�>���>������+��Լ��ｨ��(��yl�c#�c�F�"��GlVפܚ�5�i�ȷ�)�������E��U���w��6��!v�^ÚɾL%Fc��/.��΁Bw�nJNU�6M�Rs��]WO�G��gC�g�~���\��2|;��$�t�/=@@���'o U ^�6�Z��اMX �k�B��M���*�u*8M��;p��ሇ��G�đ	�n1P��%��q��0��ɍW-vÂ���8�*���.�JM�v��;��6{S���h�G��	UN�X#f��֢oKk�@�W#���hcb�o�<^�3tS��t�P6�'�WG���{ܳ��Ľ]�0���aδ�i+� �~�@�S�9Y�դ����i�n�M�ά����}��X�v��P'��h�h�>��bϚ2|��DU��ˬ�CAM�Z1�#�N�f*��\��F��zm��7�T�h�/�Y��(?����J��ǂ��"Jk���GJ3��Nn-�E�9�N3Z�9Xil�5-��iw��������"YI�����Օ�|��T[�����C�Qh���]�+It|����ܕ^��04��*�,��\$�mT�Z��^V�Ȃ c�<���&���b�ޑ��Q�a��
i��p؟?B};Bz��������d8Wv�J�7Í&����Y��N��hS)6�Sp�mU=�a~F�����h��!���Kr,o�n5��0OX	6��v,=�
���`\����������!�+O�6��w\%c��08�9]/�!����3�w�q�Hv�u�������)/�fH�y#�sŸ��D�{��O�@2�e�F�-yф0L�U�jd��`^v^��VU�$6���m���E�'�uD�[vi��St�:m�HHG�F��T�8"����?�¤�B7+�D��3?��p�9�G6E��3'�K~��$V��uW �ƽ����"K<��t�]�dr�����8���-��B�������k��	mB�����q��&��xP�: ��X7xhb�H2�9���x��&�tg6�;��$�<գ�oI��o��gs�$q^O,;��K���N�Fv|S�5�qU2|�d6)��h���~��ag\F��{�s��e�:��l\��T0�N9+���/3@�Zpĺ��J�4˭�%O�86',#{�Ҧ�hȨ��.j��3$���X��v�����4���ϋ����{`���&�z�X�r��Y#�>,�8����ð=m3A����y��A2������	�0��+9)*��'Y>؎�׆��]�ЌPP?LBpn�q�p� �vJ�wr�����+;���"����^R�\Z�Ac�餎Gu�q�fb��z9�g�G��������O�@^5)t`I 6݂f�=J�I��1�tA�*1e���dA�7A�fZ����$�,RIr�}��e:D����M�frg�k��L��i�)���nR�-&�z��������Y�*O�X�ݏ�	�<W�	�rN��~�E��e��x<?�ogd8 ��O}j��k�l��@Z�i����,�Bp��Kާ�ih6��C�00WvYI���R<�DtJ��+� <"��"�	�)�fiٛq�X�^ζǯ'T_2+6�j;OD�pD�T�Ԃ{p��#�2�_;t��szfC�9�@�\(��m-3��m�i��H�b��T��g��	����P
��6)�9E�y�:��J��"��q|����~��eU�U��d�Q2Lޢa!�@ۯ��֜��ܓ�8"�|��w�$'JG)��j����<�TO�
	9,q(@x6�rA�TW��vd~4�`�3j�����Lk#l�O�D���)Ç	���Nx�d�D�I�J����3U?J�A`����{F��˴�빳��C�F��S�#���2`@Ç�����'��.�&����S{��ɣ	�>qb��CdY��d�C�+���n���?�)�W�!�tkr�(ɡG�'L!&��G���]aL;�9���fX��ܰ�
��`��y�;�%;qx�975Ab�
<K7��w�1�r���Ma����L����a���PO֤D7�XK�$~aN�m�*�R(�
��.r��q�W��Lf�I�X13�c�y��G��0�x�?jrq�:����G���;߹M��JQ;t�	�v�,�Kl���={k�x�y7����Oޱ8M��M�A�a�^	{͇���q���G6G�5���f���s�窱���Z�M�c�Y�Oz�9v��p�17b�3�Q=R��6o�ݖ͉P*�=���?1���&"�k�U�md�_^_5��-Kϑ���!P��PɟO�a8)[x�V�Y���mЕ�W�~bN']�4H"=W�����Lg�ho��+3o"��K�,O����BWZ.�ى�i3�2��Lg�G�����B���c��J��G�ϖ��ܼjg��wDt�m�>ʀ����5f��[��?��7P�f��7Ee]S�I�?��E=��R�?g:ٲ�V�|.�C�i �����ތ��������3*q�<��Mz����4�m�����}�aCێSM�����pH�|�2i�W�6;����K�����'�%\#���}!WI���Q�O�	c���t��
�Y�-S�����2����`Ţ����K���l����ĭ���j�<5M�쉇���t#��}<����ğHH�KF;����$3�=���;�o��|�
1�^s�6��᠆L����,����[BWw�Û�2��bm9ꅥ�[��ǽ5�!>\�n��!��.<���9)�B�#� 2����h�<�.�\ �Mt�9������G�n!~P&���k�r��C%���3�Øh��Zs,u��E�]a�hv�䠅�����'�7�j�#K�i%y���FGa��U��1y7����t=S1�������}�U��3OF��Ԓ]�I�PL�(X�Q�Y{Ƿ�W٤�r�����	�\n_�2�;��J�,p0���>2����6�b���]/��%�@m���y�P]�dhX ��E�L��So���'� � �"(̕+�TUդ�����t�|"�����a`E�졩av����kyNO�W7�1��p��L{��G	'Y���w]9XC�����h�� �!ikx��uR�'�L�L=�-���[�S<����(A�?M��A�)Y���Z/�D��x�щ���`�SM� F<8E��^��	�0�(�[��]��������h{�+� �3t��{d9W)y��+P�*��5�<�ë�Z'= ��n��]$�?��C�!�y~s(���6Fe���T�/NQ�5'd"�i��w�w *��@" ����6��������Y��k �?ZR�!���!������pV��B����~��<,���s��e�Wuf��ω���:C��Z�Ur��╄�x�@s�aF��x�#�T�=܍Q~!�@��ٓߒ#.�
Y6jB6ҊV���P�b�n<���m�b���n��qd��F6q�Y}��b�LX+��Ɋx���>�3�	��{K���J�+2�|F���ە+�`�m�T�,'�g�@��W��W���Q����O���a
]���D��������|]��13�a�3����o�NlV��L���b��M����t�����۽�}��y�����ת�?1�������m��s��j([�s��ت����6�o�2�x�lwn�J�fؙ��CnW��Z��U�o%F�C�%���+������O*�?]([�o./��ȠB��Ǖ��x�|�J(�.���@YE�M�:�`<FZ�o@�Ln�{�"F��HSh�J�S_D+<���~8��.�)�*K��'��=vbdx�����I��_�q歚��B�Q��$��oi��;�h�N�]�Z��7� �mj���ԙ%�pGQ�ص�\�������3Pa��S�#�OIԬ�.D~㘼$�͕s|:�P�[_A��w~�e|*�c�CP��8/�R0)�Ne�2��Q�]���Y�����?-���B�I�&�����=�4���M���#V�mH�*�Kz`2�"�y��ȶ���/d׬���!�d��7���/��F1)�ޯ��|@֙��Ե�N���J���2j��2�����Vٺ/�N4c���T�r&�_�x���ئ2�$xC~�/k	/����n��7��D��%�k��5�P�gD=a2Ȣ��� fG�,K]�>V��n������X�J��b^(�0G$/��t_�Uz}b����?z�}j�$�@���ɋ�2��ۿ����8�m�����r����4��X�Ћ�UdC|h����Y��{���	���F�8����䧉��GZ
M2�Ǯ+(�wݝ��b8�^�x�y���fz� s��1@��Д�M�fHD��g��1�r��I&��B<�\5��8������k�] ��~��!�$rv�����gOl<�a���ٵ^+��0�~lyi��q����oa�
L���?򨸍2��˦c�0В��%43M����`댠_��Zu5�]�Riޜ ��SP�"iyKZ�M1X��Pd�>`�|I|���p�Ś��X9�N$S�ڠq�8βC?��O��­lW�;����	Y��y�-ڳ�o�o�G�|<Z��w6���3��G �mҭ�ZA.��xG��fӶ�Sķ�xr�6��2�7;�B�#t��/�xfaV�zkg�ڲ��
�^ j���תC��Z?&��Yl�_�~6��'ם�xޡR�9���\{�TC,���do��X�A��*�1��J\�ېOD�,���E�T����:�͆԰t�{%��nר��D*�� 1:0m��>��Dv� 6%ʯ��]�<���]��q6_���EU�⒯�c���P�Dة�O��!�-���j�w�����
�s��?�\�(���vQ�f�,�wƞ�e]N�4�{xp��d�S����a +��L���֏�#E�m�1|叨J��#i�\��)�����Pyl'����+�A���N0�:�
�#��у$�w @X)��qha
c�3�a��59v;�8tga���[kX}Ks��${�5�F[��
H
!��zG��q�	d9I0k�6%��%�`2Mr��!B��RV��ft�|�\�d��n�0Pi��CPCY��X �(�M)��̠.e(�Q�0^Gb��i/��%ƕ��zƹ?�"癳/�I�&�[\��c�zS58�,ȟY[�+�s���r�J����B
��0s���부+�����S ��'u��ʥѐ�nu���� %B�z���NiU�f�J`Ex�p�2E�mw\�}��k����3��ui��tL��a��Γ�!lg@��-�k����Z���>�I��E}]C�#CT@�`�~P�2sz�G��s�7�]���ö�۾ӣ|QHt��L<��J#��B»פ���Z{���;'K��71m�R�sU���
]��d!10�&��x̀�R��hm�d�S{yu�3D=���Ib+�]�L�S��l,�gF֤[����t,���#����hz�ʔ*m^w�O�G�P��/AC�����K������0��r*�S��[w����ϑC��h�=�#�R��9B�%L�N��#���o�?�8Q��k�ꎂ�Z���<�g��7����8S喕�;�?���`�*︿���K�Ij
�mG�o 7B҄�j�i���h�כV&��*�K�OAQ�%�P�み����3��[7��)uXH���w�#�=��N����:�F{��$�SJ�;�@�1R����e��D)��b$����È��$xO�d�%��Y�� l(���r��:�YXNHԣ��������5�� A�1�÷]�FRy�NX�-�K],��ȷ�ܲ���f���*~�rЋBp�;�����!�<���]C�#�d��\~{�XakOD�lB�<�de�巼�)y����ֆ8���g�P�R,ݛ?�>�y�(q��h�U���{2k�2���齱1d��ƹP���|I�(Q���n��~hD#���å'�^C�92��K`"�%^����4�Mwif�X� ϖ��+����'��-)�3�C75���^9��F�[齶�LW&֚�"^�=�F!�CU5��aC��Q��w!��ئ�Gޠ�u�m�}"Q���S�t�ݥEx��� ��S�@����4�LOo:�BC<�(H��3f	�y*���͌M0�g��aJ��F�u�U�0|T:�*����ע*Q[P%8�?��)|�)r��«���	��ה�/~p��#!ؙ5C�y$�%�W��&��Tb���d�-5in�&���斚ހ�Ϝ煯Ma�J?�Op�ý��/}̚ab�̥~��.W�BtOa�.����Ee}�B+�hD;���B�
F��]~�x�]�kq��Y(�~\��u��^�7��Hp_���6�EE<]�%е0�JGC܇�!in����2m͸؅(:�������2��'�F�]��#Hᕙ��S1�Uu��Ǝ
���(��p�!�R��ד������9�̞���!�ر���1g�6pS&�!(i/C�!��e����;@�T�[D������� 1����!3R-���/�_�����Gkp�O�ﰎ��P��y{L%��� -�<I�����6�w)��Ѱ��Bf�jÊ��;z�@�ro��r`C~k�R��J����kÀ��S�+L2rC.�bPz|���d4�"1Á�V�C^{�`�ź��Na��9@��y��r�ƿUi�?<筚x��������ؿ`�e6]����EY�TT>�������d%kSҪm��c?��`E�f^S�0-<L��[�z�1	�	ȯR!���t�W:�2C������h��~:����/ί������Y�^�!�m���L��F?j�1de�-}��T\�	+�-���h�u�	���d�AJ;�;u����2U�|���U�����[+XZ{o�}�J/�i�ob�(AF�h��C�!�q������-�DU�%�G9�Z�5Y��Ű}M�K	��xГɢ@��+砛���l�*��>{���l@ :�f�������Oy��Xka��(�0��x���J�����t-�Q�'������z�!��v��Bt)�!fp�4��d<΍G���m6�SA@?�nj(���<]?��Ԙy���5g�2���홁���4(��Z�h ]���Wd�l<��Y�\u���_x�H�o���K*L��CB����(jz��Xֲ��M"�KZ�F������t#�~�@��
��X��:Tp&G�Ё!h*�z�>�'�,��}~��y��5� s:Ŭ9%�f�t�J|M�\� ��+վ~�!���w�R��`k
y>ܭ������n���Bj&=q9�s��.'�tH���^�[:/�����^!q�GN�[�G��v�f}p��ΗI��*VQi�u��w�����^��uVT[��e�7Z�B"��(
�8A��=>$�X��, ��P��v</��z"���}P�ܚ����IQ=���Mn��`��^+����0R#]�h�t ْ��� :bo�FS`F�$U����^A�I�{����r��?��+�D����}Q�9�h���;���%��TԚG�8Gi0���^{�#�_�&48�G8���~@s��n(�e� �j~�9��	�m&;��`��>J?�`ͩ��Z���2l@����?Z�P7a���tT�)ćbJ��= {����(t�Jk]AW@���U�8��u�gV���%�p�	�_p�gF��_��T'1��̒����k+)��v��0���u�o	�8Q���.�t0Q�������G)�0'��Q�"mvΧ����l.,��<�hIt9���6�dr�3Ӿ��4k`���h%��\��4�4�]����}6�f���m�O�p��cA%�c��(<_�&A\P~��
\��V��/#�$7	!�`��E()���6t��4���]��G�A��F���|������}o6��E��~��V�r"(&W�|?>;���Y�qy�*A���&]��<�m��T����OVDj[F	&I���?�W�d���@�����e])r*/�a���.4!��	��#}��e��5��X_�ޫ�����+{��dz9(2�A��Iz��wqm�kh���z%���Cڄ��
k�6�t����5��ۥ��q;�M]����«�7�1��Ӳ/+��a$ �v�E�*t�p��.���,�������M�����aL�ܛn�)�d�yꙍ�5�oW{F�_)Ŵ붠�Ȋh���G���-������.]�q������@�����H��d���.�2��mD���ru�+���^B�D���� �B�l�1K���*tKV2��<젿�{SRd��]�*�w��@�ل��4����xE4�P1tܾ�(^j���F�
�ݨH���Յc�V| 2,���C�4��L�Z��������8��S*Q:3�c�v���a����a�S���kyJ~'Ȥ�1,TI[A�Z�a^��JfLl�T�"�!Yap��Ul�#m$;v!��L�!>�x.w2B�6R�ä~�D7o�a;�J.3gjէ�Ո[���Íѕ�v�Mh��{��e����wΗ0?��)�����ũ)4��E%:/"�W;$i��-ͣkT;�Ĩ+��k�
ê���a�����O	?Wl�N��x�4ˍq�b��ck�?оH[uA���Y%��@���fB�� ��Fg��W�\��ڧ�:�Y��)�SK���X�+�<�z��OG��.���� �A�0�϶"�]��1VV���o'�R^FDN����)�2/�d�����	+�r�w7N�J+4�S��^GY#KhG*M,p��:��.]�z�j❽�Ŕ�l��jck�TmYs���g{�L�P��Ƹ��LiN�hA�ᩰɚ� _��A��1+��[������!�v�@`�7Cvm�Ft�Eki3��gr|(;`�HHh/A�w����:� uU:U;)�Sc�a ��g���|�B0�Snt�RQR�!�䇆uxe(�(�B9 ��
�l���1xC�fx�/�8���q;N�WLtEe͆�杯�$��H�-qz�U��*L��"(�Mv�B�谆�C�B��F�N�Bk%ƁXs�]2��6�7Eyl����`��t��M?kK��X߹�V��֬��`h�^����5;Ub�G��8.��hu^v<E&�s͙� `!'���}��$���I �������D���(�*��}��;������������:\���f�py��j4/���,��� �Þ�F�˿��+�~�?XkA�,,�����/ڔ��a	}q�Rh����t�s.�:��'��9���j�qh�v��Z�%T�f�������Q7 ������1@�逭�g�>�B�T6����Rfo]���p�cg�[&DS%�{ǧ���V��rCc3���^�j`[��f����2�U&Zld;�Qb�*��4ϙ�ͱ�O�4����R]t�ȩk�����	��౶���d�'�[��� ��u�./Q[����]�Ⱥщ^#v�SR��<���'��O�a�M�|��8J��3/�	�Ua{�����'�2�� UH=B�׉����% ��iD:}i1s�^4���j9������ug��?=Z�Q~�&�i� >�Z����D5n�:������\��W�����4����N�#�������Ʃ�^�OHL6�Y^�r�5�fzD����,��'`����Vi�W�>yL+l��^8X-�g
g�L�0F��2K�!o���Xp�b W�%���*��;�7�9J"@�[Z~U@�}9��I믧;��P�P��qC�X�*G����;�ܑ����CX��i��UEs�t<�o�0��d=�/���D�I�ۿF���)f�
y����ا��\(X�B�Tn�7�AWvb��n�h$}�߰E�:C�jF���KCG����0lX� ��+8���x�'�]����ޤ�?I��3
��":d#��fʀ+�]��yќ%˫3�"�h>���X�+��s�sS����Urbo���؟��Q����p���зy6^ZT�c\[��9��U�e���ylt�h�F`��̇�K��e���0��\3�Vv�篤V�Z�Ⱦ���9��vwA�����Mm˔����|W�����
�#K=�3�}l��c���h�tb�
��sz'�/�mh�_C�ۃhLSs7�+�=4�l��f�X8�F��!�����Z�����?l�?̋���ܶ�~������\a΀[=����E.�6��@A;/��'SX�ug���/W;�PdD�P�W,Q��m��7zd�����ޔN�wԅ5�V:$[����~�ҒP�V��w�j���e��ծ�L���ӥw8�UԽ���e3A|�S���l�w!G֙l]C7�� b���~�7ED�pp1�K���b�ݲ������k�.���[;i����a�i�O����{O�e�'2;���!�dG7\�������==~G������S*]��Ca5��+�A�%�|MУ!�b�gݚ��;��LY^�����Fl���D�@�BO��0�թY&H�Y"���`dwvk��1����o���_�����i�=���l*:�Σp�%O]Fėm��i��ߊӴzП��}�h��w�G��w  u�RC;i]�EE݌�n}_�X����H;�?6�;�Z2�_�i���y��w��#ן�	w>7c�*���%��	
�"��I|4��J�Q�FR�F�g�A ;��N�!��0�u���&��;�V�m���]Y<m��RdJY��z	�7ۡ�mj2Ҿc��|`ֿ��7��z]��.��?�b�Mn J�56l[O�*~-'��8r/:�aW�.�8H��|%	�lB�d2	Ц��e&2g��=��SS�(q9s	}�/ï��n^���/LЈ�/��dK��5?�u�o�DP�Nd�����n#w5W)��-���08x�\TX>�1RG�'�� ��L۝�����;`����2��f�>\�egN��R ��x�քTy�A��Q3������RS_�ZV�?�jjl����|*+��N�����;nǐ���3c-(��|SF�RR⳪�PA�8p���-�,<��a��	�,�y8��T� � ;�ʏ��"��4�~iv6�ղ%����]���O�9�
w>���`��1|魔��t� z���U,��I��[�+��՜�b��?r��'��/PNf@��Yս�wI�%)��[ڢ���tX�o����M�(��rO��pS�ߞ��^Za8�� � ���)4'Lw�gÚ����Tw]q���	�΃�&>�M�ٌ��c��)T'	�k�\ƙ�����I�����I?W-�!8��?�b����i�g��Qf�ޔ�������;SZ3�I? �p:y�=�^̅�Hd?S�Κot��i�B��6T§w�M��-�b�4�N`=��%´�B���Ѽ�
+Ӟ�i)0��R%�������lE���z�G���,�{�Z"p�"�\�-g9�K� D�[>�
��,M|Q�'��ɦWdx�V���O�� t�0��W�����N:�d�GG�VN�`��B�VezR,6"�¦��5��Á��&�	yf�ũT��@�,}������1�X���NV�&�H*ݼ���v)�*н�]!x�7.J#Mh����h�� ��Ӳ|�ɮQ��BWy�y�3�~C#*�m�n��r�A9�4}��|ᵣ9�zM�d>�iP��GN7�	(M*�:����,�>
���,�Ł�/�̬y��lp�kY�o:|,�.156�`d(h*����)%q*�/YL���x 7S��h�^��++�����NW�@�=W�ӄH�ES�?,�݀�,��5��`.���*��A`����RJ�ٖ�|��ف��������)�A?I�Ըʎ��w����E'�r����@乥�Q���T"�������r�f�"��l�X�u�Ց`�"7H4��U_	o�`	�a�K:;�1;�0X�N�Zb�����JӺ$�2������ޘ��>c.��_A��:~�2P�F�%j�����0��lq^�'�{��>��X@����/��T.�}t�gWs�m4�W���w̭v��bҪ� j�)��)8s��]�r�=�p�lEu���E�=��l�n/�N���ll�Wv�Ѳ��I%1���3�K�[0'X����j�0<4cKk3���6��E�a��?�,�Wm\'�ut�L�l7��\�+�b����=`af�~k���%��߬mD�K�����Ii�'�ݑg(Oi,a�@�Љ:�v��b��N]�b��Bv�.>�?��rc�U���|����l���ɉ�B�ej�%(ʗ~h0QIh�Z҅�[�`�u���G(��At�q��po�L��O�|�P΃7�]��}+&�UI ��� ��z��mB�a6���:��ő�e]xB��4z!>�m��,$�wy��A	Y,*�$76K�vKA�D�BP^{���J�-
��pR�uا���g}�4X���p?X�lڞY����������2+x��j�	m���D;�w������>${z������$2Ff���' �����0�i��A�v BX���YZ!l�wT�� �����C�5dj��&+�"G@�����/e�T���t b�%$$�_�mˏN�Ԣ�F>�,�� �UQ�����Q�Ĝ:w�9��9~n>N�|�r�T�:D�6I���D�W΂�$`jU���c�\�@�9 �7��ɂ���<�O��4�Z���
;T����E	���ۢX�}\��$��L��<�����ՎaK�.�b�{5�yv��>���$���ih�!fkq�[�=i�D �KȚs���o����NÔ=�:j���R����\A�'���Ln��	o��e�:IV0�f눀UC��K�@��5����Fn��\�6I1n�k�H�1G��[1֊&�܌^�ʥ(1��Z��8ڦLz�\�((�+7EM����ME*�����8�˪����qѿ�k\�)�����v[͘�jX��Ė��� ���$ԭw��K�:�]��oȜ�:�G�Nz���:�
�L#��� �j`a���ZeC��J��H �i��%R�2B�J��GFd��n��������W^��A�����6;�T����e�SZ��+�A���(���g� j�c���A��v����������cN�JخI��2K ?4��q1nH��:�&0�K`���	ϻ��������J�!��y�sI@�C�~�]�p�Mp�v/���d�@m�R��_��r�kU��%h�
�P�x;���kȣ�5��)7�)�:�M��wN�{%d���*��;�KϤ���0���{e�H=	��B��A�t+t1��I�O�B��5��d_ ��o�Vߓ\��_��=��4�T=}%X�/���Ʋ�b{x&�@���E�ޢP��^�UQ��v�((,DZ'ADs���.��.����7����Z�H
A)OG��9�]X.�b�o�*����!0�~�$�2;���xRT������T��CA5��F�lĎ��s���O�[Y�6��r�?��������w�qW�Ř���2+`[l��8y�a�ŪdE�i��%��J\o��+Gڞ���9����<���kd*��򭩫]/��9�*�?���`�1T^UEI��G�G������k��BfQ�i�����Na��9�yh͕��w$��Y ���I�K[�����Ya�9oUi���~�R�t�*G�R=3���b���n3\֣*o��2]�r"��j��[�Z�����d䰮)����v�8���0�MV�܁����k��"������q[m]ه]��	�-�����fL��[�P@y�����g�G��+;�4f��
t�]f%J�D�R�'*vk-����)G ��r*�
3��&����]�{!¥$o�n#l�8�:�0ʥ�4f���6`�s�5҅/�H`���~ȡ�|����Qٙ�َ+:��a�I\���D�k����_�/�c�Ѧ���h�ZT�[WY��a���Y�ɡ����n�t&uILz��C��O�#�&����\��AtD���=xI�XQS�Tys2 -�D�AP�3w�x˚@-~u�y-b�@�����WK!�7y{�2�F���0�].W%d�s�A�\�J�Њ�<���w��II������Ȯi�݄ɰ�ڜ@H�����å#\���YdR�Fw�$�ؒM,�E���c3֛�@V�[~����aT�>	�K���__��U�}�I�����SXL��r�D�ʢ���$G�g͕
����Ly�3kݧ����,�r�By�4���%�n*'vƓ�
�7���w�Y�pC��	��_A5�P,���}�D�p�DZ�M�b�����莔�pDC'��P�!-���/��&�G��O �_��L����"��6�y�-���Q��e�l��Wv9�6w�G����E.��j>j�PW��17���`o
�<�����*�NNO�<�z�:+=��4�ش��R��6E���fΉA*��=���V���[����N���H7Y��Ob�y��*�W�B\�R�Mfc\K�Z�J��z���H���>���I�;b��3}nT��zz8.���(&���6*B�����kБJ������W�K���(9r�����h�2Z�S�d�������9������A\,�h�=]���'��+�xJ��h��b�Xg$M��Q�>�g��,���\�ي�i�]�R�Hm�7t��J�˪kJ�Tbޏ܌ �}S�w)�eѭ�ö����g0D >�*�N����>��sn����G��{��m/���"��\{�����)qZu)S1B�����I��w�qx�z�.O�>�Fh��l�&�{L������1�B�P��r�e�=����T=X�t[�%�L���G� 3�?�=�?K���#�eÆ�Mp�z���i�����QX)ys�݇����?2��.%�
7�8�o�A�^TŒ�3�����;��h6�hӄm�ҟzҭ�wRtj�I<�K���x[�	��>/��=T�-��*�r��W?��� x�����A4.Ԟ��o�����.=��N�?�^�=�v�Q�W�X�rv���W��I�}M�/�b�I��]='z�l�Q7���=v���צ1a��)�,�X~jZ�&��7�L}O���{����~R!��r�Y�� �o��3����]$��-��/��U�NaT�T����@7&��
1A ���B��A��u�Μ30j���n��ޕ����[6���F�Rì����̣��lڀ�説��(���Dw0a�(��Db"��!h~uu����j(�$PF��	����Z~�K� �����/���\bDA���$��5�v�>l��p��.Y]O%���q7�7s�#	��"Sp�c׮�UM^r��)Y�f���0
�� "s[H�FX]D�+U�տ��Lϡ��sg�1��tK��S;�i�'/�� )�K�4��\���lJ-/�u�vY��sH��/��,�_\��i6uF�a'��}�ؠ|���e���?"uuJTޣ;��*��]s���o�*�F
�1�$���o�E��0�f�	l��N�u��	���p�uc��,D�L�����Kh[������}2&D�@D��dj��5
렯��3�@�<T��MkZ�<+�ި���<Dd(�(��������<�F��d�t�>Zl5t����q�/��1/�O�D쯃���)����>�-���<)���v"�a?d8��u.,a]�	�@� vӵ@Z��|�[���U�gf�t��u�tZ�Zt�l!C���Q��ݔ�3H-RԒ�$)6Pu$�9d ��儧���y�8�V4�YDqq���H�݃}]�@H|3�QЎ�j��a��x��|�~	�Z��P^���'k���8y
�s&���>����(�Wb/Y�CXG��g�؝��X�D��(֭IF��0P.�q�4�ii'��[ӻ���ۑE���"��/R	o�$.n�����ƕ���u���;@�W�Z�@l��[%f�k���	8���9����d�|5�
��5BH�jr��03R}g*[J
w��7+n����W����s���=HN�X��w%	��Q�L ᷣr_�f�����y��0�D����/g-q�s�����΢ �M��S���'��*A��z�D�f}�qo���;f}U7��� <s�)%�Vl"'[�A�f�Q�T���5d�%��'����~4�[/v}C��ko�5�o�:�퀢��6��ʎ�aҮ0g��O�F�`or �e�90.~qh|������w��m��B1+ ee8kL�WRKH��7����\!J�m]Mm "󠏊VO����k�ߨǁ���2�u�RcZ"{���B6u�X���w�=!a�h����zr0 ����I��J�'��sJ�����C�
����pR	z0I�yZ}��֒�j��}�7<�	a-�yk�gh�$������f�0���Lb�PJه�h��;���\/����4��EB���8J����������Bz������}�,~��D�p[B
#x䯸U_N�}7�π��}��c$�{�`��Wq|P>{t���&!U�*�Ѻ�h���x��д<�,v6{G:z���D&�ii�y^�S�L���l	��e���}1Ai[�J�Y�3����.]�3�uA��,y����At�h���m����-i�1���E�[�(g	4lEB��"N�eI��9m<6���3�%_�ߧ�.N�;^�4�ϝG�Ӈ���7�f�vҝ¤ǐ��Ml��7s`T��l:�=8�����H��r�W���`���吝�?ԆG]��+�~H&��^04�X���Wgq1���1�s�?����@�n)r:͌o�n>�{ޙ3�ӲPO=�È�S�T����y���0=T����Q��XL����9�\�~����Y1'�LɊ�nnO'���>	c�ǡ
i��Y7�""UƔQET�;/���ΌL�<���"O�1'���$��{���օp@��%�/����-x��#g��Ѝ?v�1B�8S� �`���e5�,�e���U�cl8"[b�����S�S�~k36�Z�'i�.^�<9�Yg���F��J��s�·��OE�><qbO�v*�=q,��8^������"�~
����J��������Yh��ABha�AX9*�T���D�G�.gA4�����}���oFH=S�l�]��\�h1� 5b*��?P��WDx���V�.�c(>�g� 2ٻ͉�>�0�ìy�[�m^���^g�t}kGO�\�]e�Ɏ3�@��K�����@i����#,��4��?�E����hT��"fH�ᤦ��?����%�r����Ek�,E����G�G�\ou.'m'��L�()!�A��� �4�|��?��@����jv�]�E|��1p��� �t/]5I�↎�-��7Ǆ	����;��M��^.�MFmU���dQT�l������5kΝaǿv���μ$�[(^C�/�ZJr/J���T�nu@st��ͅ��k����~������9���[����BYǵ����`�iC�"#u��^D����i���0I���4��N�6�%L
�D�+�ߍ����Ri�\y�²�9�*/	�݌������Ї��3���e孻������U�iլn Z�+є6�E�"�C%I�fks>�_Ʋ��e�:9���g���,K^�S�UX$?rޛ�Ѥ��@�����gjԻ* T��n�]zB��R�� ?J��r�Mre^o$�2*��Z%^L�:Q8�����ixY5<s0���oݗH\�[0������Nz*��Sۆ��OX��.����g��0�Zco�h�zc���~�7��5n��f<a��X��I	}N��� �D(�5��U����i-$2ލ�iU�"�"�[���*��d$��r��@�#�ͦr�zN�%�+�hB�a��f�i�@,F�8����k�x�7���b�}2l��L���Y&+=Vu���o�#�'E��Y�$�#C�1Ms�*qQ��$<	� �tQH��:��V�W�I&�@Ӂ��"��v����S�w�h��� ��]R6��;psZd懧fZ�r�I�X�o��%u�#����N���T�t�&U=����V(� ��� ��LhR4vﶓ��S�C%�2�1?"���P\F�	m��ShA-��$�g0��ƺd� �����4ƙG*`�f�u��l�@�ja2�ZV־�8���>=E�"�Jq�,l���0˔����č
p�CX�E��ǿj��1`�Vs�ll����PT���6qe�d	�O��Sm~�K2��S6K���
��'��F �M�[��'��<�6�8��r��?��3�jS��g��l��p|_�]��{�O��&yF&I�E�L�_L8P=D��5���>&d�b��%�_=o�� �
y�~! ��Ӵ��]賭����Dor�nk��.ʔZw��rNA�ߌ�,�26�6�D�(�鿮*�� �y>B�y���5�f4�����yN8q���(�mM�D"S�WH$��;I~��"۾����]7Mv��J�r|c!S��� B�ɗ��Y�C�3��-�d��}W��4:�?r����(!� �՞`1K��t��0��b�(� �컕����?hy��'�ȳ���P;-���qRr޾��O�-5�Z��<vGb��=f� �"�81\�_��h�z6�c\ �-�W@z���q�v�N��L6"�;	5� Ν�~;~�αSmސ��mގډP�8WC�,E$#�{���<C�F>��;�G@��K2C�����[�df����פmr�	y��>�Z����,��=�"<��+����T�q
P)��[2&9w�ʕR���6��(S�=�~.z�៬���O�����r\"#��ME�M�}������!{��\lR=��Ch#[�`��=C�dTp�ڂ���8~�5i�4@?�L
8�@4���ʓ҅G�x[�-)�4 ��t�������|�<4�5_3�.��9Axb��<�_˚��g��(�v�S`��p�C糎��>uR}m�	 Cc�w��j�S��mV����*��r�J��ĖRRSـ���f~_�*�a#�9z��@����f�Iʩ� ������Pm�co�CO?j<Y��p�����6L��0o���"���~.@��Y�sZ��t��Q;�I���j+�O������>���XSZ�Έ�?�Ȓ�?�)*V�0�=y�3余��wl�������V�1�Pdq��V����?�Ҽ�tbr��!+$�1_yC��ؖՋUp ���&�4�륅I*�.�ʰ��D}+���nz��)�ѤBG>�ΑR�0� �j�R8��.�v�Nr�&}=%�ٸ<睥\�juw@L���X��p�v� E��#H�<30J���W
��b���wԝ�0�ƏMcQ ��SF�z��4KM��S� AUQ4}�L����+�m5�&>�b� J��.����QnXF��"��F9�~#��,>c�1�F��5���b��UD&S�!w5^t�"����qe�XȽ��P{�=_��&����]�ޅ/�x_/���<S\Kq��o�:Y;�2���)�[���l[91�/��~n���������L�<X��%;�I�P����$�6���x�#o#�j}AJ��|��c�X�(��P ����n�s\IIV���>N�v<�߉���{�Ǜ�;��Z�1<=�NH�����(�X�ivՈ*{'��_�=��E�^ey���p1u *���ݛ#�Y�v���hL�$~EmP�n{VW��qnK���s��u��D8��>�~�vmy%�hf�5o<�����߼w%�;�XT�zn"��O��	�1����+9�_�k����^A3�~v��t5�$<����o�D)��� �qk�����y�������UL�b$
4f�k{"���@�dstڧ��}j��Y��.�#��R��͋K�;ď��0k�h$i��YZ3xܴh-�]�/H��Y�K:CK�x?n��Z���INE@�e��/���������!�"hB��^ڣ?N�VLXЃ��)��A4Z���r:���"�%��k�l}E��@]�� �x3ોB�{�hyQ�������mν:���Xg<'j��dd5'-�9W0�Y+�Rn�欈#��6��T����-mb����� 9nV,��|C�5k�L��	ߧi/�<�ѳD���G�%�H�|ӽ��y����6Vz�BVp�4;��+�YJn��H����N�9�s��򔔿���/��o �"�g�eU�l��-�(F�3�ʅ�t�j�j��IӃ����tٔ��Iz�������u�:����Ҏ��b��� ���
��K�<˜q�`�8�40R�b��y�,p�/�2�A�jc7f�f"c���,���3B����8���E��$���+��E�ح��^��D7o �9�Kf���i|�Ш��c�� ��&�o9�w~:3����-a��� �f�g�hz���VP?*��B����Q���o{���Eȕ$Z��E���� $݀C�#����!1���4�PW�p?�+:d�@��_'��Ϣ�ºѭ��[d���c�ga�%
I��Ry��4����T��>d�_���c�e�c�j<�
�u��t��u��������>Go�#������\)�xVcтVڰΊ=���蒀�xehc�/��@V�MM���*J���9�����+O��=6�	�	��`u�H��2B!4�e���;�j�r�&������n���`�f��t�{��� ˣ>�hߦ߱��*���p��q�s)�ò�+3-|G�+�l�l־��+���h��g����ƿ�~pjiț����������瘚�S�������\Wl�!/�7��cc�x|&��L˽V��و+��@Էx�G�J����"��t�ڽ��aXW��Q�[��B�j6�8�Ϯ�*��-���:���!��i��c�:��%�.0�Y�u� a�WB���f^����m`'t;�)fo{�5��B�&f��D�]�E�m�7�2�]w��Y�%�vU���1�p���%�@��
S�*\�9�m���N`���E�-Y�ei��\ß?���5&L�HS˓��㳃����eS������_���͋�bۣ̌�^S��<�{����b��r#yҳ'�>�N�ׇiU��2�R��~8Z��-�a��A�����˩��;m��=��v�+V�O����R�i�MG��1g�-�EB�o��/G��,yk_�+���`�GŔ$����@;6�t9s�y�� L�AE���Խ.Ru��@`�͍��Q��we_q�p�'�'=��ݼ��.���Cc'�Fp�	8�+�߳�0�&�L}�-g#O�ߗ>n5��IE�m�֥n�
LK�2��q5o�9�L}W7��S�xx�"�.gf!)�J�Ǥq(�ş��7v:D�#�3>��?l^�[�F�65����+)Y@��G�Z������bh�ғ[����L��(����3�Ֆ1A���*	k=����G��N9����fiL�f`�(W26�ǘ@�+�BP��k���y���?~|t҃'��]��g��<�?
�����^�SN�X��[��Y��[JV��<����\���ty��Pԗ� z�]3y�p6�?-�3�����F�A�mD4��m�+��.�ìHLB�mz�ȍe��ˢʫ+�����Y�����ٛ<�~f�b �`�K+ӡ-p�R����!���|`#��_X}+wC]�op��\B �^Z.���(jH
�8�@��Q�8�N���z�e�
ځ�K�Ʉ(�c_V�u�K:i1$�WSMK��w��1W�����}H��2�"<�BT
U���Rg��M�����w���g���ϴ#[�	�&I�X��`@�V8;}��%q]R^Ķ��۞�6���N�@9�k`r����90�O`k�e�ȮV����4�5�Kߋ���S���á� ��t}�(:�-��\��o�5z���ˉSྶ%�^�PYMt �\Ch���ռ;׵���?�:���Q<YX�֊�1gl0V�@�2���r�gB�&��m�%U����М��^��89[yU�0j�P��m���K�B�C�**}[����)��M�ez��7
�B'��sy���%6z�+����AU���w�~�B�� ����쁶��R�wr�A���n���Ǭ�4�/�;�����MA��ڪ�&m�Z�	Z�*i�$	
�}в#�sYM��R�v�/Y4�e䪯�>7��&��V(sU.��} m ��,�S��-DB�t�݇�]���� (De�?ȿ��v�w~N�4�����������ò�Ľ|�-@'���m¹�/$E>&O=�Hns/�)���M �D;�@~53��'�S������!�(�'�0�e�g�B ����D����d]ETa} ;U�ǽI�a�~C�i�f�z��`�=��`_	��ޠM"��h!��JT��$l��U|� 7�em�1�|�K�o��p=!mF��؀[嵣�K���I'w*�6-��$�����<��F��X\�Q�I���P\�(1�J���-rM;�57a��q![�5&�@mZ��:��y^&�����_��_�����uo~�W��D8y�k�4�g��jɃ:�ٺ����ـ}�'��S���#��g��7�SRI�}N�ܺ6�%E�჆�{�+E�bk٠�/�$��h<���'2����e���,��U�!m�_�{6��{`�;�{T��C;Dci�#OI�#��J��$N�+@�1Ay��P�?K-�Mᨈ�l~ ��]C�U�Npظm���m�A�Eمa�b}�lg����݉I�s$��EX�}��2���pM}A�7A���}�[���E+� ��9U{8+f& ����N�P��5_z�Az�7�	e���^�	�y����Y��0.�h����̌��|S�W�r'J����i���s���'����OnP�}k+;-���3J�ǜ�a�W����dk#'��!|1�;�s��̒�4�򺖌nAR� 9"՞愵Z�Q���Ś�F�ʯ+ ��HsNH�4[�?�7U�q�)���m�a�W�{���.k�FQ����5���=�N����HrOr��t�+/f���S��*���u��^9es������t��O	�זPr�U�Ͳ�;|�,�Z��q��G���pP�0��"�n	��u<�|�;tN�k�K�����Q��O�M��~.�W����/#�G�`�i��Ƃ�1�x�a��t�N�#�`[����j�!��9�g�Y�q+��&�4tg�M��=���pq�Ы�L����6���0�e���s�xhM��z#��A߃������ �z'��A#c�p1�@�g��ɤڭ|/.��0��(tJ�����$~K�):��z��G/�%n�����9�|8�ܼ2[����;%#š�yJ9���T���
��c���]������)#���z�-����4rm�)��?�Q��U_왖�.-��?����`��"yg`��@��ɟ�9����:ى:K����x/Ituq>�� 㧍M򠸌�e�|F}�T��G�MH�k{�?Ui�A�˸��;���қ$MN�����c\�Ai��'�~���c�Y���lD��[S�:��>B�t����W�$����#��Kպ��2��b�Z�?� ��6��N�-j�,�Ž �֎���p�͝KK��3��k���	��쥮IH'J�!����5��fC����k*
�a����'��o�U���,��׼��Z���yY��D�`"o��,����=|kH��*5���i�-=s�8�v�So�����y���+(U��������A�ͯ�iX���h�a��,BU^��:�I��.$�u��Vl>vU�2"VA_~�Zz���w&�o�I,�OE�lg�1`:�..5�eԣ���`�~�=T��\���ê�r�>/dJ���WE�.�6}�ݣ/���%��Bdq�^������Bxn�YO�m��Z���?mP�u�%�ٌ�A��<t݃�n�[ٷp�$���W��~7*��zzܮ����D��7�.��Q"���.pk����
����zwWjs�˲I�Qf����aTc2{�]�r�F�C�}�ҵ�Q�>cԅ�:T�t���珓��hu@RbF�����������j��c-�����C0	�+[Q���,q[~�-vH坝���w$Vs�ۥ�G`>��!�4��3�-0#���T:�l=HRǩ�Y��iK���d�{.��L��p��9.��γ�U�󵢔�ȑ��ӴQOSP�{��=ԯ؏X���cOF�
���\����9�L'�h*F^�����7���uj�=�H� �H9C��U�h٦����70�Dg�Ĺc���@O⨮qQ������N����*��J�g�Z��^���H�}�aWGR�~�����wo�L�d#I�k�s����J*S�0}A�����1<���L>�,�5��<��x��d����}�7'��2�V����;��aa�h���|\��X��r�b���lhVS���>��3��z� &ϳY��vlٮ!zO񇜉.\���#�4�����:�w7��"Ct
���5�b> ���?�
%&d��d%;��R�xl��"(vO�P!���Onu�]��cfa��[C��]�BB���������1I�;��i�$��D�&.ŝ�
�xre`%΢��]Rb�o��t�3�F@I{���t�� ��? ��-�2UO}D"x�O��JF��WS��UMY�Oo=���&��?!�V�y�07��(�+��ir���,�6Q� �՘d�v�́�4h�׽3�U�/�N{��+f�S������꿐��~����!ſ�0��n�;^7��%2�7 )5"٣{$��1{_����!7�ԻqK�a��x��3ޒ����~iU�)�ϰC������i*�������@�N��)�_[�LRnN��QC�@P�y;j̆���M�g�pU��a�Q�S	�|1ݷ���6���r�Rպ��7�k�d�fO�0�db?���1w�HQ�cK����P/�FIk�>/M
v粇gE3�j�h7�,F�Rd����l?��4`���{��{+S����&Mo+�e҃��u�O�_���=��W�	���"����M�����rN�q٦{�3� �r�Q�Q?)����؂�f����Uf��Y���*�!�[�J*h�j�[�$�����	�ɛ��A�1�����p����&g�DTS�s�jZ�c�8�C��Q��I�v��*w��W�-
��bR�h�e�
�X�#+C�K,�;7��J�|�������Q����+��"���Z�	�7S�|��$KD�ju"nn����:ɞ1�޴���3��?���g�  N�ї���a��d����Tާ�
id
�)�t~/��)���2n�mA����HB�9� �9�q�%��ְ7�f"�m��ɑ��p��ֺZ$���0/HC�%jR�?�&G���FV�(3*X�.��~�l:��E�\1~��Qˣ��̒&��nB5�6F�Ն��m�b��� 7������1k�t��[�w���(RD�X{�  �_0r�R�����L���	#��V�.ܝ��:��R���G�h!yE��^��)<�Kw˖�5���r`J��sB��8���4G���5���sK�`�j��ɠY�k�ol�{�8_ ���?>�V�=H=X{�l��zkfؾ���:���-�;�mj,�Xa%�	�!�,ZOK��%�=���֠�yzh�d�՝5�5��;��-���Z�S�T���u�"v(d�+��~4�ɒ������t����K�a��`�If�JI�;�,�D��@`d�^�,>�S;�=C��e��H�JKkUv�e��"|�/�u�Y��vcȚO��)?7��ɌhsMN�M^M�Q�����ȫ���X�����wP:%	��ԙ���<C�[;�f؇�U�]ܦ4[hm'O���
����wc	�ļI#�~�7S�^�i�C�5�R��X?b�!��q�e&��!�`v,l^�! 	񀀮�%����r
(�m��R�
9��Ne��ga��|�/9c�߅wnH=܁ם?ܩ���<��Hv��ߋ��<���WX��s�-��!� �l����>a^�j�oV.\��Y�hm�&p9���5� �V��w��#@��� 8�0)�� �jզ�t��=^Fp��`�6�dS��S%":�*'�g�rR!,x��5��&�,Q|�H��k��8G���Y�fK��@�H2xH	���{E������;��nI��܃��D�o%/�LU�E��xh|���mq���O�#B�/�_s]h����ި!\�h��'����`ւJ	�d;������4�:�c����25Ia�^-��xoO�qd�1u Ɓ���oɔ],� 죃�+�Ĥ�>QOz��C_���k�(a�����U�����(T|��������!R�_
�Y����aq����y���i��8���4��{Ki�^|��r�F�Q��d�33x�Zt�u�I�<��I$Sȇ4L`�Ӗ�7�H��Pe��pTCn��>g�9���'������r
�A���e��3��++����&�w��Ѕ(�t�o@�s��ݤvc�)�I+�Bcw�)\-6J�~&�s�t���;�%J���}������d\yS�+�af�59��c��^��	p o�E�*8|O9.�� ��*��OS+��a���L��7� ���W�@�n�]���G�Z�	B���[А�P� �7"C7��W�Kt���)_�{p��c��)���	s��R�'(n-I��!��� 6�����Ghإᶁ6�n��:CG_�L��|�pT���!��`�"����;��Ԋ��@�tѲ�=��,S�j���ZÎ!f�I�V��&g<�@��;-*�����'qș��;<~~k��u�'Qs��9��ء�������R�{M�"�Z�-QB��'�bJUQ�&z�_.`ʿjU�	�3@k�O\@~��Y3�Z5���%8�a.��K��8�c���L�5�i�{����8<8�������E�D�i�F�PcM��*;-�5(H�{V���%I/�}6���n�WJ���aj!�lYiA�,�Ā;����,��O�yn�T��k�`�4���&Y��@#�{L�*���|�d�����Ҩ@#ŁO#ˉv���E��%����6z��wFqξP��_�^g�V��Y��c$��D�;���~��I�m��!�&ܘ�Huf�LT}�O�t�))��-���|��]~G�|��3��B&�5�E\� �*&Sz^zfL�p��~��6�Z�&Kq	*��G�}�5Cp�!�{����Y����\P�b@e�0A#�u �׺�����R���&h`E�@O�!���l`�51D 3����9p�+]�y��*k���C�8A��C�GU�#�xA_?����w��9̵� (&������2�&O������	_��p$�k�kh��G0�23�+ ��TQ��sW���q=ܮj���n.Oz{	l��8�����
�'z#�3�n0�+�b���K�t�P�O%������O,Ug�N�\�_���%�kL<Gwb�2N����ݏ�=�܏�U;�hx��6,#��
o�w�k�%Q���(�G8��M�xq�8���+��
�ܯBº��`x%���������$b�P���AJ՛:�p��W��N��D��Z�}���o�mIr$�N�4%C��(�i<Wg�>U���d�w���e�W$e�ؕg,`DƭNy��"��{��+e����#.����}��-i,��G�K�e8�>�=m�V�Uڢ���
�j��]����-���]_"�h�z�i�����o�f��K�w��H{�l�^�8������&1��s�[ru�t�lXI�Df��[����j9�����v����M��߇/��h�ܭ���x���E"?ޗ�:]�VAS��`��v���H�K�2�B�TD�eז�����L6��h��7���d7��.@���F;ӎ�����P4���3�Zs�u��iJt)��J���G��DQ�T�р�N������8D�9��7�N�"�dز�/���� "d\��)��|*[A��7�&9�X��A<
/\�)W���V
����*n�:z4)�����z@�Ό����-��q���~
��$	�����&hr���`r�U�Y���/&��Z�e�0p�}h o`�<�EY�˗}����l�:������D U�e����I�u�au����h���2c�����Y�E��|��c�;��t�,�.v.�%ۧ9a�뱘�L�����fAD��cB<�D�'5�o�)˘�3�5c1@~�E��L�*���~�ECN��A�R��7'�Z�M2��%�j�7� 2����s;�.��:A�q��% ��B�󎠏+���W:S$yN�%Y顐��V��!`_�v*�V��jLn{�M=���8y�"�/"��q��= 9��'���s,���=�c`�9���g��*�^��D�����G�6KAai~�s�VyX}B��f?*~�Г�)xuy^�@ �Ь��&e�+�9/��>z�����2}��
sP�dI��g�"$�8\|H��˺L:O���+@�c���k�bŮߒ1�<�Mb��`����'�W�����Og�Gm��A�f�2�	��x��̬����J%��۱�͵Y��G����e�3ֲ�I�r<LqDU�e|�O�5BA#���d�e.���8��*)Z/\� t�s�jF�	���ۙ�!����"7�Ԯ��[�dBB`[A�N}��x���N�t�������Ֆ�Y'�ZN����;�޾J�����L�T݈�c+���p|�_�L���@D�8C�u�S9M(�*�H�K��%e�[�ͳd���J#��6������-�mPUfZaB�r�ȵ�q�5.|�6�Py��w��L��?�_-��`؏`�#'��+��>я���J=�U�3��?:���ۇH��S�K�ņS� aU�|l��Ѻg̻=&�y���yH���a�%Jp��Ğ�يA54�]�_Kh�� : 5�U��_�V�6h�d�&���֓|�4������@���*��<v�^X-ʬi�
��z��
��޷��9�sj��9�,������Yl��#a,]S:Qؼ���¤k����c�<��5r$�x�0E�Mؓ�*�q�̽~@d�M'�c���==eG_uP��n��
�N�����w���T�W	����b�=햐O�wR������C���f(����L�7�x� ���d�Ï�ywk��Z(�꽇���d�5Jb��:�O�nu|��<s��Y��dph[v�N�&�RL��@�5�+�:� L5�e�[�����ɓ��8{����lyJx� ���s�w��c�*�A�:i��w�'��6�Z�o����q>nO�~]�o�?ôh�Y>Ĵ9J����Tbb_s��� ^1ϑH�%�ǼF洲h<�i���Q���pڕ��*�Hz)� !����?�8�-�����6��r#����7������m������ZG"��I���[�������	�p��>< �p��ȸ6���
B��΅|��K�`���ѣuX*T�e�qZ_鲥�X|�`X�.8c%���^�,�7�/�[&��Ƴ
>���9�yT7�r��?Q�*�7R+Z�>��}2v�4(�)ͭ˙�$����L>�=W�W=<��w�a�k��_�[�h�5�tZ�-C��rtZ��j�u^�Y �!G�g,<CI��&�d�}�¦�I�k-�Ӊ�4����`_+y/����܏�~�4����
|`�/�X>a��e��:[��A"��+��sL&�;�&�*���c�F~�b�]�u��ި�fk�Q�j�ioh*7"��u{�����tq}� J�j9-	�w0�"j���*+�?7O���GLg�4�/���K�~�CG*�P겼B莕C�U>�ʨS�R���6����39�jK�*�J�P�Ӂ��x,��ʂ2���fqTW�Xc��S�;@�����;�9!�����L��%��A�,�X�oBaW�g�Rn���&Cb9�9$�s��ֻ�fe'��+!H`���aH�N����6����Rˮ_P��3��>�6V#�F����/�������,�KU���y��I�=%4��S{�ڂNc��ʷ��8�fѸ�\��#�5��	���笐�)��Г��^�b[�K�}���B�I��S��s?A�0�J���o�
��Q��O�H���u��#|�#�Kz��B��߹�.J���34db�k��S1{GƝ嫹�Q"���T�@�-?3
����K�����	���W
[H�x5�X+╁(���Cw�}5�} r����b)�sd�"k��'%!L��#�n�/�3\k����Jh��n�x�r��>�U*�w�B��p!Q��\mzWh�%K�`kr��D.J�<qh��zJ#"V��H�:�W�_�Q��8��7�fA`��rbrv�Җ�l�`9�3d3��FR�^ �8��<���r��b�x�E�������h�:�0%��᪏6��d}��E��a^w�R1�}{��#  ��L�楂�X��`���jf|$Tu����ݮ�f�"&�ӡ뀾T�'H��_aӻ�A�1������޳AÝ]2���Ps�H5�Ҫ=Jg��Q�﯎$��aaHx����n�q�ђ���C�.Jͅ���A�|����Kc�W�,��4А���4tI��V;q�3O���?VQ`"�	����D�t���w�'�0�_�@��BH�����
�iV�N�i�=�jr��&G�?B����'@�%�O45|�5,�������u���1v��W�����r���yq{�:��xwDR��C���Mp4D����xzZ��)�CSG&�J����^����K�C?' ����3y"x4j4|�}{X�������w�|��֦NAS���E�<��ԼE�X��+�?C�a��ir2�K�U�!j�Zw��Q7b�ʽ
Z��Aξx
�����8 |��6�阃����S�d�* ��%��˳�e��j�+_�톟�'�;���Fm*��L6<��/���
$A�7Ym�Mh���m[�4ss9�6��fX�Bi$�
��ep��C����adf���Rm�����7ͷ���!�"&��-[c,sdˡ�׋����s��S�ױ����٤������]{~�3UCWKi?|Vc��4A(��f%EmdOl%��>IK��]���H/�vlRH4;��x; ��PJ�0i�X� ���, �?�	x3�9/l{eD&���0u����?�R�t�U��]�Xi�[=Gy�lTd]BHd��djP\@T����+J���TɸHa�oZ��s��U���7�8����
[�ks���N�!�CcC���8��A�o�3���g�S?��u� ��tb�>�"�{�N�r�Z���yki���D��&�DC��<���ܝO��U-�s\��f��`���	&P}��M���&V�*����� Ɏb�([�G�.X+��
���/���=da�,*��8Ia�f��E*Ճ�r"Ě���:���':���G�ֵ��b��x;+~Y�tF'Wp���K���/c0���+U�$�V�Or��}��w9lل�O�o�\>|x}��n!���EC%Z�Nw�U�G\&9�}8��8L��"��H~W�q��$�އ`��l/?���`\(�1�#�:ѭC|�=OX��n���Xˬ�:�\������� �p���m���((��=�ի��_�=�5)B��T��T���x8��v�t�p����T�9;d�"*_[!M��>�� LM^�&��	�!X*�;�S������φ{���\��-]�F1?~�岋6�.�a4*�6a~(�W633
�c�V��۬"C*`�bu�Ս����P��@�H����"]�O�Ь�C��m!�9y���X�ʸ���WH(��2�3%����x.�����Z�z�cP��!�6�~�p!Հ����g���.�G��[,�Yv�wP���<��~��]ZAL�?���D�DP9H^7�:=/EF�[JF��]Q34c���+W�VSQ��ɷMgd󝎽m��x�g!�4dQ4�+�Xև˞}4��?h[�o�?0h��%7�y@�Ar�17�(�͋��4'i�V-�y?<�35������$�P��~ɒE4�O�~�v����o�
�#�c���T�3o���C��	�)�Ꮽ��?������$I�#��ز��d�r��l������OK��t���1?��<R�aO���Y�du��r�<��j�wQ����nCy��z��|�L�ڦ$ZgՑB�+��;��a�Ǿ��"�Q���R��Xp�Bu�5�&yl�qC&��շ�H�N�q�܋㑼����U���Ħ���}�j�w:�aNg�Q�lO�ZY�!q�+�4 �P��x�5��e�oQJ���s���0,�5D��J�� e����U�K�C`�\���1ze���(.c��]ڈJD��m��I?�JT�J�;�Ɋ�9��I���6l�&֜�t�&G�j��j�s�?�mE���悎������.�,�Ѡ;�E�X4i���6�#�ƧƕW]��RJx�����Z���,�`S~Ċ>��
�M)l ��Yh$Lp�&�S����;�����iVd@��㼨�y�<3���zpM��	KQ��R��^�u���VI��AiA��Ub~
� ~?=@Z�%zP�By#]��/e\7S������-�J��ZT#+�˒([�hv�p�?�U��B�>��<fI<#V(	:;+�dX����y�,��];C+�ߴ4����,��l��9�J��A횞1Ƃ��x�$l�FO]m%l��c���~ܸ��ې�XJ�H��*R~��p�k�����5H������s�0�s��=$��ۃW��Z�1�~�[F��t�]��"텑D��z2s�݊�+�[@y�6Gϰ�è����NwsF02΂�Ďb��L�21���F�j�r9��%$ ��e��-G�l^Ste��i1t���X�������h ����<N�c��H
�r;'ĵ#;��E�j���M _�{Z�IE6!˽D-P%�����@"xf�d�v:��]�`�.�E� � ���9E��a��a����mKL��"iXa&�����3I�a����V�z3��k�l�Jl�y���8]
E�F��	ο�4�A-�T�GY�:򂠃̅y~Gy��k�M���]T�"ͣ�:U}�y�LY
�tuS�
p�	|���j�Am[���mRuYPBG_�7�|sO��f���7���N*"��r��n j�Qb�����^͎˘"I��q���j�P%����[_EK�z�F�4h��G^Dy�l�͜c���~RT��wg (��u>�y�w�QM�O���}�R���nHE�o2;�5���ȗ�h����?yDפ_�{�,*��N��}�B��
l��FY�X��m���%*��̆�IgU8B2 ��&���a��o K�Q�5g��<�	QU���W81�s��#��DSr����}�D����!�+���'XUߧ�K�'�n^�Ă�6�G����#�)�e��b|�C/MS �z�m5��}\����<v��qg�]�EkF���K�'X�܀ ��k���k.����`�G\��5���Uv�GQ��x�ӞK �<$���J�oI1�QC�D("��쥂E 	�j�L�>x��;;�@)��J��x��I0��+�͌T� ��R��7�N��s���9��qu��?/V=�hPƻu?X��C��ן�)�B0փ#%q�������h��m��^X3	b��Ѝ��L�nT�1����a�@>��оN�S����9�ޔ'ӽG�H���.�>+>�hY%�1#c]W�}.0�����zt.�z���^��;��X��h͍��3>-������J�e��4#��7>T�(��@�9v �)A�B�!O��Sj��7ޯ��L/j�;�*�*Ve���t��y�I�dh 1lczb��B�A�k���^߁j���k՗�)������W��!ҫI�P�u�f��$wP��j���-@5�1��������Ii(�l�s�D9م��-�Q���J6�.�?̪R��;� Ƶ2Tb�fՎ�B�s�^Gg�vN��د��xEb{m�=�Ӽ����uc�\��� ����+R�ݪ�źVxҹ���P�OHy�"���r�879Ug	]�����6��@p��K�5ɘc�ϸ/0�t$���+�r,�ˑ�n���p��ַs���y��]�b�h	Pmp�J�������GK�2�U��$��	�܇�����@lt&��t4�}�Y��׏L�bzb��0zrg��C��5eR� �������/��^f���]�[�5�3��Kl0$�C1��k��W��l���2��@���]�J�d�%Kد���<�Tc?w�C�Ct��>��y�i�ۊ3(|(rW�.ʁ9I�5v�%�$��bϐ�SY��`���2I�$����,Kr�K��@�Z�X�W�����ˈI���\�Z�	��[`�Ip�D�LJb�u�PY��p�/˲^���ŔjD��F8"��I�Ch��)���V9�g��8�������O�^�-��ÁY]�h �܌���? _fê�M;N:U���tZe3�,�+h��8iO>I�T��U 	���@"N� f��r_���g��[�f�k��)hdէ�R?Ĵ(�Li��8��C�w5����}^1Q3��}�����藂U���X���p��B��k%G�p�e$�~�$hf��ݧ��M���[������>���')�~S�e%��9R5-8˧]��ܖr�mUoֲ��jۯ���~L=�M(H��c8q�8�n9�ϛ��!�>�(i.T����n&Y����W�^[�H0dV�Hg��z���#�6Y����.��;��#� ��fgw�وK*�����IV��T�N#p�^Cj���MC�n���~�dp��o14�����\u��X��~����uנ:6�|��	 c����9Kݾ ���f��"'�a��)YQrD�΁t��j�+�l�u@b�8����n߉��`�nO2@�LnHU�����M���(�1���\�j�,�Z��6kv~3aD�L ���=��i�/O�w�E��W������]����t���DGA����<u͟�Ӄ6,�����;v�A����No9#���c�>7/$7�/k@�	=B�I�.�F ߔ#�)�Khȹ ��>����%X0����T{�*��B���u�j���>2�z������{ ��*�գ~Wy����%�W_�"�����������\�߁�����5���Y���o�ke<�A�
BY7������g�S�P�էW��pX~���E�_�o��ᮊ����)�5�sD(<*��<I]��Rwڲ�կ�ܾ�1]�{�Ӈj���zU�@8�q`�ZM:�����@ő�|��Se�]�V�
@ފ��C�X+C�^V���R��Q��O?��[�v~OT�$w饏�#�H�RtI9����{v�Vy4j�J�c��=��`����,ˬ�h���Q�lC�~ �Hc��S)vL��`IS��3��Q[~R`�ܹ*�*�d��;�Udhq�?U3��i��J*<��6ޏ�lf,�/��_�� �-��⏷kP(�bp�(!Iދ!��+��eH��������a,ȳ6��T���@���788��{�ƥXo�X��7���Vl���Ep�3�91JԸ�h���D���m�(''˗^V6m���w�+�_�\-�/$g���Y���9��LT�a$�|�A,�i]�q]�I�)�����%N=I�
�gޣA��Y!j[�qu�(���>'t���I�|L0U������O�<�4i%���j>�3pdV�2���	Y�W�qnО�ܺ,[n��w��	�P�U��<b p<�0�@�����X�o�wo����_^�u�Iԥ�`T�n�	������\!U0�h��j���Yf#�0I�8EY>��ϧ�|C;����Q�F	�b^7�f��Բ[�{���p�9Œnt)w8y��?UFh�f
�Ke[�"�{������X��,=~�8H}�ECϗ&���F&�?x��v 6��X���-w�B���a�� <2o�ib���62dR����6Զ�"ϖ7��?�OmY����D����l&d��ð�ڻ�-�"�j�NNT1k�m0v�l�ڈ�^�|a>�
�̪x���@��ҵ�e��^��ǚ��fr�|�ϰ͔L�-�5������{�X1Fz6.7�\�.,_�����o��Yާ �տhr2m0E��mֱ�/$��/\pb�O������ҝb4�������?����$�GW΁���C ��,n׊E@f�NFg��;��Lq�J�OJ�'�A����b�
$� .�`',+kXᔉ��%3�����,��k[�X���f�2.��6A�>|a�-.�`��[�dN�f��Z��NV�H��E�Fyo,(rc�,	��W������#|h��w���	�ӛiZ氳��/�_�Ƃ�dٶ���'� )>e�i��z�7�.����I������s`�	Q�+۔%:Л�\Y�$�|�䛮�e�U#d�m6E�B���{�W~j�U���|���}]�q��E�x%�_�����yM�Y4tyw9��_��X9an=RNu��h�	!$� }���=�������b?���/�	U�������� ���N�"�+ 8�>ՈP㋄^�yxB�f(���b�즾�yB�!�������f,��k�L45���������k�m����ĮI�7��}/h!�D��ZR���#�<� �ZkMԘ"�)!�qL^g���F��`� pl�<�3���vK�O~�ϗ�O�1 ��&)�I/���1(��'#s����r��{��U��΀8=jM�!.k��
��Q1J:��	�nG nk��צ�F�}@���L`���F5Lc��_��1u,o[8hs,�f}��x��������8�J�ݯd \<&��U�6A�۪�t����ۻmn+C���oG��Z�no͉W�/���n�.�>ЅOe�p��Mv0�i�|u�v�]����}��A�i��M�:2�xJ�����}�-�������_�������d�p�=�<�Xkr�+�-T�Z��4u{�)#?���!I�87�~�����fI`;K��XL,P�B�݆��FAo��X�}[�g�����k`�$'��g/Z���v6�/߷p�)�NU���p�g���(L�e�z*���)"�؎����sѹS����σ/�3�=	w�)���w��d*>6�(rO���"��>���eV�m`�0� �G����%�(�<�>��@�4� .����@e��'�n������ָ9qJ����\Q�'��s�彼�Z�&�j�c��"b�.,L���1�K�=�G4��;I���&#� V�}NF_�r)�x!���r~�*�Ȑ�Hh�jŰ��B��V�	+�B�W+
�`�)�+�[m!f�5׭b$�$�n&���S�����\�[�@��=��ۜ�#	�+�!��@H����
3C�d�<�T���p����r�ʬ�T�Sk�q�����-�n�jbn�h|��&�͏�J{fxPc���9���Ҹ��X��FN�k��\Q1��!pN��t��~�q#ov�.\`��� ֣<���� ��g'�z�j}��l�LP͐�q-�=?0�$�F��?_��։;6�\��~Y�ZZ��Q�t��J���w)�N��7+�(~O?�*�h񇰐�{8{�!W�]�2�[D�P _�F+�LB�xU����	7J�_��`�����0�h+Qߗ������n��\��*�:αK���P=B�s��[�������-M����[��x�r�3 � ��a|BȽ�)��Z���~}6��0�
���&���ڌ���Y+i�5w���Gۇ�$K^

��P�~�1mv�pF�k$�z �$�V��qL���*���-f;4����jZ��U��Ck���\��L!j��P9�C���=�.�H2D��;ӵ\�?�P��#��s���1�.��/g�OO,6�����1��j�+�T��7���"i�m`�9�oĂh3�zEK���c˗��?XO$��}��� o�͢���Gj���枬{�I]�6&�L�S�^�Z�a�7`Z~��S��T�Z�ۯnƳz<?��8��S�� ��5���l8��4-B�7��Xuk�w�:dTs��?�?mZ
Lcs���w�x4�f5�)J���S%�	��?#�����ᕺ3���ʘnl�U�*����s�Ќ$/j�0�s�D0��+���8������;��/��{�,)m㹓��ց��}å��(]O�\�DU�ۺײ���PBH���7��O��_LelQ�6��
�l�s�Ĳ�a<Mr�6�Ǽ����k��6o����J� f$�I�e��q-b`I�y?�Gr}-J�Kk��iN�m>^߹���ǑK����ł\)P�\�3�+�@��k�OqM�4�rH3R��1=��i�x쀜(���3�1o	'��_�=�S�c+���7̺ƾ3g�ӝ������Jp ��=���X���P¯N��9 7����p��[P��>�ϚYl��o9V�!Y�ZҢG`�ܔ������6R��|����A�Z�!���٘�����<ea�� ��s��F�?3��vT>e�z�r��\?��o��^8�WT���UЫۊ��YV;�	�@��|B��΢��`*-#�Ko����:ᄾT����ϔ.���G��z��P�*2����ö��>���١>�/Kjp������iQ����P˿��_�p�A@����56��b����ktg�ۙ&g��Cn/M���\�Y,�{U�aB1|e���O��=��Qm�[�CZ���4z��!�OI7'R�YAj���)�<c���sb�g��vZ��Nzz5��9��⸲���M�SI-���l8*�${O��t�W/�-(��]��#3�f�B0dc���[&��|��j���/)�&?J�G��E_
�oc�r�7K�G���8*<;�D̔-��j�(�e���OWjXZ"�C�kю�$#��d�������YHC�RF�h�K�	AAIE�7t���������5��e�6�{�B(�N!�c�b溈$�LD���� �
8��Z&�f���}��
��_�[
�|-(�N��]l�ֲ���6��!�o�=h���n7�~]v|=��o$�?<�˥Ykܺ�hm+j��(�!����U飈��l�="/�ҭ�X�A��ad�m������ុt��)\��JE�V.u��a��� �S�rk��q&B�ժ��:@	��[��a��Wu�3��?���%�}��?��H��z{+=�,���ۙ��A���o[�)RP�UXy���#_6��}��~4Q�\��nz3H7��Q�c��`U�(Ǆ��#�����h�|�h��8�WC(�4��8����}�DӠl�Oa����f��g��pm<#`��d�[�_h����b�*o�Z+���;+U�S��gǐY�}��CM��V��Y!�E0�9x�ϲ�|Iʻx����z�K1�Tx٥(\�L��h�=�ڼ�@o������K�?Rr�%�jLLq��ocS
K����ƌ�N��h�I��l�k.#�m��waa6/�H&���=����I��G�x�>��9O�4��8��M����_`ҋ/#Hd\��F�?+{����S��=}С��l�t 	��p����r�`������'r��xe|Paja�3EeHv�jQ�(�t(� S�^Q$]x..e����b�8��ƌFhs�2*�)c��C��u�1[q���(��f�*�5�fm�Sc���R(w�	>yd=�1#���j!�� ͥ�;A����؋&�̩w�
*�0+�C�G�@�U<�� 9���8
��^�_,�gN�@�L>�f쎇������J	v����c��]��ͺ��V2��Hj��$��=��`tL:jZ�P�Zgr�nF���.��S�|�]p�v�up!&*���s�s+�ȀIi�/��x��<>6�17Z��OP��/~d����[��6��L<q]��6��+�k�5��W��8�S�j��X�0����OZ�E}�رoÜy�T�Z�N�;����M=�Hc����C�h	�C���aI���4�=�:f�PZvxN:(<¿������*
�F�;�na=���$4�G~I�����ɶ�FU�Nq��q�Ө�
��/�mѤ;4�J���I	,&����彐	0�>|�����i�ã��˹@l��R��|���b.���Tޝ��`��V]�1�+BԍO9��F��wʄ��-���V�U2��7x� ���ՅS�-���n�M֟�ip�=�r�HA�z?�8V�ny���[.4�E�(Ua�ɴ:�J#9\0��O)��y~ �rH��������HV1w��1)��s��bRt/:��JN@��;v\� *�ǈ��L�ܬ-�b$C�Wq�ʷ+
��� �_,��	��!P�\)�K��;r"���}�r��L�F�5
�j���.0��_
!!�P�O)8���ddT#K����J{�K2����A�cG�LT�{�PY1��s4C�K��18G�7QK�����Ę��¾�.1�bD���p�蜂���1�
p��/Q�N�z4P��?Q~.x�צ��R-p�;���lF���t�=/
���B�]�۞%�k���D��?0��x�����l���F�UhNi2l�'�X�^�f*Zر��D�;o\�0��T���86�aE�7��`��M���:%'v��o_���n��u���S�I��r�V|>�T����nd7RQy�
����/	�d �J%%4o{Qk���g�������1،���ö�w˱�Ş�0F0�<(��2齍�?(.��@q�tP�aY~ \�8���AI�!���a�8�+�wׂ8%�f7�9�x��̩d�'����e�$������ѥQ�PG��LT<���ӌ=+6�'�3b�d��}��@3��f9�J�F����h�K+(�'Eν�7T�8�/!���������@��� 9�u`��c�(X!:#����3��D����*�v��ׅ���2�e�V�!B�/�f�I��o��
O	T��z��|�4qO��-�oe�>���s��h����o(0*J�֎��p�D���hM~3k��trfG'��@N-T�SW샸�)�k �o�
���H�Z�$�S<s-_g��L�1Rk? nz�@��L���?�ڰ��C7]m�V���7ǯ+�[��'`�}�F�%�나�
5U��Z����`�%qr��`�ܹ��
9$�i� /3S�L��nmXn�BE��UDO���0���ߊ��.�P�%�6*�H�����+�����6�1?\��~��-��ձg�������ٓ�,a*y�����o��N��/qد"ʓm�[(ϲEz-L��M};�I�}ޡ�T������,̛���B�o�PP[�O��ٻ*��\�s5����ф�~�����`�m���P)|S>�� �/8�E�E-�LCӉ-��
�8|�^�o�����0"G��lY�L�A5J����s� �i+�C��	5T��&rJ2 ��-?H��̓d����hiu1���Cj?:��u�x���[��|[r��������?��b.~m�Ǔj�o��Xw_чc
:�i$"��Sc�I�.��@��		M���a�(.���Y[�}��~��L6�g��$�V̹�tN���V�Ofk��-bBs���[��ԑp�����
����<��v$��.���W*r(��_����Օ�#Y �8��u���j?�ٸ_qrן�D-�޺�UԱ��/7C�öJ��)R ��P�~^<��3`�󕃠8�7�S9&d5�ה`$ۭ�n�ߴZ�w29�8�u��%��؜kK<���*+��U�R���(�kځu�'!f�	���_��Ap�y��ʧ ��FO���M�O��\��*`WLi����T�'j��Wƽ�U]}:Q��i��+����ԁ�]�/G���ʐ�O+�¯!�ק�P\:s@6�ĻIs���u)��Y�Ap�Bґ�c'~߾��͹��y
�(�@iX.ox�M�N��"�u�O| ���Wi�d;<�;���h��+�/��X&��x�ʁ���@ �_�t�BՉ^F�L�n��DY,y������y�*�@��(��T�u�1vl�}�\�)R�b	�U7�}n�'$b��q^�2	�q���S�j��s�K���8T���H@/���ˠh�P���sU�~U��{�3���K�}7/����:/�Lq
C=r&X��������z�v�ߜ�rz�QX��d⤯7�>e�M<�7~���Ki��l/���t�J`#�eC]*���4�K���ph�Z5�{�/�p:��!�r�bF�5���C��!�u��_���Ux�F9!,Nʱ�&K�`�1h����y�3\��a��#�az� �o]#�I���	���S��(t��]�a�������ÖV?��F���<����:J:#�nr[Xt�}���~�RN�g�z�M"��%Q�M���²ZG���i؀�[����i����m�3/��4_��� �y��632Y皷���Ѓ���2�v�-Q� ���5��N�~�.��6�]����3AƠ7Eop>��6L����Lۆ~KV�i�HlS2��P�
Kz 3<[���4�4��ZJiy�:В�����F���,^�@����Km1��oo����Ћ�>y[j�[�fM,��YP����S�s��K?��&5ep:c>�Њ��<0S�Ĉ鲮��E�����*�y@��5	����/�1�h4����~p��S�5��ԗ��GE��s�H0����vzy�����gh~c����CPj���;g�%��hi{t��--c�Oy~�2K����3Yg�IR{���6�[@�D��S݇�/����q����&���M���Sa�s4}%T�Km��.�]d��,A�⸥p��i]�=��V�XRc2��_5;��,��`'�q�=�TbkX�y�D�K��JO3du���~���{�6��x��%~��ȶ=1�ᶬ]��X{�L\�	�gw�(�Y�9SY(<�� pj�s�O!&r�н�(}<�w��64�����C�eY+� �d�_5WC�0�p^8���w�	����#t'��n����͠��,��;=����U���d�(L~��"l� N��+c�"~z�J~���g1�gāV/�6b:V�i��I�r����?Gȧfǅ�����gZ���P�"/*ٗ��P�z?��(���J\HMf��(�-ɒր*��6�cb��3_�<(�s�\�Ѱ.΢Z�dI&�MU"�iԱ�g�%���=����'�W��PT�Ǒ�L�sJ�W֦Dmk$\A�a�s�1�8�E� 6��E��ݪ�k'�qC��Ć�a�)�&����I�����䂇�+hP;�W�սz��X.��nNĿ��elZ��s���<���JQ ��N_�����c��%��8����� I
�����_��:k$�F�Y������Ǥ���Z�dD_vӕ���*9~��ZX
k_`o���d	��c�֣��Dv���Fo��sX ��$���s�&�z5���cO�V%�N�ч���C으@fV�[�MV	�s��>cQ��:�vV������#��Z��t	�[0������]��H��Y��h⸹�:	�8�\a��a���}W�O�6b�N��e�:'�	���3�Q:�^�7�t$�Z�[�]������Rb����{��:�4��>���;Lg\��!��{��4��Fn9���ɳ)fh��s��˂UlK�dƚ��~�+7p�/K�Ծ3���".�����·^�qկe��;g�YG��O��03��Piy��V��3L:j�'Ɖ>���2��$���h�֌Jb��M"b^�M#����~>��oF�j0#��*7��;}�vMG�[DM(���,��Xn��a�?~CD�X�-���$3��(�������nW�]+�{T6觵�ZEK��R4�јƶ�.�֏6�g�L��5�nz�k0ۑ\͕w����y��M��͹r3�pb���"�=A2F_Q�5�o
?ԭC�u��|���U�*�v�2x���@>5�< $)�!n����ַ�����`��`F�G8�!:�_�	/��r��9;[>ɑ	ar?�b���;*�g�e�R���4��)��^yj��X��D(AOKx��w{U"�R���by�<sͫ<�q��ө}ƛ4w����B0�C�V���4u�/���U�k�N�n`y�c	�]q��#)�����nO��ب�V�VY)���K�n�D��g�٦{`Q�dX�!��=S*�m3>:�
�&�'���r��QQW7��/�8��,��aĖ:�d�DZ.4��0�d�^�*���1�v����2��E$���Ϗ�-��y�5흝���C���)Q��N����'یK6{�{�� \�pb?���"@�2��t�bRA���� ��� y��8^w���?o5_���"�IE!���-I�o2�A�y��K�q�����k�XM w�-GR�XU�j��|�*7�#���0B���*�Nڋ46��r�l8AU��f����O!-{��Wv��}>y��^��4C�Sd{O63L�lU����[��X$9�x�*��%�[��	H����O�x���A����Vu�-Y���Gh�颱s����6F�
��J���t�Yq�V>R����{ˌ&��N'�k�ׯ��~�2ub�s6��X@��t��Ka��E������[n�79�>6��M'��K�B{ؿ��5���YNq�л�"�Գ�T}q�;&��%�gq�����G�YD��"}�巩��.uD)Mf������Ê��)�AGu>��}`9�H��>�t��oa�֘�-�b�(�!�mp�P�KK��g�OC���|�l��[�s|آ�ݑ~��1�^�Mm���J�x�8ݵm^������]t?��Zg�
���g$gRJ0R��2o�Q�	��?�2�t��;���^u�����Ƶ�H7ҥ�eK��8%�y��*;X�yҐ����7����9?���Ί��B�J��֥����6y�T�3�iߒ]�eK�,+б��~Dl�#I��8��U
zR�_ӆ�^�/���ܕ�<<��5�(5aF����R��
�{�N���/��ʡ���<A4��Xʜ� �	��	W&wy#��}��kkѡh#�^�&�d�2�e��ր��T�Rx�������L����q����%ʛU�p?���X,���?��O'�!�q��!�c���ڲ;c��\rx��5NѺS��͜B��5A��p���L~���x�80��{�s&J,/�M�Z;���+L�����?OQ������FQ����/�Oiz��+�ȧ�����G�.�n��u�������^8��L�m�_ڵi0�;T� zP�kI��R��>ܛ��M<#8�4%�Ō D��;��B�h+�a�mL*>k8�a�U)�V�Z�̈́%">ֳ6���7�}�m�p6�e_Y\�c��b��֦������zu�<8m��,���$�m�+G�.���	���[R����)M�����s0�����@%qp�5E4&l����)�Nn'mUW]D��S7hHP���ƃr�Ki�~_������ �ҽj�T����(�7�uugL�Ծ�f���@s��) #Ғ���b�4�;��<�2s�AEp�T$}�Lw��*�*���א6^�����+�1
��)��59[�oR��*f@��[L��<VB��:G�{!�A�:���ʬ�.<�L�o <?��ˎߑr�ۚ��/���M$�)Fd�f�1�'���y����u�f���Ʃ��A]�+���tNk26�<���G~s���⻘��7#Y��3��7��f�̪,:0�ՊD��[O1��~�Mrn���?Dzҥ��pvW���*S��W��1���㤰�.�͆�Ż> Ӭ-L"��s��)	�f�P2����B���P��50��!+���9�`�I����0o�l_�)F��l_]���+ȉ��6f��s�L���o��t+j�ր)�񺱮:�l��?�frH)¿���9;(��Ƌ����o�����ݥ#�|F�\�1։���V�4��*G
� ��,�Ŵ=` jH�� w�G����Y��؞�0���A����}��(���]�(ߌCn懱��i�lէ�؄��s�n1�Ca*�
R[x�Z5c�7�#*;f����9�ܟbݪSI�c��SYm8b ��4� Q ��r`mh�9��`��z��n�l�Ŧ�� ����[�B�~ !���S� �w K�D�oq
s��A�T۔������w�f_M/�=Ŷw��e:S:9��y�!¶�����Ld�bs5�N�~_)�����m��|���}5�S�b��V���Ź9�M��z�s�J������ԫ�C���.e�SUY�XM|�M�X�	y�e��$�>=���mn%���|��Sk�;�`�z-6���\�g�"������~l��ԕ�]��7`M�qEE�;]9Y�)VVD����sE�����AP�N*��-ɭ�i+��%����{�$��DFQ*��I��!=4&�GU1p�b1T}�C?N�ޮ#���
�RI͢�T��dφ\�_��iO�QWTc���O}9��bh�_��Q�٪G�??rY�Dş䔲,SpYj\S����Sc#��k���(vJW�S�.��C�Z�G\��@��㕼ƍƂn�>��hr��Ѥ:-�����p����F��L~%=+�mD��|�`^�>��wb�%K�)��'��3u��(����bW2#d���S%��e�6���"�v�$�L���\��޻��M�D󕜾ol_�E��Y^�ky���*����W�8w;����K��GK��j�T�),��x�:� z�g���^!��?����tU�M��M�/+��p�Q9�X�=�6�������p z��x����%�B;v�2 �T�=�0+�c>Xu����G���A�hgöCnv��Rf�ZttG27M]�@m�C��A��f�!��D@�Tnm���Z�5�X�uBcMN�K�0�-�8�:U���ɬ���"��|�\�آj��wK�6~�H)5��?5Q�W>p���R�A=���^/=a7�z�z��E��J_N?�6��X-Cb<ks�ҦNƢ>�C"�9�
7�fT�Od�R?	�n��%R�Cǽ�G�.��f�|t~����\KOބ��Vꮩz��[��"�v
���gB�/�n3C&��OZ.O�G��@����*�c����g�ᾇ��#�?�}�~�y2����@�}�1c��������!-j���� 뤊G3?���R��9���I.;�EA�k���4Of_�.�9X��a��9��NU=��`.s,�e���K���r}�ҥ�b��_��<��@��x�(� n�@�.7���#��@�3�́c+�!��*K��Px�P�ڿ�{��js����ľt�ң� �8��� ;����J��8�F�����E~(k���Q֦��ݮa�2��>~�k!���cp�G�7(��w'�;f�b��S���v��r8&RLS�u�+�J�y4��U�6w�)af�E���ݑ���{Z���Ų� ���d�����<�B1���p��*J�}��C��@��A��G1
��c���i/=�u�֚����JG~�)�����X�.�zL`Skr��P���8.q� ^�#�zI�K�#���?ʟ�=��ҷr
���+5%B�	r�C�~"ިu8����Ih#d5�� ����,�����Q�C�5��A���L����ha	dY�&ѳj(_��UY�+b?G�*6��pq���$�<�����ks���8��!é�f�[m��d��A�b�9A��Jmq���
x�y`9
�K�J�Ӹ����ج���W�#JHSu��5iS���$�=�L���ix��︤�) ��BZn��^^���sJ���e�6!�&p�J_t�fk/��� 5ϕ�j*�N+J�V����}
����8�NU^B��jnU8�(7L5��Ñ}9��O�o;!����A"��Dy&tDg *��&�����$oQ����րBO��� �9�d�}�}|�ot�� �i2�>թ��U���x�{���,��SRo��n� Pw��/,���h�D���G�Gv1U�Л�Ac�
�U�;v�}��4�QBƹ$k�Ӄ��W��kX"K�[7k��؞�A�B�m;���#�1|�W"����a^VxWV]�sLr�`$��eh����WY=!:�W�"�BW���v��[����?��GS*v�T�͠��"է~��w%���rB8*�������:z�#0ϫ<��:��I�p�k�),7F��R��[[�{��ͨ�E�0
�������D��Y:��
�6�&��0}�a�q���]�x6�S���p�{�_��1
p��W[pI*���o㿜&��D��zJ���q�xӒ,�j�l30�L��p��'�6���ǿj�S:�[�츻� �> a��yUH�����Y��4�En��)w����Z��N��GA,�3��	[�6h�K@�&Kd�ok�v�Hr0~{/�L�!�"�� h�3�vu>@a�k��pV���L�4ɑ��S�j�-�����g���DzhB�����9��-%I�s�����%"-v�/ī�-�=�GΠt=�d�k3ʃ�*�^�	Y�!8i�%sy�k��|�[�9d�}ޖ�Y%�-[��3e\���犼@�����R䲍mtrny�n,��Ã����x��O�/���E�#��T�i����*�%⡧ۥ��]�~��y,lQ��	�1M��*�#'����e�+�l�f�(9�vx%���'d���9tMKd.���J�H��F��aj�I��K�)���x��S������H/��p�9�&v5m�C�(E,���!��ȯ�1����+�r��nT��W��[!ZZ7��;s�z<Z�g|��S�MGMf�Qw@�V`���}Ѽ�9{Ћ���DuTv���¡���}z-\�w���UsI��J|u�=�5bv�. �Z��SE'��3m!�Utt�%T�R��D';G��G "H�����:�	�g�5��"�����A���	:���=W�r2]Dm�]��w'�Tބ�����$M���
�����Z�G����z�!6w�Po?�Xē�P�m_��u�_�|�w��E��~�5�֬.f��9J�11�
����ym�Bz��֟V�!31��jJ�����L��t��S3>��!ϕ��n�YbO.j��͕�n�)�瞀O,��V�:^2�� ��s/x8�!�8��(XC�@��D�Hz�%���qN�U�qU)�w��*X��t���\|5��àh�qհ����|�;�C��SA��[�/�g�C�=�S(�2��Ȇ���ӉoM�'Kn� Ϳ��L�^���������D�\d�$20��i���6��ÉMU>E?KEӟQ�zy�P���1�l��п�u��0�q�%�Km���D���ʶ#>�c~s�(E������$��Y/%6����5l��'9 :�/*1\+6�1�3]Cls7t8a�@�_)IV���W�ٜ��{J��E�:��^�.!P�&�J���K��x��.�6��up@'^�z��H��4�s����A�6�_R�	��Cvu �VP�r�0Ցܞ9k���^�6^ۤ�����]�� �I��c�Oq����� M�`r�>g"���@�c�2��H�J��̢��,c�V�¾	E�<�cK1ﯭ��D�-
^s���j�
�;�/Q,�(ɩZ��3�M�k��L �}O2J�ZgE�C��0b��������=;���Ano?�p���"��X��y��6���;�����1����ރ��>o��쑆�� &*�Ktv��]�r��f��o?"�dJ�1�8��]��{���a��	�n�%�!��da%��F�5]>@P��Dg�J:H����,���
)���F�ݪ�^��
߂�4���Wk<�|��k�t�J
Z�9��Gi4��:D��䥣[�I ����F�Am��UE�~���N+:�y�4��=��a���֏6��:؅Oj�R4 �Ҵ[�g�-�͐��SÔr�k]�����>���-!������l�Ƶ��7!�ɣK��M��sPCj���6��%D�=l0��,��5�L9=8#�r�[���7�5��͝Yn���6�"�7���0�R~\l?d=5BQ��9j�G�� ������ ?�o�c�5c���-�L ����۴w)K���Qff�k$�C�.�J1�A��ae��T`�������m����Dâ̧��]\RϬAϼ�亂o[�0��S&�SS;���A_�}� ��a��p�����-��虂�&�ηs���h��5�Fό-�v�b���_D��{7zꊟ�4V�o�,�
G8,��9�Ҧ�z6l��Q���N)b���
/�Q�9:�x�(,�0ɜ�J�ĕ�k�-,q��H��JK���؋x�>�f��T����>��f�Jo�	�l��Q�� ���՜z��]?=�`5�?�h�0Y�ѕt�"��5k��εNd�ʾѵMOb��^�?�W>5�X��y���&b8��V�097�K,w8�<p4�Y!�s��$�� @���r��S@r�������z|�k�~�����ݵ얙�6|����=�A������
�2�M���W�9�!���3��F�#�(�X�6 ۱٩n�Hጻ���=8.�(nbyoQ�LxG%=����v�� F�]e�_�YS�=I���$�ɤ��Q�5�]H" ����UV�t�E��A �G��5]#98i*h%��P�f0�g|�T�� ys%Je�� �*�^�� ���V�����DD�p��4��Q�s�ϒ�(�3�#`3<��2�A��M��Ӷ`�-�������	��6GO���?c����ԏ[_��.������Y�f��0bOwҨ�h�9EU�x"�3^>���q4C��q������}ca��`��/
Duk�p>�m�	��d�"音>zř��`�Ԍr:;�S����Z4��Uv���-N�Ω�+�u<�@\�C�Wr����6����>O�¡E��"��\��S?��:�oo˥J��5�G@�4�s�c�0���ò�X��lvM��ʲ�� F�C^�L97�):�|>g.h��5�_˛�w0?ɪA�D��{#k���7�mry��A�5	RqP^�2޶��,�Ż@u~�s .����8 �[� ���U6���
�z� �vѴ����pc�����&@�72o�{�sj<u�!�U駇��
8��Ԧ"�h�����E�TE�r~�_��kQL�?0�+܎}�Q~����IP����b͝���H��V����˫����0�:�G�D�j妠J[S��k-ͮ16`j=)����v�AP��o�zc���O�����s��`����*���� ����UZ�0�a��{�l�~m+��� ��7�9u�p���/�a�2itPk�hiJ��P
#@�����xJ��Lp�[���Y/�&:zo�e\RD�}<�#N��s/�M0�g����غ�6h'���G��+Ź��?�PN'��w6�댘sƴ�S��7 ���K(+��Cz�ghOw��H���i{Z�ރIۏ�%>,�K�Ѵ���;IW��g�n�|P��\R��Jʑ���� ~��Y��L&ٕu�F���mV����(4
�)%j�")4�I<Ik��Xqw\������iȖ�����U-�Qi�I�(�aA�o"�L��MT뱓�o"	�N�췖Xw;��~G�}fDJX��q<>,�؅���RK`���U1$�`Ҽhm�����m��OO�A��G��,�"�\������0չ}Q��������RR@���HQw�B�'�67��ۙv��o�J��U�' z�u��?����J�ސ_p�6�!lnpS�!-��?���k��uoYK9\�nFͰ%}8���\|��j���Hζ^V�#g2�����n޷Q���]��kTP(`�c�8v�ƹ�z��k�^�x�VJazk�a��@
4��/�;�w���LO:8���S�gRQ杋!��^�Y 2���$�:�o�z{��I^9��|˔/Uʒ�ՠ�<�k�<���8l�>�Ɗ�);��'��&-���wﹰvB`��TUT�A'%8�T{Y&UV�9���5;�3���"����w!�����Ə�����>,<az�UIhN �vvF�=�ʽ6��m�r�+��B�Ay�j.��~Z����J��!Ɩj��:�4�н��'P�;HH�XXG�64I�*vP��Ԣ����T��m���BD��y�`B�&��U8�.7~\�0'��޹SU�#�����H��ޭݍ��i��ly�g���"���P�U����ǭ���E?8p��*�;Vܨ>=���\W�f4TRO������ ����a	[�Y]���V��	*��T�h��El���!p�4y\�o�'��t�E7�:^���!�r�)��#u�{UÖ,�bՏrA��g}�B�k��p��X1�Z��>��݌u�Z��O�[;�w!L���Ȏ�a�su����dF쒨�q �+8 ʢ�N P Ur�v�+��y�w��H��Nce�8,�#�c��6;(�r���mi����<��}���+`�NHnV��*��ޥ	��!����i��Z+,Վ W��pP14�����$�VB��f�Ϙ7�c21֌ѵ��\�Ap����U1���wu��mW{G���S�:55�B�M�,F|�67��`�d�D��=�p�qjє:'8wx��֔�6�B�:&�ۥ�8K�(�׍�ˣ�m�����z+�ٲ��p�,'���>�/���*����kD��]�vq���m�p~�����"��vp��H�G���/�Ct�X[�3����>�_-��ap���Q��>��_^��p�D!p��t̵�
i���k�)&j���\x�A�l�M���]xEF��	�Yg��YcD���+�X�uOX��M�O���9�#j,�R���4��s0�H��j� [Y=)��+)�@:�1����ߠ�	�i��E�s�또�U	/@��dU)v�0�������{��'�{m��~V'gj%����H�%ي= ���7K��O���h]TdK����n7k]?U�"�%��H8����;u�H�8�b1��`n=�.M�Y�ɧ��`����l���j�:=\�a�]Vo����ן�_���)Ff��������{	���H	�i����f��E�(����İeV�Qv?I�[���>����}������+����+bA�����V��R��ڭ��J� mۋ��]@~�Vg�I�;1#���Ԝpȿ+	�%8�A��w���|�E�Bd��|��9�8�?����k��# n��iRo�&E([��xpt'%y����f����\#g�>Jl�f�P	���n2k�󵢑 �<�'��)|�%�+�J�ynw��I�c��"�xǵf��� ���©���:�B"2�*14�,���"����	�F���!Ճ�̜{oH4��^Ǯ)��L^�t�>87@}�{\D~��]���,��D�Iq	����yS+y@rųWV��N���%�>�0)N�?B̩?č����y������EFq/|H�k�v�f���L�?�&��g���F���PM��w޲�w�ePU����18��G���ʀ�|;�,
�W�ۄ݁H�?GЄ�S9�e@�L��g[��;s��C�h�=�$E/Z
��4�;[f���ӜH���Qd+�Z܁.sȣ�%k*#�j&^5d挂�4�&l,���.�LvK���r�*(�{����!$�A�{|�<.������qL�(?�N��8�S,�1�S�8�J�ed3��PHJp��\�`��'n�..��C(�h���~�g���Q�7&��B�6�U}�wM-�����%�9>^�+��3P=�q�MwVP�ô��(��v>�?�x�f��Vť@Y�I-����d�g,�"�#}�{aah
����]贯����x�5 �l�z�׺��"�[�j��[���?�+�;��c2L��E�O�Ŝc���ՒJ�,���K��:���5���e������$.�ܡ��ب�Ԙ	zbU��{B�G��۷�3j,O�;�ʴb��8n'#M�(6D4�Q@��?^���n����`����¦K��BO4�`
<<N"b�f{R|���EI��@_��L��Y`>}���4Ѩ��"�V+98vǰk�Ô�ޕ�Q�|��75�tɒ�;VRdk���j�?��O��h��p��Fcݸ�9�)�8^Jq��=�m�[X3��`O��6�79��Q��x��7��a<���m߯�eIp����F����"ډ�����}&�C�˫��c��@�U���	�������vۉڬxBLccBƨZ$x���|Ӑ_4��A��jER۬MoM�&S5�jI��Y���q�]��h]"�`���iŪѱ�j�n��`+��q���8��PM~L���f'�O�"�����_��'�n� ���k��G��l������2�w�=�`����G7�^+��ܦ�����d j��b5�ʺA�_!W�D@XM���mT�,(�
��y�:Hj�_X!�q��(̛�4#�p�_�:�I��R)Û�{4w·T�~����m�![\�W��.h�ǐZ6���N��'%��C��][D g%��;+A&��Խ�'��ȸG��#�-V���#1Xj5�8�?}�^��7{���FJ�9	���p�?��he)�E�U����ĒL<��$y�P��A00��B�BF ��V�`��I��}#]w�:x9Ќ�<���0z�Z6�L������n����w�L�8��a]r����������s�<"��p#�؞qgW"�V #����"� �k�7�C�O�niR����vL�� �fk����=)�D4/Y�7�G�gurt���'9����1���~2zm����4_μ��0�-;��d�k���'w�p�j�2I�w��6t����ugE��";�v9n����+sp��l��D9��>�����Bf��P]n\����B������?}�,�l��L�t9q� �j�av��*�F�X �CGM��ӹJ�G"�L��؏�Ak���@��bZt�:�Z%�)�od�� =P�:��{�4��]ck=,��)O���۱�Ȧ������3Q]�C�N� �_)�����ya#oV�6CCe��%��lC#��2� ��ܳN!����NAX7)�CE�&V�@�'_��ǛP�N�Y�(Ŀ"#�p����YN��ˢK!v��Q��CN��U|�oٵ�n�C��{�J�!�ʣ�:�p����?�[�Ԇ��YuR�U)�����hڑ#��ƴѩ��.��W�i��R �QT�>�;&[+ߖwI�¥
>b���?m`���ZD��P�D��$t��U�L��*��p�{���_,�"������S(���g�]�8)��l{�lm�8ˢ/�`7+*;�D!�h��#�0��EF�H%���k���ܷ_1��I��+Ξ(�{��}��6+�0G�oT '��E��
Y�:���o��ivS�*`�pQz24�z����/��}�]�-lb�S
����a�삃~��E[��_�=�0��=�O�������ߖXj�<?)�_�O-�l>�Q��9GZc��Ym�f�HM%�K�AL���n���2�J�G�\�<L)�T0� �z=[�w^/5j��z
��_^�.Q���Ol���dh��Cl��e}�{���ң�G�8yaU�UGz��X]�UEjs��n���a��a3�8�h��{�q���TN�]�䓁|�ҷs.U��\��)��,��ZNC�xcbl��8?�R�H�y����=����W�,V5h;N����l!%o�Jz�kj���9l
��j�ͬ�6��u�@k�H85ˬ4����=�(kx�봸2�������Zoy�J1C��:�вB���ICK�U�%����>�f �P�^���Q�[ݸ��Q��y=��,��� H,醘�J>#���A��Z&	u��_��/0	��u\%���|�`Y�?;F�̂2�Q�pOni(	C��
xQ�$-�n��+������+�r�+6���~��ax����#&g��CYy��K@T$x���J�6�і�H�~{�R��hY�~��B�>s��_�YȒ&�"�7 ���q������FS+ښ+^��L�����.m
xT����~��C�8���2����J��M��À�I�B/N�3�.��.Sђ��m�L��.�m���w?K̸�,4�6����x�H���uojʃf���꒜]�G��:�d̒���Q�Y��P�Mw?I�Ѱz��\�x%�&���Q��#z,a��-�9o�M�����ڢ�lM3BZ��Pi �� 	�d�MB�����;�/=�.H~8�
��N�ꨓ��z]�\g�YnAQu��W�ժ����wX��z���l�Y9A)�>�c��4�sS4�p��|�e��(��yl����"X`��� >\�Q�jyG��I�Q�ꢊ+�>3<!�C^$Os3�-�e�%���x�7ٛ*S��4=��>�j��,Ჴ|hF�ɲI�*�B��%,렉�GC��Ed�j.'	�E�c�CLa`A�AC��~z��3��ڏ7x��1f#5�p׷�NJNS�������=#b��ل�$����6�iVq�&'@����ƙ�%� ��g���0��w�g�m��
@;M��	���&��kء�ˮ��\� 挃��@���)]�yf��:!���0�8� � MB���E�ʬ��M&�v iI�_܀Y�!A���<?i���3�,Rg%xxތ��ik�`�v�^�jZK�d���F�i5�6�k3�J�p��+]�ѐ+���֙:T+���î�U�"-�1Y\R]��Q�ΠW�4�W���`�w !�oY@�-$����k�Ԟli�J����u�[�Ow|�s�~R{��?'B������L��`гk��,�����|��N����axt�	k����4�yP�~PCIҬ��tp���t�`��7`�������*'w�65K�,�K���\�#\�1� -��&�K76º��}�`@���K�`�E�`�?9������U���@Թ�pp����HJ��u�7�'�F��.`��v�i^$�F_��
<Bm���\�MNYGʩ=��Gpl�3Q|l"/BOv$f��K��f΃�R������R�G�� :��E�,Ʋ1#?���I�=i7��M��9����5y�-�Z6���[�ٛ��k��|� �NGA�2����!7��5a�����}��t=�>���0�a�s���i�����m&�4�Ak� v�>dP�>!�uߍ�� h�x:(�e�Li?���-;�X����w�	�T~T�0�cr)���ݷ��54Ȧ`΂��ǿ6��ic���BD��/�6��s�ʢ���Q��CX�qVfNK�Y�Z#.����D�C�0���8�`/��N�H�4��L�Y�6Se*�_O���-5#J�����r��;.+eӈ����_g�i�"���+���u]��w��ur��<�*��R�n�J���p��h����T����R�I�d��2Z�yP6�a�n/���V^v��M��1���6�V�]^���FT3p�k��,��C�m���Nd;�Bq�"��w�Ȼ�b�%	�!�'�禡�b�Ψ�	�B�̰+�?�wI��ɒ�sT�Q�m��Z ϧ��q2�	�/���ɕ����k�V�;�俷����$���~*�{e{��Qg� ��~d��7J"Y-6�P��9"�!+`QR�>fD4CKn	��Ky�ӗ2,psZ
����dˆ�$b�VJ]������0�*��hdc�������e��-\��YDn̒����M����>��e���R0��n�fp�����A)�>����m�����ޭ\w̓��`Z��t\�f�3{�ḨUO��
6�-�l�[���!���*�N�����Z}�2��*7��0e������d�#�Ro�	�t쑯V��)��n!������+g��.7�e�Q���n�'�O"4���;:��s�'..��n~J�=β)j�Kj�	� y6�_B|-	�	�Z� &���,�^�y�∼��W�L���,?�W��M�ɒ���B����·���'#�����m~O�K�Ԏ��j F�Y)� Pܛu+>���^}��vֱ�ټ5��"������	
���	����b\U�0����ztr�k�Rh�k�gZD�*�G;)��^�;�yG��F;����v>��#6:���큟}��k3�a"�	�����N�ӅT
��IS
VtĞ3����
!�P���l�e�o����Ď�gBпs������&��w����l��:�%�X��=���tD�dw�)��[�W�'!O��%:�@��H�⑊g1f�z&���PyT.�������=�~%�v��2����fkʥ��F;��
gǘ�&_��$�����/܊;�!��*p0��#>2p4t�rfLYڣ�>���e�yk�Hq_��}rYs�xu���xi0,@����٠�n�`�4Bn�׶��"��;��[�ȿ���u�YN��2�}�na�T��0��c������O�T�§ݠ�,���7��bs#(�:������ez%$�"k�j��&_�2���kBX�wnk�w�J���Kk&� �϶w��	71�
l�_�J�o�<�!��Zf���חTσo+�4ϡ��;=L6��f��l�|�߾�w������ͭ��9];�����`:0�ܯw��V��ˋ��������F[kq�R�/�t��(��v�Xi��O�Jψ��*&�VJ&Z��̬[k�Q��1� #�{fv�b��)��\�"MĜ����c��`�Le����1lK������Bt?��A���D8�B�E:���:�� �g;�/Tֽ���`s;����\`y2�ȇ���z\���h�׸���T�t2�a��NC��V�HA(�M.W�~� ��|yKY�� �/P�@ĺ+��$��`,
�]���3�LG���Ov-]��CcK�Pk(Fj@�@�]��%��]�_�ñ�I��#&��MZq*�ġ
�m��]˱WãҨM/L�4"�2�R:*EVc��)�����ႡM�
�`��#u�e�|�]�<2�:��� ��U��|HX��Ud��#Yg�#�RnK�h��P��h�͂A? b���(�]�U�5@i�w�%�yS�,��oQHʄ���u�m�ox�sE;���X[��}f�E�\^�~��=󦓢+�"i/�gՂ�<���n��
����L鍒{L'���P���UR��f\fp�Ju٠�s�ScY�B� �����:��/[ϭ�wGA5�G�MZ��u��L�����Oq'?#	B?-<]+�Pj�����E~6��٥iT��y9�t.M�������¡2�c�������X���;"W{�oo�pfK�-��)�|V,-����:�t\�Q�8�t��E?��6��{Q�t��"l_A�\0X��2Y��\lɈ7��Q�ν9���63������fKK�����oPe���t!�te)Y}f'a�d����1n6�3�v��h.�ve�Z<Cz����es��7؈�s�X�V���=���M&�lF�C�/��#�E"�I��B]+QD�.��آ�4�"A�D<W���[ٰ��-��-n��C=Q}F�˶�L	K
p'˸=����4���wN�7EF�]�MT��:���):$i:jj���;���>k6��"�J/��_��Ɏ�Q���
-���E�@����O��0J&�h���D��>1oB3�
�p�cS|H߷�'ve-2
�o�MR�����쬁�j��ǻ2����	�n��q��7��[�;���ւ`���&x�0fC��,>S���?y���y�B^�A�R�o����(��^�2s[�;&&��dz�j�_m;�+Ѧ���(gٮ�4ٚC��D��^l��G�h�ώ�OwN G�ҏV�FOޤ)*��#�#b��,:�J[����M�cƏ+��@LP�T� '}�b�<���?�|=ɛm�u����G�!�È��|M�I�à�-�F�Z����h��'�rQO)���Z6�QC ���@�-[INBX	R2!�.E��E~u st���~����|,~�& d���!�=WP(5�<�)�^�l�c=���L�'�^��
��0w6�J`zc��ƞG��V��.C'���h!���d�ͺ�D7��7ҟ����+G/�`��c.R�	��7T?6P0S�:�LAY2M�j����Ĺ�F��B�����m���LWb�~lW_i`�TB���s]��ja��bf�L��Ī8�>�
�_$S�������Ln)��o��G;��%�+=�<;9!tbV��λ�˺����[E��r.��Eێ#W����h]#ۗ�4���_9b�K�Τ[Nݷ�_%�Kc4r�@��o?)�U�fx 0��D�Փ[J��'$��|��ˢ2dn5�.܉�'����9�|Yz����tܯ��ݕpʂ7�:��䪆� �z00��m�c:@��U7��U�Gίw6����Hu�~#��NU�3��7h��-6@�m�9w�{u`;���/��צ$b)�L-��'����O��Ixu�;�L�a��D��.]��|pB����aC�O:f�|Mdʌ�֝�f8�z'�T�_8��h��Qm2L)��'K�oYo}�]i4ߑF������C�����kF�GS�C���d���k7b�g(N�0J\2�U$]�H����3T�*�O���`A\̀��f	S��{f����|	x�A�<�� ���ֆ����"� ���爭ϿD]{a(��/?�=�Y���/�(��4ڂ��a)�hڦ,�k[�
�h`����`F^��R�>���XmW����0�A��	����.܎��⇟9䶚��p?�(�w�=��l67�2�j�	�V�u��$k�wó@��L�i����	~ˡ2��T.�a�B�Mw�z�|��]�c�գc-�j1�2�����EN[����i�%ǀ�xa&����!j����Zw�d�qru������\��qG۷y�4��Nߒ��X�L��)��B�+���޻��Kcg�I�}	�س�����F�q�^�r*[�T�y��2jHP�Z�G���'7�N���N,ca~xRQ4M��dh>�}h���8{?X���r�/�1<gf|�-Mg��ů�J8k��a	r1A�O�o�xӁLm�Z������Q��QH��ei����˄*�g��)�F"g����)j�U�+u�e0�p��8�,F�w{�ڬ�F�(����J��j_�R�C�����plː&-Yi0�\��s�h�)cF�	�RNf�߸w{�m��H)@��*tdO��%XIƏA<"W�}Z��Mͫ��1�H�X~�tO䥣��я�>5fv���A_9HPWF���&y�G*�.i>�hf�Y��iN����S>���NU���p��WT�sQ��R��T���twE0ِ���%A�qzǯ7�dD��IXB������������o�H#H:K��1-#�d�b1�G3j=rp����i�� �e�IP>2��o%�1�Ş9�	��#f��-�A#��ad���q��VqN�[&h+^�$�լt
��pHi�r��`��Nį����C�Z�WY����DmC�v�
F ꡚo|)�VZI68Jt+6���g=��-�cugi!����~�U��!���Ym��"A5ƙ#��ԗ�7��u�da*���T�=����Ȋ�Z<� ��y'فW���sD��p�x��� ���F���L�c�x����wƖ3����MN{,���88�K�3N�K���&i-�5σ��V�s�Xȯ[�D���Q��iӒ�������V/V�Hph;nsl�?�����������nQ�<�_Q�����F�I���B��Yff�g�e4a�3+�K��0����yV/�F>�+n?;جB���;�"%��=��D���q^jG��_��9������c��������_�Qԁ��O�Q+-�:��1N� �<��4}eI���۪-bnSqVڅ�����,qQ:�6��&�wA�+[�Ѥ*��F��GE�v`}K�j��s��Jٝ���ht���j�0& �1gb�+��o���h�.׏���5�C_q�nH�q$��S&e� 2������c����ʮ�h���p�n���cXH��p����(3w���<F,t����>���
OT�zmXD�q�����W�-���ye4X��'�`�dx)��[V��޸���I�d��=�ښUJ	ʖ�kρ���44���H��⤁I�3f:���lF�7x��	П��8��tu�U��{���1+k�P�����v�|�1���|�y��ܹq���*�ȫ�a�B���0�^dnT�p�<P��"�r�)pn�˫>�ּ�VӔ�<r��er�G�a�t�n����[�X�1C��M�ɤ�ͻR���i�͡Yi��ݸ&N�Qnx�י"52tq�^�vQ�����h���1�>�g�Ku�p#V��!>#F�}� 1JPɤ��������&����qE����;��nMT���:�(6ƭ�O�P
�`�,�<v"�o%n����\�d�>	otIy�sJۚW��B�[A��+��{�?X�d�==��s޹̳XT�}"'��S^�r�A��n��_����K'�]T�!Qzo�k�cv��(�̺5x��p���E81�;�o�Y���f�P�v��X�fg{;��6����֞L���$}���mJz�����}�'l�?B�V�#0,>r��M
\X?�#����C�we���A�1ܖw����9mu&q�*N�����픻Яq&Ond?}i��x�} 9i�U
|�,�`�@��w��Т1���r�w��P�����ߟ�����鮘�z��W��U$#�������\쳔�k*޾��72��c�l��ѕk��Ϲ��W?�0u���:�_w���H��*��M�c��P2�����ɛ��.�ά����9�K k4Zyw`*�'*��	e�b��[��c����/d8�Ԫ�1ʛs�8�)6�p�%���+�Y�@��l������Z�N������/&�S��{
�"V姛�I�|���r����F� �8O��p��8f����. �^H���y�<�Ϙ~�\���)A�O.�Ӻ�<m�-.F�h�#�S�����2JpT�Q[Wdf!��O��D�Ѓ����i�OױU� 6��XN邺 �D3~@��g�
Ã�Ud]<��zl��Z_�"1�|�ٴ!��,+2N4ư�Ԉh&>!���ֹ
��z�8k��h��X���).�����xɝ	c�3���Uxkp<'��$�} ����3
�3��X�N|�D�3�@E{+���!�.��<�8')�`��!s�K1{)tf�گEx�n�=�G/'I,w�N  6��?H�)�_ǭ�*��+���C�(�d��c����1��ΩՅ��)�y�� Ԟ�%���  v�ଅ\���R�o�S-�5a���oe�}ݑ���ͥZ˯&��������m�����y ,97��䣲Ѽ�v%�s	j8�Td �@3�K/���_\k��E���0�fp�Pn�z{�dp����|S���Tby�� ���nezߵ�z�78�f�V�Y{���G{Ȋ�R~7&}���\��ҭ��a���o$�&:���%ϕ��\2"�Z+����r��sVg����-�x�N]��;��l��ș����}���G�
<&-G2�����]�����������3���_߱�{u/�En[C�<����������F���a`�R�EH��ء&axi�u�e��z�O�%��"Xm�}R�yLV�sA�+0�ѓ�������#d��NT���Z�{j�/P�Ê^���ep�0แ��cJ[k�T%��ꗟwKL̖_�I�O'냬��"����'�䳤�j(��<U=�f�{%�ޒ�p/Ѓ�A�Č��Z!Xg˷���a4xߙ�P��x�O���]�~�p�ĕ׃�D��/�_U�,�%J���/H������yM�U��0(6Y*�L��aqr��z(3�#V}�u�Nx �%����o􅉡�V��g�]�=���M���6uQE-z���=t%M1%"F&�4�[L:���2[��:�c�zqj�(z>⦡+;�V�:�_�{~�M(�2U�p�-���i�����N�X?�\�1G�����5 ���&Y�oe��FE��.u٦�x<
��Pԁ��f�s�<G��b��i�v�[7�T��q�Y<q�����{�]�t
�@��"��u��*�b9���|�m�;R���"���3�1I�
Á�����n��p==�r5�����ܯl��&��9lV)j �d5v��<�
&�K��Z!�7ٜ��A�$�l���%;iZZ�����@�_�m���ם�}��c��C��8��ыH�X����9���?�T@p��T?�ט/�I����!�Ԅ51E�Tf<�*�sI������vF��L��*��@�z��]'�j:�Ȕ��^9����C�^� �C��I|�)���{6Ow2���b8��q��N1��}���#Y]��~9��؈�C=�yJϕ��	�h&�������I��hr8�Z�[���wCސ8�����?�҉zwk"Y���2}57,�V@���6)��ѣB(��((�\zÜ��p�!��Mc�>y��dy�LZ�ԗ.���ه��fn\v��`���qh/���!w�J�?ɚ�V�cރ�J���'bسdVZq�����%TJ�|B	 �
�Ȧ>I����Jl��A��T�4h�&OE0W5�Y���&>��fy���t��.��jK;�3��E���J�;wC��z .ӝg�MO=WtW6�xg�9��a�m��ˋJAWI�1H+ٹ��zmp�W�Z�TD' ���Q���v��)&q��yL��B�J:XF�Za%�F� �ȴ�:D�|\��+�ڱ�2	����j��A�>�JAF'Yg��yF��J�cj�����g�= ω��RS��sR-i��ghѷ��n��͊	-�>?8q�$��֑3���f�Ҋ�D@ �jCP���U抓�qD�m3�|st�mV�;е@Se)��ʫ�3Z������|����C�\5P�f���Wz����1	d����'u���d*{V2�O�Ά?�{xjX��
V9�P�k������X3���4�������}Fa�%���R��=���fK�1� yF��H��<�w�D'�dn,pL
�w�Q�N��u:�� �"���l��3)V�Je����T�����{�~bC�U��_`���|{�]^
�c�i�'�vRqu���k����Ѻ�ߋ��1��$C�$	g7�:?��v?�|��4��K�mle+����q��*�w�t��X��l�h���<46���[���D��G��(Q��B�=�DdU�K�&!���֝��67��$���qiX�)��5a�y?6x�t�WY�B�,�Vj���?"kOP9q=�kƗ�A��P�/�=���|p�OJF���o�3N��1Y�#od�´u�t�^����JT%QڝrL>��@��k��-'�3�ف@�l�@$���l�f��
F	G�8����4��#�ͰX�z����[J5���Ҿ��(нj�=atP����6��J��`Ks��"��zyOH��q��FDh:G�0�B��a"�VVMU��R ������� �(���|35Ԅ�ej���wxc,�2�$LO�a��MN+¢�'�Ҝ_��s���t�0Ҩ�WD�6�ګ�_&ɸ��Od����z�o�$S�|/�t��h��f�A���ťK�y�X�����\��%!d�h�W)6J�C������ $b}�-�<�U��O�2�'6o�ֈ�8��ς \���s@0�d�lv�G f���*��z�%��.��N��<�ߺ$$�א	Ϡ����6�?�M{sNbc�eߖ�Z+�z�Biy�PlA�Ղ,?�W%�К���Rc�ؿ�&�4KT���4�Sɲ�_D�t�d�a�J>Z�<	9��.΂v���[|6�M�[�����vn��fU�UM�D({P�Fis��ꌎj?���q2��_��r��d�bEצ��N^q������9�Uv�.	Qok�����}���=�:��&*-���q�����4��2��ΆTlv����`��"=-�=�}5��f6��U���ٲ	0i��׶n(���n�
Q��O��d�#jF3�m7o۷�S@o��.�	����AW�"J����1ѩ	8�Q�� �y*Cl�K;���Ə�؄�,%�����ǻ]��^������W8ZC7=m�!n0��L�%�
��Z��y0{j_�u���;�\�� b�5I�-!)>晴��%�����cB8���,w�J�
�����������`<����и�2�$S�[�Q2;�{����Ap�:z�δ�jO��j���k�C�m�+�ꪼJ�a?�=��<��bÈU���1H=��ּub�)��az�"�����u��?d�EVG Ǩf�ĳ��
*��8�hR�-e�ixz/	��9kB��Wm�cH�X�6�O�k��1�lD�)���_�W�1Yⷘ�^l�e��g������2!����N
"�<�q�l�g�L���K��;5s��!��҈l�I=�+�>�ꪺN#���R�-�53��nxd揁��Xm��kk�t~3j��X�}uޯ����I���_����
���zĵl���D���{�fN3�jy;�rO<?��:	�E䝐��:���48	�(�E(�&_���RE*t��R����a@pI.DX�M��A��-`���X���u�����q��^H��]!�}�{e�b�У፰.���+r-�����Lм�ѣ;�mzL��H�S��=�r��FE��T:�?�9ir�?g�૸��f�Ȉ�r�r��-���69U죑���T\Eɐ.�>�����mv�
�R���\�kYJ'�!l�UMT�(@Tޠ�I�?�d}K��<��DIA(<6<�W�15Y�]�=w��ũ���灂 u�P|��xe�du1d��)�`N�M"r�ީN㸑P5������~��&L���������<�Q8�>���w�V�޿j�K��v9�"p�����	;��A�d��#�c�q��8�:
���"�~:�����R�o���m�9[�
�[W�j�hr�l =�)���W��4#'����ڣ\���#�@X��+��8[��B��3Gĩ��m1�I^��g�|M�:5c[�YUDơ�II�43�%ȁ#�.�� ˝�B�}-�"�W��}%b?;}����Y�άp<�NsH&���A`�{���p,�Ly�1b�i�Cq��8W]iz�$+��8���f��a��?����>0�Ʈ�}Z}��<qV��ƥ����Y\�.�&e�C�e�& �erB�Jt"]!�L�����>99Ad�Q�槀d�Y ��|3�-�wu���rs���E�� 1J����jy|!v���P��`*/�o�4Ll�e�5]e/i���&V�Y�A�T�ݶ�	��Q9�4������,���Ŭ������mG"3��N
2�m���s�h���;�*�_�:����J���8��W�����.����l�e<T�(���Ci�G�xݖ6���\l����8S��	9Vh@�s�S&�f���%l�B�T���%���I�l�0���nX�(��s�a~����u��B&+p%�a�C��B��t�!�aAɺ�F�#|a�j��Qu�5����1��+�
��Ƀ�� �,�U!iFW��ß�
�H��2C�����}�}|C�! �� �H�|�#'��m��
��c�#%mfӑ����H�kM���� �z�D�鮚0?sD��*�}[5KV���Ϊ�n������<�#'�7�.�rc���X/�j� ����[�}�>�R'.ٍ��\p��;cs�� c�etߥ����P͞�Nآ�����0�Kh��B��E�:h�w���PpOG#�z���ޚD��g�K��K�ģޅ͚��!�s�Q���z�����G�{�@@��k�̍��c"ȸ٦[���7/q�@E?��T	.T�N�4eT�DKY�'4Ev�rA�s�5�~х�N��T{Q�u%�ݣ����A����e=���l�]X��=S�|[p�T31h.Cu�
N��u���=�4�����Z}l���}o�Ѽ#���r�,�s1�̚��sm�F�1�:�5|L���>�b܁Y�j��S�b��j�$���G-{_��z�N�Ǘ'��'!Ļ �7q:�D����=&�ܵ6�ȫ�2��yT�;=�Ha]E
c�.�"��~.���Pɻ�z�7%A3�<��L��G�s�s��)x��/E<�cp�R�R�a@�!�����|����h۪�H�Z!�Q��/~G��d�Ǎ�Jpb����s�y5��	�1(��yvoe�e� �6`���}:.1L��#��b�b����m�+��}�#`�Nmc����M�> "[*�A��_r��V55g�?�R(rO�Uc��f����(�H1�A�^�4�N�H5�wp�"�{��)�Ii	=����p-�`I3K��x��M��x���?u}��
�殙����Nf�VW��&��bђ-\�)�PeVvY�����	����3
eny\�Zʘ���谦W���1��fbt���8���k|���*�O�7���_v��ZcF�b<:S0��� OGj��tN�9��Sv��ƌ"��~!��#/}W��;�!����pl?^F8p�u��p��B�����IY�1��u�7��Ymk"�8KT$
1��,�ƺ5�Eqc>�Ď��C.�HLz��۫k�H҃'/*��ݔt�-tlR���i����H�������	��ב�&���T�H�'m�-���qM�,S���c�m��GEf	?Ǐh����K"�'�����-��1���zV?�Z�V>ؠ2�����$�y�VY��p�k"Q�rо1�oL�����Ux��O��8R�ͭ�&޻*� v#ϓ��?������ m)�a-��9��k|:�=���0ߑ't�/�&&�_��H�HY`�[f'4�&��A�Q�((�-�䡩"]&�pY��<�jN�V1C�Wx˖%�4�ޯ� <$�tV�����!���^�H�h�ĥRj�����0�:�qŻ����E�|>R�z(���o�ó5��j����uͣ[q��?������v�P���-�tp��A����֧��XQ�k�B���,�e	��%����<�*�p��#�Ď����{36�wNȃ`VS���}J*1Igc�i����$FSp0�t��]uM�G�!��T�%34����\�J�$�|�N�s�8��xW��IM{�IC���i�j�[��8r6	U��RD��Ӿ24��,�������yq	���)����4p�l��T����"�n���Hn�#:��,IeP���o������A��5����:���y�n�j��a�,e��Nظ�h���	���-@A����
$`]�t���ǟ���OEk�NK6����0��{�`	o��I+6l ��B0� �]���?�\Ӧ'ҥa������e� �Az�K�",׭Q�&�j/��\�/"��:(a��531�C$g!;��@��˖U�~����8�QHn`�0`i��`K?G<�E� fC���{�ɰm	�T�~V�M��Y�p ��V�Mh #�u@	@N���6�����O��cɴ�4���؃LYis_�%u�wZW6a|�qj���p�A!�����8�L��+�Ӡu���\��})�֣3�*�:�N�m���-p�\g]�o/��r�)3�ղ"lm��x���J���P4��P��γ��DU��S��i���{w�L������ !������*`�t�[J�Iu@euG
hq�0����|�{z�o��7ك  ���U�ߎ��w���o]��Op��C��m��h�� �~�)����oq�a*���%l�S�A$h:��Qޞ���8�%NPC��-2�Am��
�8��& ���"
+}�C�r �pn,�/�����5�m�n���ঐ��k�0%���ӎ���2^l��!v>	I�=I����Fѕ�
�y%��A=3��SY�HP���X�~lf���5 -��1�h��o�:Q���FQ����ʉ���|a�(�%�$�����c�\,�6��
�t�KZ�WM�Ǧ��{�v��Mkr�Z�3\OA
W���e �-Lq����{#N�ma�c9��7 ���'$��i	Le��c�@좧Ct����`���+��m�T�Y$�!�?���F���� <����|�)�����{��r��X���OĜ\����x�J{��p*9����%�el[r��LƎ�8��6�+�a��Y�|$$p2޶�m�+��[��4(�����e������?K�A"0��\I��F̻�X$�k�#ى+X��Ծ�<��^|�� �������o��؉�t����a3I��&|8�1[�;��/_uI��6h%��ADK�j���Dw����7����Ȩ����6`TY>���h�Q{�ߑOz�A�Q�K�"Y,�+��n�ax�C�~L�5`����3{��TH�|LY���V�fB������M�KƦ�-�j���$R����9�+z̽@�ǲ���E�3���[��p^n&BY��<3����܊�9EE	��FӽG������P��M�NX�~�tR��x7A��k��P�: �n��,�*L�0Ҕ�R$@�{�iֳc�"iT��U�i�A���[n��XXb(lP7'������NC��=�w0_��j�9�D�CM�9M���jv��3{��Pi?	�?� I�?��9���roz��h� ������0�}��_�ލ��,h�T4��u�P�5�rv���g��/�W��&�2�x8�Ю%I>Mn���S�S���_�'��1GV׈�z�<>��(������P1M!����ɽ�B�u�z�	���5k!�=�@Qu+�2�����sP~�4��X}怃a,,����2x��;]�V"i�
"�h}������Bm�\��Ġ��AugN�~��5��M3�![�P��f��H��7�5ڝJ�z[��ԣo-_�P{T��u!H8���*�'r>qA��j׍'o;���BZ���'���@S��n��]�G,���%�N�߿[����A�|����B[��g�o{�e9�G�e�qQ�{�~:�$!K�xB�nY���8��S�t�_�c�9�4�b��7��������p���]a�����3���I�b$ʜE|�EW��՜�4��S���,]�VB��@Q��,68���6|i@���[m��>og�����PPPL�JH��I韜�H��餺�3y��&�""��>�1UX2�q�Gy�W�do^>9?�.���`��/���\g�ܹ%$vС�l6�8n\Z�#]d����H�+��[��S`L�c�O2��=�X�Ed<��ȇ=X�ZAx����"���F�<N���F	��4�+(����/Ɉ։q�)bG����(_k��nZ���|���k��J��M�DC�٭���,E0=����>J˩`��en�D�D$9���oDu��Z��,��3����=�U\��e"���o�5���<������[����3�}D����9�eIp|o|�ۤGH{@KX��C��o; �o#����쨐8��T#i�=Bz�d�žL�d���қ�M�<�ܞ�Q6.ZQu`W>)�,�eiu6�ܔa���������>��k��_f"�䥎����ܵ��u�~G�D�ܰ{"���F��G��S!��xRN���6�e���EQ�C8���c�>�+�>���`:+��hKfo��8$p���z�/�P��d �&�F� 0�K3����k�ж���crt���91\���S'��{�N�"bQ~��V+���2�n�f?\2:�]Ym8�}:�B_K���a5��{�(�M�;�c�iGd�Tt����:��f mFg�3��\�2�ddPj�������_�U��@��u�E�dO�D֡ߧ^�d� Hxx����p��n��IR�H�A�NeY�?��pT����Գ4fI����}ߩ�1Cf�b���R$E�J�q�6D!�\��[n>��~qWy�߮�W,`Df?�a��&GN��O2V$�i���x�6[�e�@3h�'p�*���T���E�����Q>��F�V�s�OX�wm�]c�Kt!A�߿��+e�Qs�A�[�L��i�f���Tz��,�� 
UO-���=�!:�o��?�n����6�#^����ƌ�<�ʻZ�Ui����1M�/�D�2�$��Uz� �;�����^�&�<l�����F߯�6�Vc̪�����t���teX)�-Gl�������Ѐ\�6��e@}s�ml�Y������<lgt�ـ�~���ᮻ�pR�h�\IىJ��3J�m���Nh���(a^IlV���J�����]NXKm�m�c�y��:^ �0U�N`��n{82*�H�ҲBl�nN�7�����j�D���t�:x���u�@�������u�b*����������ǲ�p��!>ǔ�����^���U$N�
��C?0�|�q��O������-)`^ɲEHD��ĔB�8�@T	Q�}s��/p�LS�-5?zO�[������@M{o�u�n(5��o��s��4��;�^f������Z�l�C���o�$�i��Zl�<g���4���Rq��f��Q�gw
iIL�
�;����V�w	�=N�I���dB �-���%���@&:�bf�$�E�\�]�#]δ�����z��=����
��
a3x5o&KLWW�G�ۂROD�-�ҹ�&_��Os�d�x�0܎n�edӆ���y����3�h����4�*���]�<V���>�𐳛�n ���1Ȣ~�z���I�"�n�޶�t�54��[\�Ư��U��A\��ϣ���6��8X��v'J@�B����aa���9=����@�+��DN;�Z��C[r�>��09����ģ �rk�	'�p�+Ѭ�'�ľ,!�����Y�`1^�1�Ftp�i�,<�t�Q{�s��Ą�[r�{��"��yV�7���E�W���'<����	�$"�ugJ�m��|=��9.�����K灷.�Cx�S�J�a�y����)�S+Gk$y�V��Ǐ	�c��@����,���=(��	�<���=�T^��d�H��b���KL��� 90R�5�=�/zl�v?�.����pN�|�<���h�qE�!�����VƲV���Y~��P_�����x%�7lY����~��\^1w�����:�q;Ѷ��,"��P���Pa#�p�(z�����G�h��{�5N2	^^0��K<h[֫B?h`�]{�6�%ͺrQ!N�66��E;RoF9��v��ul��xd�4�t|ZN>M�0�G�Ͳ�߄0^e�Vռ��.zʫ�0G���oو�Ϊ���U ��o3x؂�%��+U*�Cd�:&e,�|J�,G�����w���;� �1���[��r�,�P�vt���}���F�p򜺺h�w/+��JgJ�Ukþ8n�3��Uvu&�'elA�M��ÌhzLd����󝊄.��lzH�d~4�`}:ͷ��|'���J!���.n�V����i�Թ�1��-ܬJb1�F��a�ؗ���(�����R7WM@������M-�
�<����8�=����h>���q �/�Tn}�(6��R�sA��)t�1Y�V�u�Ҝ8QhF#�V�n`A�ϐW����S ����~�WR�'!e����<�U�o6�x��n`�#��4���z��Et��+/%ymȤ<:t)�nv������De)I�x��HA7�ex҉��ӣ,�ȫ9J�x/`���Ew��iַ|KO�W3xj$@��(���?y.�������ĶC������ƫS�$vޡ��r�/��l��U���\��� �����՛�D�U�,���z�c�d2��]�R:���4�h��<�1�� u�1��{f}K�0��>��6�9�7�P��9����9�WK;�>�:�m>��K�1�G�:�.�Α����H]����w��ȗ���X�ʂ��Z�	s��]�����\Dǡl���'�y���)�*ȩ/��!���R��3F��w��b@'���v�tb�<�~��*���D'��{!��'��3?��'�,,�Y��1���0(�#�:��2��G�e���88~f���U�I_��Я�sg_s�<뼨޸�mr)��𴂒p肵�|h?�7�c��tFFt���GIo��hx�d6y!�Ik�ƽ@�R�F�z&�6_�t7���\��YQ��2=6x;<����xmٓſ��f3���+p�u͹h��,#s���� g�6� �q�kr�Gmͽ6Ʃ*%Ce~F&��]���vγLw4��Dp�@H٩��d>�������Oݘ����خ��#\P9�a+պ7L? 5���4��jw2���]��w����ōk�� ���۔�������*O�4.��`�3�����/�,u'Q;��Q��&amB?Q�T��Y��o��T�X��f�%�p�� �!�~�C���ϱ�n����&��D��ԁ���u_�RJ�u���"�
I�%[F��P�b�f���w�/lGVC�p.!�~0 <���h7x��C���A��������8��ͫ
�=�v}+D�cp=��!�NK{;:�a�$��d��3�D���*

�g?��쏝i�0p��?�x����(������]}���/ˮE���l���I�5���l�1u�6�b�H`k R�J�Bޢ��!Q�i.�[�.3r�Q�k痚��3�sQ!��.�����B�8�s�#:!c�L,�`��}`I��bD��Mxc��z�	�$kku��(Pիڡ�X���-Y
f6r�d�-� Y��8i<
�S��`0�<�1'�0V��_!��>���j|g��U�)/ߖ�6����[��9����|(��9�U�b�7�a;��E��\἖ߜO!D�ˉ�M���c@�x�r<z�����c��Ɠ`��m�Z.�߮BAQ���uס/sS�n#I�
�Y:����������.�x��a��e�	��s�%T�&f��\I\t�s �Z���ٹ3k5#S_�X����b��s *���JEK��p��9J�S}�'�>��'n�B=-�$V�M�k�NO�T����[cJ�H�*W�HP�2挼5����k�#��P�-����]|	-�%Пk09'èA�c�ڏC~�k%����G�[�*^�����b.�8�Z�[��n������&�g��Ly�tI�gZ�*ǸE.�Q��\��<��?���"�l���~�3��l��y*�z�r�؟y|f�S���(F8����(P�����}vd_;+�z0y�zL�x� ׃�����xo�״�O\���N ���xe����b.�fޮ���{(�
=.n�����W����S���Rwqh���qe1��� �C������J�J.܇y��-7i<)��d�.}͠����8��=*<���V
2'iө��V�
KEk�P|k:�Ga_�B��bY��X���J�����y�G�BZ�f�:�y�8/QD���aW���V@bP���~��,�m���s+'���B����������������f��¤,O����NF,��uā�s�&ЌFH<�bn9�\�(��{&&e2\hN_E#3�����Ln"��n�ؙ�nV��g��i6��Z^,���Yi��A�6fŐf�%�Yإ�S�vA[_S	N�"�m��T�x���C��[�0s�o#�R'�x�y����IC��~(���)�}�R0�"�Rz'IZ-<����)&�4L�9)π���$a���6\�1ԧ]�C�*�ۨe摷r�Q���J�����bE�!	"�$7�yV�H��Wq3�T����c�O禧�R7˷H�p�$�K��%�k��o�rФ����2��Yſi��!`D�{L�%�`�v����j��`9���$v�""�u%	�BW�c^�/bm!�ڮ�S�9��� �P�~q�HH��|s���'�}��W8� -`ϊc��|L�P�ͅ�J�1�␬X�S�:j��8��.L���?�/�|H��*���0����2	�m�Y�sJ2����z������ 8��%Q��)ƹ��]K���s�fg)�tՋT
�����1�
����G�f𳮨4��q���o�<���/��j=:��c�4�I�Ή���GMk��-B7�!����-�U��v� H�<`���HD�����i�������̐?)�VxL�ǯm�6�����bp2F|�MI� ��]�249�I�^�Hu��6D���RB2�����@G�=w����@�q�!{QC��� ^���`YbJmAm��@a셠pн��S"��L�ǝ��
bNdv�5x�3}��v��a����"�������#�.C{�vql���Mǿ�+�
��K,	����\�G�����xg<�c�$[-�6B|y=��*�E������U�hC��đ��Rq~h��J���(�����Y9}��?��StV����}�q��Q�+��!#��c����v����*;|ώi�YI����Nt߇A��	�kȰ�~��ô�+�Wf.���D��S&�Q�����rǎ3�H�x9�>^c��^q\�>�2�;�3A�z*�DnVbֿC�"i�(�U����\+e�Ƃ���bc1*�Lэc�(o�1V��e:6l/�J����CI��%�F`6��$��V�VL��3ֺ)w�y�U���,��*�G/��k���PY�����O�7��/m:�:�w ����`�~B�\���@k0z��ѸujT��G�2t~��E�6�!k�Aq;���{I`>��J��6mLB�k��r \��3��l�wM`E��E4�N��9������jhEʊ�s�% NԵ�Cz]??{0��Z5�Bպ���Ť�iQk�`R�>���U�C�os��b3½��.��H�<u��s�rx���E����ژOV2Ns�$�i��p��i�Cx�a]����Y�)Ej4F��@�v�2��3�H�(�ߏ8�-)rij�����ޮ�
^�|C��<�a�@ھ���@�)�ȵ�����ڤ��2c� W�9�K�;|�**l�������d ��f5#���(�͇�=���FJ.�5VXS豹�R��7�[����5���7?�3�tMBDtl c���C!mP/�rF�zF&�T���i��h�|F�?�+h��<�r[�<uw��pMaP4��fh���;-ή���'jE8?h��-�+�;r���\�7@��Da��	G�$�k�[�GC��,�"�.��k�yp�����(���%��T�$C�D��h^&�4ag��3X�$��+�^d���r�$Z�9D�I���z�=@����[C��xV�KZ^��t�%�kg:�`fH9/:Z��񷻵l\|q���(|����.��Dd�G��b[���L�6~W��m,)�ͶՠV6B��	���P\�mPo1����^��C<�f'zk���2׌ ���Y�����t"-�\�2~6�c<_7 :���.Sa�z�d���c�L�Hw�!4j��O�G�+Ѫ��㾠�H���)T���+RuS�rx-R�/�t<��"���?���W��>�MMqH�`^-A��;}9
�KY�m޺�I����� ȎO��q�;ı��*0J��������d攝�xdU*����k��^�SM�f_ܯ�q��*)��BZ�9r��<�8��Ә1^��N{�<G��T'�f����H���hgp�����a�p����5�ʎ���<.I�y�P2��4���`
`쪁Q�N1���+�0Da��h�IU��TSH�d`,-�v���fP��WZ��($sv=º���`�o��I��{��weA�j*LZ�G0W4): b&��?$a�
�����(ɒ�`QRسc@�m�&�gn���R6Q�3Vu��܌�J�D8^�A$��Ko��K ����,#o�9d0�C��}g�[�ˋ!�W�%W��0]0J����ѫ}W�o�H������)���j���i�̤\�^�g�˷"<-
z.mþ��!������R��АÍ T/f�m�H�bm:�s�gߵtI#W��<�xdۻ����FP!� ���1~lŘo�2�U�J�&��C���0�u���~g�t܁U+�Rˏ�UGv��E͈����L�%��;)�� ��1ih�0�:J��`ԡȧ�q�<Rݻ����*+XA�.�V�d@w���*\�r���F%k�e��$5L)#Y�	ֽ�2�m�L���ov��ZD��(�<�bĀ<���2 Л��x�h@�Ҿ��%�T����2��9�:u���*u�m��eRi	)���o����IW�@���&���)�����"`WI����M�9Y(~��������~_���`>ӕc4d�?�2t.��a���4=w
�n_���q=^�Ux��c���m�.����̑7��"��~���aB��Xd���K�z:�l@����S3w�t&k�jq[�-p�jD��D[Y7b���y�i�sc6g؂]��g;����9�!�ǚ	�s}-���C�4=�-������IQ9��9j�����Π;���?�#�cS٩�(�ҥn�e�Q���> �l�=��0ꋵn8% �����kfK��2Kb��� 7�����!_�C s{@�S�Y3���=����C�ʏ8�m)ʁP��j��7�5?D����*��qϼ��*:����'�X�moP�˺KxD1�T��]�u�-�0�e�ܹ����iX ���jZ���0ʣ�R�/� լ�-����=Rb�̃�\r���=N-�JVق!�ʮ���^GV��%�x�d�v�%��J���ц����B!a95��(�#O����1�#R�����n�f�u8��g��i�h߅{P�N
�T8J�y�R����}B�q��D�
�?�]��e9�Ry��5L�P�~��6��]r�`&q\���kG�@�>JPX9.����I�<��G���!�'�#j�g�\��2��^�����䭑�'��?�:y����$Y��6�6�(������6pF�x,j��5�k�ZuEm���ԭ�_T���M���Pu�G����� w�)��q��D��qj��F+��s�R�[z�\�&>̩s���G{]��c*(˴nH��~�����rЅC�+U#SFvV�rqUd��)%H�
�5�,\�ȃ�*�����+�����T�$�r����Җp����sͿ�f ��V ����D�徉�d>#̆s��S��DykMl�ƃ�7��~����g���Q���n���0F�r2�9b�`�k��'��>T���Dd�n��*8�xB�����(���3�e�����z(������4hN1���c0u>��Y���ެsO���Cݢ�L�h�#�*�������9�&�i���Ly}ZF��.�Z��w^e����oVx�@L$�ב�]v� V_)��f�_I���v��{���	��L.7(�h=+�>+줚s�2�{&+�%��ө�=z��p���/���i�ܜ�Q�� �~7��?UT�"���Ȫ3o�Ւ8�S����j��1*C��8�;:C���2�w)�S�bE�Ъ����!�x�5��#�V�Y��In�M���l�[eL��~<�kcR]�u;l���>�G�.�r�$�."���D��t�i]{�����B@C���W�_m���&���=��9KZ��"��Ѽ��,c\�"	Z�َ�K��T��� ��B(��UͶ��ښ�X�QP����U�|����<I��g��o�ml;�Uý}�|��� 6B�@���A�iu|��Aʥ#2�**�2�f��Y1AA����[T�F���!mB��ÔR�V�΀�D<ˮWv�X2�'��΁��~U��c�%g����n߭��N�����?P�W��|<�)2�kY��n�xe�~�w��]V�뭢6��s7�(+~G��H�Qɲ%84,R�6��E�w@H"i՚JȞ
��]��c�1.�UɌ�4� ��7<��X=�eI��?�E
Ah-�2ϖ��p�<MTG1��M�H��u�`ш�&dSy���U��`E��j�0��LN$5&�ca�
_r�*�@�0l�9�sĿ}@��KpFmE��7�h�z%�~�ȁ$)����cU�,d�4wc�4)�Jb���>������� "���m����\}��K�_T�	���K�SF�GP{aB���	��}_��y ��ʵk0���\j*c�q�}*0-
3�e���A4��;Φm�񕱲���L��ۯ����n��>a!8�~őN`~CE1R?p/���N�u���.��]���&�nR8��WUy�G�
֮6��2�"w,����Y?�VY��!�;F���	������F8���7����n^
3�I��4f������{O�~����Ïz��h�&��dysv�����9u�Fˏ4�=��FC�V̰�"�%�Tt��qr3oL���;�H��*˭��N�gZ���>'�+i�=q֨C������
f������dM�g��/��VG������聦��hY�c�а�_��{+�܌�H��u�ԣ�O�����l8Ű�o	�t�Og�7_��0��5C�8:��mb�k�bu�KWk��i�qb�XbB��L������u��3�/X���Ք��T�z%�ܐP�L��װ�� F��4�{��aKC|T=iC�M�㴹�'e�Ȕ/�};.�,���e�_)�v5�Mm�>�9^��naY�I�axkP,*���m�b���T(�n׵�@�V֙�+9�:��],.ɑ����EO֘��~���Ld�}��*���@WN��|�n�[�-
?�7ʳ�𪠪PZ�e��e$�kd&=��7��|�R���J:,���. ��ItT`�heZGg����2��4��ED�n�A'n[�*a���4G��V�_,`"|�X�?���GxЍ�Z���<����N�~�9����7O
�����y}�1���upe���>/�Z�c����	v��'�1��\�#��rg<�rF��/����9�S�<"��^"+/2ܜ�w�	�N� �٠�32��g�����Hq���O�h��9��z�z\6�Vڌ�	����"�S�8�r�K�X+��nB��˪S�WY͕}��|]�{����4:��ZY������"ӣ�_My�B�UD��|ϒ��M�=��qN�i3���%k�xI��wX��!`υ�e��Ҡ���9=��{)aB�P�{'������3���f�k$��1v)u��{�-]������@/���^S�f�$1|�v-�_b��JN�q�3��3|HX�;հ:m2s@�g��	�Qב����]����W�$��7�h���O���SӦ������IW�I^5�H�e���?�O��dIpz%Lw^	n��ik�2�D��8B)��BS�D�����2&��{`����F:�0t��Wʩ���y�J�ß��p���q���U��R��]��{�H�����KPl[I�pxxc�����0��H��(S�9A�ףK@O57��/f��1�-�� �gCVV5p�	9�`�f"��] 5�/P߉%�)$���Sz� ��ŲA�\����r�G�Y�}݈��|Z�m{�z��:a�����應Ld�QN/x�����i�*n�a�nb�_L	�2Ď0��<]]���ġ���f3�2I�8��~�R�$n1С���S�uJ_�T�+9L�׵�}�|��3���}��Yh\r�����D:���SK���z-���2gP�b]V5Gm`�&/Ngl�dE���i�f��l�n(>�H�ڴ>���S������2<O?������̛x�erNDT�<�Ne�H�t>�o�ٹ�X�it�C�5�Pa��7"Q��1�<�,�8��/�x���\q���?�n:��n�(�}!L�&�������o��+�ce*Z#� ?w��`�y�X@ǃ&R�|���`]�/@��!0Z�C�a%؛��U渽��S�n@��S�31�A�\�X�Fz_0ɸ�(��DP��PN����	bxD-ϘM��\�L��i�9.s��	���|�dY[sf��g��~s3��%��DLZ\Z��{����mzz/C�SW�������ߊ��k�\3!\bC�?�=C�J��J�d#:�0�h%�v�����6�6�պ�}{x '����H$u���ZY�C33�)����Y>�#����e�j#����'?p��ť�}�f�ar���y���>��k���g�m��12#p�*`z� ƌ��u�[T=Ydc��5=ʺ���s��瘆�a�>ɮe�;��L�-s��z�1�4��h��L[{����2��H���/b�K#w)↓,�`I�j�oZr�J��:̻Yd�YQ$ûD#��-�O'�vc�~9����U�č���°:ۈǘѸ�
����)H�u����~&|,���t芘��r<��S@�pH>��	��q8u'���X8N݈�|P��n���)����QGz����J�k؀g���$�w#Md~[����*��l�ܬ�Kt@�@>|�wK�p�-���Wa����࢒�e�%ْ����|7���|�5:>�ڒ�'(�~P�s���m��Dw�����4򚰓�L� �?��G�?�f�����hs`�z �{�w��� �/gQ<>A�s�/a�{��H.��'�;*vxw����N��=՜��F	c*�;�T��Z�#����#��I��&��t�Ҷ���6i8�@[��&]ƒtf��v99!U���l̆�&�'�����Yl��f���oC�f@J���V�QN�Kz���^I4JlN�B���1���c�f^���)��<��!�IŖ�_����5"�L�߱��u��"z6{�п;Dن`�9d�_�]J�=C�e������x3q-Tbk4��w��xm���\�&P|���ׯ�V��+��p�7#i�
1�:���)\�@o
o���j�0ɿ���x��]XO������e���C�����-�=�+��g����I>я������������q�Z�$�LĤ�b#m�w�ۺ���(��g�T�����o؄�Ę��B�����3�.�h4������0W�-A8ߵ��_�#a�
��?N!�|����߉���#)�9��c4�?�ue���+,���hhO�W<�<���F`�gS��O�բ���}���Gͬ��)x'6��u�+�%���th�H��a�A�Ig��s� k4���'gA�dw��;8@D�w���
ÑFҙyR\��s2�@̓J��^d��?��S�[�O(G,j�����'�� G�Fk�N�qj��c���?�գ�D��yr*Z{T����(��k��o�Z���do��IK^��s#eg8+a :LR�7�^׎Fz�U@���{�5i�T1�XAm��wH_�R�j��][4:�\(I6z��JM#�U3�@et
]��1z��8����u�PC¬׻6?aYT�t6��G����!Ŧ*�%������}���~c���m)�j��}�]ȳ���GC��QJ}ld~��TB�l��ˏ��@�g�K�)i*�=�a4㋠�g3@�p��XN�F����F��7�̠�$�e�⾗v_��Y��PG�3h\>#��_]rIJs@o �Do�R��=9o�3ސL$� (A���Fʎ�>�;�}	�i<�d�W�~zNIp魘bd��O�Q��6Ԛ"]���=�R� Z�<�e�"�0o����p�!5�$O!�O��6>>-[���n�E�Kk6����oWac�Cs��=�G�*u� ���0m@�詛O���+�M��$7���,�C��/,%}�Xp�f-3�E�Y7 qo�V��1�R�F��O��lE�=>ElB�t ��p5#�,�a/�]��`��3nh&�-2�"�ɘ�g3}C���G6'��D<��|�S&mQ|�F�]�$�'�L�*�<[>Oz��}-���jіN���fS;?}��IcZo�f�y+;�?I��`�e���0�/5ѿ�m<6���8�~*��7����	[*��ү�n�G�J����|C�3nxHXT�X#X�U��~o;�"
�.R�7�,P3�âi��Ŏ$t��_"�԰������9�jD�@��i_(��Vl
����wtI�,��=~�&���܈}? &N�=,����B'=��t!Q��U���o�w
�!�Ϝ�:s�{��b# �n�o
@k�U�8�U�|cՀ�&�c���K�׃�J�L����i3%?6�0��!��SV"��5|h�!s��N15�G�|ñ��i��M��$i��8�
�&��V�^&2,,��$R�ń�	r�֓��3�U��Ӣx����+��-Vp��t�&�<kO@�\<��X��S}7e��pVE'��Vm����;|PH��nG?�i�/���#�Cڞl;�����0-�E��^��6�)��q]uq��OÏy�@US��(ÜD���|�M��@a�3G��)<�b��t,��fc��]��F��k�<���-w���"�7[<�+��Bd��o���M\%��-������3�j�Ļ)<D��з(���3S�H4J���j�tB��$�k擅�:�}�����R�����L�}Ňa����<���Nەb�~����HߕX��r^�#ȶ��8L�E�y_�NDC�7���z�`o�|k���6PKvEh�j�PE���$�����HAt�	>N�'Q<�.�ǆ�d��U>̞��$d��W� [����)�Տ�}g���?蹫�K�y(D��D�O�$?�|#E�1����)�^[�eo�ef�,W뚿;r
z�dv_P���&�x�7��^�U���i�*p�ٕ U��-�cs�ế����
ЉŤ�q���8�2��Y��QhT������a�z'�['�����_�a�{���u	В����k�� �{1hN|�%|�k����`Oe(oD-��5|ӳT�H��yE���m[J�S��ek�f4���y%�����<b�����z;F����(���^���I�HoP
c�����_�Lg��^�>��'H49@����
��u�-q����L�ꄷ���:�t��D(���s ��?��q�wK�;�뺪F�{A>}�FD5զƨw��񱵃�HZ�v�R����2�WE
�L>&5��,x��c�Hwǃ96����V�D^SŠ�~.��_+�&�$l��1ǫ�6(Al&
�D{���'0[���_�BxbG���P���(��4�����GV��Keg҉�'F�@k������gD>���^���\���˫������j�燔�_����Y8�=��T��rcGuC��²"��ϩ��}����>��18��A�ɣ����z9����vl(C2A��-�,Ն����9�AY&�
�=W�	�����}����B�1)1i����,GԲ;�yF�x�sW�$6��·�p���H1.b��0�b����g6���Cn��e�iY���b���Jf	$D�5A��|.w���Ny�x��if/1��9�l�.ml��eFvY,�uj��h3gd"f7f�ͽ�����\%���|rW�J���P�0��lh,��&,VR��D�ܨr�9
�N�n�S��X�� ��,��]�Z���R�"�B@?��n	)���RT����<:��ƞz}<�\i��f� D�v�Jɛ��s���;mU3�ZDɚ5�I�(c�-a3�/��+ƌI�t�"����J�pͰ�y�N�]�Y0���\�:LW�W���VD���5�s-��o�y��`]��R KeIvрO 0�m�
�/�4��Q9n
'�8j�`VQF�eg�R
��
釙��E��d��V$���[���u�e�[0��o��b0��*�L�)�K��&z��.|	�|��f
����K������6��쪄�]�]����49Uf"[�r�'�p�������Sgc���-��cxWF2��.,��)������Bf�S���w:���L<��˗���L�m�IB4��`iL,~)����溙D��c=�<1�9�ɽ��P�:�8&�^z�N�����,ߩ�z|J@����2���q�fM��ܑ;-}y��5#�藱=���[^4(�)@m��G&�������8.�Gw�9rĀ�W�F���T�FFfn�e�����^\���Ϻ���#B�k]��,g�G�^�E�6����m�M	�]�HVџX\WD�N&@�$c�"R�}�-��ۑ�7Um)w읳]��<p�a���}��`g�'� ���)T��X*xy�k�#E�_����務m2�ۖH�7��N��É�b��;����e9gj�l��_ 9�E���\ӱE�x�h���!�:�X�D��l薼!`̫{��ŻXp��L9�Ӱ2
݁^�G5��r��Nx	��eLK@�r��?c����`��?;���"�^"p�{	vӶ��E 9Q\����_dB���8j�H馘���~fs�ݚ�����L���68�F�0���MFL�7Ix�Z*1nUW.[�qC5�`�;e&�I��!e��\�m۹ئ�������m	�6���z]G�kl���_�;���ކ��
���Nևy�׍���ē-NE�oƩ�?}%�[κ�U\Y����S`o��Ѿy�Lo��: [���-&	����Y����S�5C�ĵ�SWnT�/C�����T���W7^e���F3�Qwb�<M��(�Գ"k��E�A�[��'lUMMp.���M��w��VU���8C�
�c�^R��cv� �i�ɴ��>F;�����*ن���S����E���(=�x�\��N�	��Ll���n���Lm��i�u�O���FU��])�+����z�el*!@��x\��D֢����V]p�X
/��ߍ�:�L���/�\�o�1�����4ق�S �~N����2����\��m�w��Y�?�&O�r��~~�\��9,�W"G�UT�� 7Lʨ��s�#>�_$�5?��"
v�cUC��J��p���X����_�SI�}��I�G�9����촫{�ҝ^�i�Us jTe�}���p��D�U��AN,Vv�Ǖ��b��i�l8����_��
�h"�5+�q��	{*tD� ɑp_ە�͘[G���0RU��l*D�F�����g�[�L�D$��K�Bc��{����i��g�x���-� ȆV$��2����^\E��?f��DP#���?�v�zA��e����|�l���x#���ɨ_~<��h�7��)|�p�-��>Jb�o+�SP`�F�2]��/d��d�5�2L�|�!��/*-���R-���H�)�K!9�?hiȅ�.|Sd$z�7��4�	�8�n�9�e1Z3�f�1����?V���p庉
��[���x>o�m2]mڧh���_g=�\�O_�Ə��9<H�oWT���>e�\���fC���w�YH�<T ����n�=Gƀ:T�d�/�v}�W��D�\��9e3wx���#L	����r1:m~�j����@�z=�z�g�&������S�Ě��?̾r��1E�M9Jy��.i��u1ElW�'c{�4d����:+��lo��lUz]��4'��s��!����>}���K|d���S�8a2*Gw��Pٌw��f�N��?$�ِ]~����H�JEFȵr�?I$�����P�({�D�����sR�!<8���	 �|[% �g�F��h�u�0��Q�)��jDLD0Z�9�Gȩƕ������WsXX�٤A~֝�9��$۟�.���D�������(~�w�!��LF�Wk�7
Mb�I��,5X�ʝE��"'$j=���ŝ(���	���4z��c���ڡ��;��)��;�nU��>���+t
�ճp&Q����N�(.��A�W�&,����T��u$���N|`󳡷fބ�V�TN��I�ZO�|W�;E�"$�!���31	�k�f��Xoc��"r��6�u�),J��/�������*�?+� ��?((ҿ^Ւ�d�QۨYE�L)P���O�i@T�iݔ|I\p��ڟ���U0������֨����'��i����a*��V���eh=�9 ���_��tw2J�/�m�;�|
T �a�s����w��	����v���2���Ȋ�D�h� U���}����	��������,T��6�u�vxTE�R^mbdO�3U�5`������خ��O�� �Wm��Ń�"����	wSQ�B�;�y3���q>�n��c���:\}�s�#|����`��+Gj)��
�Ơi���0����䴤����
��
L��+(�H�@�P�Vy�a�����,����(�3r�(���E���.�wW��c��q��d�o+�]3�h�����^#�bg�.&Z�XXFΙTE��I3�Jwq���{���'Xpj[a�/0`�����j��s���64���1~�gp�O!���N���Kp��Iy�!ҫ�Q�!��BY��WO[�\"�jf�� @ߍ>t�C�P��6�E�����9�O��%�g�y������j�ʈ��?^����0�T��M�P�ʝ��.��a$!���	��΅{2�V�(��g�����JM�B��*R��ߤDK���W-�=������T5k9��	������&�i���F^�����zB_y�F)�L'�O��YI����u��ڥ�4G㰌d�ko� %�v��Z����ς����
����t1X�a!�BA���a�����}��2|��a�9y��sc6�v���:�d��ᡖ�\���0)d�v� VǷ��$a��2#�B���Ac�rn���8�J��|�s�,��'�D��,#�P�Vi?�$�5�S$8�͋�������E��̓�w��\��k��ܭ�L���:��'��r��,} )^���fM*Թ�r�����ML�o�DJ�9)�B�t�������:M8�v*��NO���E��c�UPf��ˤ�|$���JQ����&�.dk�RjԄ��#���3���Y��q�}��oK��^�tۘ�&c���n��z���n?,��0��h(^�aX�V��o���7<=�8".Vz�C�mO6.����'i��c�� �.��G<$$��u�(�D�ԙ���Ƞx�/0�TSc+˓��=!���c��>��(Q�p�I��x�gT��CX��@�<��=��AJ�*�1�¬Z�Ո�o����ߓ�0���0��Z ���'�&�gE>٪њ/�Da��Q7�*��ʱ�����;5��ڛZ'�c��8a�>�^��#Z���G��-x�A��Nzd�:�6��W?c��,4���a������b�+�5:�7��#���}���u�,0��s�X�F�_�Nɉ�ϹG���~��%���.�����%??[yZf����"x�KQ(Dڅ�'t�w:���D�F�5O��Q�n�mI:m/Ia�n>p?')���!�J�y�h��^vF�)�i�Z��Aϖ���{��Q�Mn�B��3.��RԤ-���'��B\�s�T�~���*U��l��U�+�1&��+_���RSa�������F?����(xqHj^�:�7�Q��l�-GsZ���Il�]g<OX��A>�@�]q���Q�h�	�Y|.�-�!�Z�;
o����0��c����,wU�_�I���Q�n��ԁ;��6�>�\�|�d�ys�at��u<��:�+ 6%��ejBEc��e�u���\n�c+PT�l�5�2ڛS�����ߍz���6s�~E���u8A�Sl䁨���9�19�����M���z�.��3-E�Jvɍ�+)h�n�^�R*?&+�%���4n��;q�Ө�z�J�z{����x�je\���d��M�}����'Ȩ���|��i�����s��%�,�F~�?~Je�N��y���E�RrI��Z��^����yе-;.���4��T�xEQX��tȝ-'�y^�m,oY̖u}���f�[)�mUm5���A5��u�5�&��O��M��v�} �
lP�W��;便�ʮ�vt��Z+�qMmy>g]��D���T�?!P�[���'=B�Csب`_	�K�s��Q�F�>q�Ʊ��y�Y���+�Qb���'RR��wtD ��UZ�ݎ�Y�ܧuk������c+�	ꡍ�H�v����:
by~�	��oI櫓#��~w,��˃����:��f��z,�Sb��#�.��^��`��Ɩؿ���ǻ ��`h��\�=�s+q��(;߄)�),�G��#ٍ���ɠO%�≔��6��ș>ƜS�rT`e��B���QhC���C����Bғdky�bLAj�2a��<!�xr�;& TP��I��� �]�� �x�ET߯��vd�ϝ\�=�i9*�z�ӱ!�_ϡ�m��ӿ�Ș�5��;�x���^-�F�J��E|�O�i�����i<���Cj����R��>�J��*Z"/�,O�FYn��Q,�~O@��0�O�w�^�7���:�j�m^��������ʌ����蚸�rMz�V�$c�c�XU<�	0e$�*-^����.+�����kAb�M�/�G�Rl���`U.��J��jAk������$�`�$�Q�'�s ��ↄ�	���� )?��,���d�r��ihS��ʼω��}'���z;:���A}܅�~X���u����"��yߵ�j��rz�.d���J"�ܞ���^�!��4�c	�&�^��i�7&�����c��h7�����J�m���:lE�Pvy�jI��s������ſ@Q��2@~:����:�%kMvGC8��Q�9.���J��!|U�@H�G&��=㽮ty�+}Hh��P�8�x�MB���vZ�1�[�H���j+�6��+��ޅ�P�6jTA�8�q*B���"}c��CՅ �f�(M���"Z+���R����p�E��#�Qw����#��OR~Q{[ G�#aP*t�$���l�/����פ��WZ��eA����e�O{��Ǹ������K���s�̥������DH+ ����NJ�7�|�rb4�i��x,� ��ΩZ��^����|ݵ��l��Veս7a��(�5R	c���r��$����j�/��en�v����t@p퍣IY鳢q=-=o�uT}�6
�.jn���o+��w*xΉể���, 3Á&���z�2�h�w�~��d� �Wd#]r�Au��V'R�C}�u�4T��Rk�0a04�ޣR�ɭ#K�=Ś���l�}�O��G�r��&�O҆��0�LJ��������7��u�;"�_��1���A:~'ē�n�ϙ�K���hV<���:��id�v��=�G��ñ��LBe����v��jM�Q�%ćw�Y:�]� �VG͓� r�wϗ+��߰���%������kQ$�k�At�T�5�맧^ ���L�U@�f�P���41Bˌsq�z���%� o�Y]�}%ΖpYc���V)˵�.���M3��y)�8�X��4�ƺ�F��B�k ��P`XA%��Y-}�O:�	�{�U�F�:j ,�i��Q�T��܍u��g�������΀�U�8����g����G����H(�^��هA����(I&��Np��[�i	��̮|rAHl������UJVmĺ��+2����* �M��=�]b���1���q*��x]�M[Ӌ �G�&qh���FF����m(�d\�Ʈ��*0.��? ��g�u���°��-လb�,�Qٻ����E��T����w�:��&�1�e^��ci �|0���h�;� �o�QI}��yl��[�7s�RI�IMD�c,H�J�$�-$����{V��հ�Q�
c�H�-^1����e��S3��),�$Vd%��I=���p�:$�jz&��Q�=,i=�4;���#���[�=���7ߜ/zQ���3�*>�^6�
�F��<ӇTs���dr������R�dz�DB�}�ࣷȲ�_r"�#�V�m?�����UȑX-��{cH>n���dL[��	��,��L�\�Q�H�y�%Om���wz�W�hZ���='u�F�߂��AR���z���?1ȼA�z䃙}���U�G�P�(�Y��%�+q�ݶ9��n:)e�<���!T0��E�׊9���2_N>�T�uE?�̡�<m���΋z\�n@��d�{$^�D���3b@ Gޟ�d�H�,� }��� L;-_Z��e�����pc�uy�޽�0�����0�W)�2�x	>�u^��O��̍t�*�i.e:^DD�J�"�O�5����D13v柟�]PLW�V$Kzrw>]@	#ETj&�+N�>���#.�)�+�:�e�e6~5.�%��ǇSfV;3�}Y��8��	`�������Wu�i�E�v�hC�u��O0�N����}h*_jA+�A@�Ka��
B��{���R4�g�w�'����|?��>��V��D�%��UK�E�+�������� P�)��:���˸6�Ī\XB����M����x����)�m�<?��X�VZ�	����wM�� �E��F�_�)_�_�v�cB��:��28�E�~��V��	Ã,1����t_�o��=�� f�.��?8��D9�*�S-���g*IW��-���F��ԛ�AP4Y�av=zݩ����-οf}K����hgp�N���(�k�P	W�:Z��u��`�u�P[vv��(�~��]ڲ����t���-����tb{�;ǁ	<}�bVG(����I��N���Q9�?$��+�pH8A[S�����q'#_�7ݍ`U���h�
�7�1H�4v,�Gs�C\[C�1�(��#'�����+�wW�&��0��`ZZ�?*�)�Q�{۫�#A;�����g[�?�@@/�//���:֚���Ovg關�u�k}�#��cvw��Xx�*�c����:TzQ�*���}G���6�d�@�`���wL���%
1?0�.��;.�%�{�����!ܱ��e�2Ny`� �� ^,"]|�4���BQ��X�lw��D�O��v�� �[���PN��?x�r�h�Ҏ�0BU��}
6��:��DW$W�̋;�
o�2~��[s3à�U��l>%\ �K���2�ظ"G����xsi"Rm�\k$b��&���+:�3
�yk�Ƃr4����J�A�|��X�!��	x�����4�
�Oa�R�A:���C���~a�h�DvГY�Ǹ�J�y��{��bۅ�@��L���~ܝ[1:�ך�i��e�d�[����^ݒ���2�j)F�
T��=��ϣ<_h�bF~=Qua� V���R���S{V���r�*)~��K���q\�<�>����p�D���8��U�lۑOѼ^C�F8lTrt4zp֖�##Z�;���wR*�/�X��"���D�-�v ߶E<Ԭ_�������J�a����p$�wa����3�&�7�kT�� ���󊯈#FU��D�^f�^BF$��7���eX�Ų���>�_�cquvaL� X�D��R�,�K���dsP�)\��!�u��`�שw�5��*�b�^�uJpG�C?�gؽ���Vbo�����N=�2�r�՟�SS��_Jé��(��W��u4dim��5$��)��/L33|�
�-Y1�⏉���k8U��uE�b^�S���4f+O�OmK��D��#���?��Z�btH4����������X;�%F��y6�S}����q�\	ܬ��un"ɽ�6�\��y�x����O����0���@m{��Ro�"䵧LW~�#(�l��c	��DJ&a�g��/�J#��ӈ!�����+���uݦ2���G��zY���['%��j�����S�Ɓ�L/�ݎ��i���qoaT*֓dF�� ��A܅}�G���4*QO�9���/�&��v����&	jّ�jkDD3��Gmp���|Y��v�쿔e��7�e6�{���p�%�-�AF�큅[Y��I�k�Q�0�����F����(��$�~渳���u��D�tiR&�a_Q��bKnA���>I����ӫLhVN�)��pg�ʡ>���7P��B�r
�x�/���i4�c���}��Aἣ�K]'�����E2�4�khܳ\j)��"���
4U1�Ծ�<��
�&*B߼������4�pz�Dlb+�]-4�3rJ!T>9��Ҝ��3��!C��2x7{��+odAZP6T��.dy455څ6,5`����Ǿ�5�J�k<����7Å�1%9���g@<$y���X*{��6I�r�B+�Ǡ	�����Ro�=r�L�x�UfR�i�^���+��<y2d�:����e��
���o��p����T��������V��~Lp��_�~�l]V�իkP�U�n� ��f!G3����"ah�̿��#mFw�0��Ui�P�]d�tWo�o�����_�,0�s�;ut �Y����a3N�*H����L�ʄ{�M�Ζ�]$���c{�]��H��2��G�g �N�B�>@��L�Q�ګ���4_a�z�F����^�H4�wI}?T���nj=)bh3�C�c4��C�"��j9�J�;^�K4jDK��v8nWk8�W��|PKd	ݠ�A���3d~�����V�HS$��M0M+0�%� $���F��ܓ08����-���ڣD.�11�6ݻN[��2P~O��j�Y����"t�G��	x�*�"H:Z�� 1��%�*���6޷8;/�5�H�Ś�ÎjcoCq����O<��-��}fj<�B�����TN;dl�}���q���3��5i>Y�/��*�CU� WC
f.�u��ߧB�(g#)���Ԁ~7i��e!J���(`$Q/�z��s�fQ/dwó��p0����<5�
Yo~3�u� ��)����8��@wB@�+*��A�=Y�*u�V��U����Гĺ>�o��V#�fh�Ywq��K��.�Ő�쵋r�;�q��J"����Ȅ�8
hˁ�������- s�܄\���BbƇkcq'Bcē�Uªj�t��J�)
A=\y����̤��܆A7e(��1�VKZ�
�z&�Xs��,��a�u~� ��7a�����d���U/[�k7V�֍��g�.k:��QSw;d������3�����d3���JLW�<*V �T���ٓ�_�	Clb�"4����ǝ0釳Xa*����;jw
������or ᪕n;)�8[��rZo��� �7�#���R"�`��U�>��{?�Ө���0qA����N�1��$��0�Q�/tBWx�����5u&8�NH�;����u�B� ��ԙ�����|�����Iظ �k�Z� 
^��<�H�%t��	'�����Nj��Yc�m_�5j;=c_��a�B<7f��v	�aV�w4�$ﵪL��U�I{��X%��y.x�:xJG���"[������s��_f����d6�o1Y�+��p��i��}k���F`����_Q���w=�G05%�%�����<u��v���F,��������n4���AT��#/\T�POf��(��8�N���ۅ�H�ސ���}ɒ�D\{���B�,0�1��ʖ�W�X���1-	f8B�XΨP�B�8�s��:waS�#CU�`r.:3Yr���:��h?Y���fx��M��
��5�'eb��r�`	I�L�
e����������)8L�V�	1�6�>I�O]{�Z#��$����=ʈ`]�Ė�O����3>������ng�1�M'����`����)�/��L�2�(��o�6�����--���_kWm<уv�s�:G?o���#)��|�AG@��%|.���Տ-�$�<Tÿ��39FRZ��c	5�j+�٩�ϣԃ�!� �����	-��r��;�p��y�7�ޮ����){A�d8{���d�0i�Q��^,�,Rtqo�A��Ju�&�4n������H�3��<�cepVG��7U��I�uOIJQ�1��>K��87B�*9��	J�'��̋Z�|�O��Q�B�k|ix"Q2Ϭ�M�r�H(!t��;=�ё�?F�HA�
4(.�������@_"p׀S2Y;�o]��Iv�_�+�;�����I�C�A�|�ܪ�n�!�B@G���%eZ��-�kjm ٜź{R�Bm�U��Ʋ>e9�jܔ&�rU-�Y^�����QL�E��m�m�n�l��nR�2�_a���dC�T]XB����EI�iy��t�Jb����uq�Ep��Aҕ(����v=Q������
��78]�t�ǺTc<!U��J.|��E�G��y��?ˎL��e��1�Q_fҙ�����X�!�Dʝt5�`��Ԩ�a5$�>+%��44N�;��o���E_��66A����'�y�#!�1}cS���F���8u��'wu>�{i?�N�С/�Eu�1����#����&v�8�T���}��w��+(�&KF7$��RVRK	�`�����ܐ�����r��-��d9�1��T��V~-�Ĭe��Ch�%`H���3�[z�uJUi=���� �ۀ��7� WV�N��s�b��[G��t+?#ab5-}g�vn�ݧ����=�ƧO���Y&ߜ&Mr%Ϻ�N\�<�|�~�6t�M������5�}�g&;s��͹�J��[�^62-D�o�Bq�c&���~�zg�j��~�+�/�.����� 䂘��U��Yd�&����pE{�FT}qʼDYBk��b��>2Ou���>Ok:n�>)�m���RJ����(�"�������ISS9+���~��.E"��*��̍K;N,�9ģ��]!���@zŘ��c�������/ؼ���ʷ�����om��K���X]��� ` ��_���������ɮ�O�\��4����]t>�.=F\6�O0�K�A�cN�n���S8Q�n
����t����[�_{���;�H��p�����&�������Х�X�+lи����O����b#�9n��P�}�����<��U�0t��ҙ6?i���R,�{;)�< !���l�P�<U�A`F\�bEM�v�����/z9�D��]����<	�8D�>��' ����}���4N�~|��%v �'�|y�`"H�Ϧ���e�K���[���4(_`_��z�Ӹ@i�H�ŎW���:<�*�C@t���7���qOaL�"��i$�'��ͨ��m��`����(;��f����I;xf)�� �?椽�ڪ<����N���[9L\C^�4�ޚ��TLSM��pW� z�א{����XT���em�����:�G�,�H�q�~�F#�`jd�m�W�@�%�l*1�����y���4v�č����7#�w.e�
E���a�:�8+*	�0ƥ+�*W��M�z�>n,#R�cM2����#);�.��%p�����~�ip�dgE����0��]�Z��&
�[�?���(�5��g2ݜ�yGa�pC�)�)�;xѐ�n.I�sۖ�x/�1�HG�4͛v��Bk�>ǎao36�w���5��nC�~%)2+�c	"�Rp~�h4���̻a1}�z�nf5�|�� J�:)տ����'�:�*�
0��N;?�!Ӷ�7��.����g�2{�@�z��FZC̏����	�"9"�m�~It0�p�$l���x {�vi���loP���9+����b�K�^���A��؏S�\ˋ�x�,So�ke�.�:&B��6�W,�q~;�Bȋ9�/K��!4��j�4V�6/�x:�ܹJ���L�jf(@t�j-�����t�>]r�XW��>�b.i�.�S�A����y06.Lj�P
ӫ�-f����l�:#iw9f�����
��=�
�sʝy:���_e�h �?�<EYz �۹�}����hcFP�B��#M]D�m�ɂ��5�a��6��{}��<�/�M�9�@f�颶�@��3�-��7�5��L&�R�f\�0SKq/z�P]:5��=x4��lé���!rE��蚔��.گ#t6��j�Vƍ :�4dJĐ]d�:g�=����MKOyzo����]!���**o���T�X��S.�	TJDl�֕≖Ӏ��M�}��{��J��(g�oi/�D�`�eJ���?��էs����F�+���E3����o���1��S�b�.�x:4R}<��2m���$29D��m�X͂l>�V~�0etJ%�ބ�D.���Dv�8`�����L�O�����\iZP��EV�[b�^��`� J�����ۑ�9�x�����5�YX�nb�>������F���͒.�T��Mt���z�[��h F�?�M��ziaz���|-�Ƹ؜oL�,��k�i�ا�I�eI����BR4Vq����z,=���M��a#n�눉�:e�b��Z]5�fJN��1;�Ԩ<iͅpC8�;q>z��H��_���ϐ�!�F� � å�wI��N�zv���^ �Q(e�� ޡ`l�a$�L��^�&�@�,/�^�FU�<�����
�n|�S��w࢝�{�6yr��S�?r,�#���LK�.�����0��A`NJ�Îd1K�<����m�F��v�����|�H��?l���	?���1v2���R��<23h	B���ښ��`V]���pn/U�����W;=\a��>N:>�:P�ǿ�*E���I�J����Ex5�s�:LH!�:�T�3���6&�
hm<_ȳ�Y�\ڠ��录w��<�<�ux�qojtN�a���$�n�BMߢ�,/( J�;�޼��M�٢bB���G�1e����u+��X����6�B�נw�/��XET����d��Kq�L����t^ �����J�R���F����y�#�J��|�o��G�)��9,��m�\i;��X����!�_x9.�E}<P��y��}��Ub�9İsA?�v���E���E���.��ů��g׹� �X�U0b�Z���6�$�����s8�����zw3��vLa�J"��;;rW�uN5\�J���ź�
���|�!����,����=�dm��G�o	V @�GG9iZ���;�q.�~�`������vb���E�d�"���!P�aX��62��x����5��2I���3�~P��5�n������bO��[��l��xz���M���9o��d$������G�,�ԖW�Ac`=�H�o�]����Vh3�|�r�A�4L��p��K�d��'ٽ����]�����T�G�
`�;�Su����������V�M�������U��Լ�� �\9�!�}�ڞ�4u�>$�з�/��p�C�����$��U3Խ1?�a���o��)����y`�@9��q��-��e^��:N�1���)<�Q$tQRX��>=�댑A�B�x�0aR��	w�n�'�@kr���>Q$�{�Eݎ��Y�|F}�^|�ʊ��IA� ��8�����+���#���%��O��l\De��I���#*��V��=3}p��˻�>��L��$�!_��ӆ�^�C���M
_��ů5}��3(-(��dڞ�,�������\lMeR��U8�/fJ�mn[8��~x���9��З�|��
����kL|���0n&��*�HfrX��e�p�(��W�<ˈ�2��(�i����
;j �xi#kz�I�R "�O�~� (yɚ�dU�n�R��n3�D�A�6(�-?3��k���9�n�Z�t ں���j��\8����̀%��Xb�8i�\�@�����в���H/��<)�Fv�c9k��0`b|�&7�@�$�s���֍���K8�Wb#�N#]b��?�������Ej(���O+?�B�nqל�MY��IF�0Niyxav��jJ��P�PYa�<�� �d����Բ���2`*|s�_�'|GU����T�_Atq]H�@h�F�� S5������C����ȷ��f_Ы�z;��Q"T�X:C1f�In�M��[�8�=Ze`w�4=W��d���c�t>�Wn$�U��uuI������&ö�Vw ��5�G��qը略Q���+���~�)��:k�#�Q���#��\�;����}B)v��T�N̖�xT���;�,w�X�#�n7cF����h?`j����sw����_�,��~���{7�M���"$�kMjgx6Z���R����2-��P�Hш0��u|U�*T�a�����w�#9��}ZJ���k2#��SH��U��5ֺ�+Օ Ϫ ���^�EL���p�8��3�}�"��:8������*k�m�n���-_��5Dჶd��`z�BAyMy��ϕ0�0<�l�E�Carw����
�(3`+ ?��pq;�LT�M@=S���-l�B��?�[>f3˘��OĘ�c)Qȟ>]+�����f���j�P�p��7s���bU���Z��}p����0DK9e�U�ʤ�
��ats����ɰ�F�vy:�D�Ŋ%���N�i����Hq%6S�E�/R1�+�<��o�<=�DN	���[�k�\y8�q=c��)R����X�.GE!�& |&+��|���'��e}�eo��v�U����KF�Vlܸ�Hg!��	�I�&��_�h����t���b�Ky�S0��n��J|�F�K�	#�h[�{�P�x�Ԧ&��a�"X|����<H�x]���H_�>�k.����/�E1�����ެ�hz��(p�>/ �y��l,���J(|kR�R����9Z��<(0�H�劣��2����W����Tq���	t� ������,N�,<=��L������Q��;��h� z8���y���έ7�R�"9�8d׫��Dj]�G[� W���
�'��Z�U�/��Xu~����pʩ/�C���IWR�'!���[�=6/�$�a.��}/�g!�v����t	�Baʾ���j޻�zB4�^�t��q��eȮXN)��~ʳ��L��/�/收j��SM���xJ0/�*L����H+.MW�>����5��r��Nr�+��`��4�����9[\��3}�^��Of�W���dV�	;D ���}GRj�/��y����4�+=�2K�.�sPG= Y��$�ǭvf�8���(�����Ȍ�H���ۖ�T������h��+����%}���l���$�����r�8}��Ԗ�M�:(ýq�X�e�9�5�CA��6!ʰ��]��(���%+7�O�����|(��ʙ��މe~%ع`j�:�˰-�b��g������uL25�}r9"����3�;�3���NT�p�S�1���m�zD�-[��2Cc=�$�Z൷���B����!nPo�7WU��=,#�1��
�V`����0�~����v�Ylp�^e3,�;�/��sv$���`��vR���]t��U�05���	�V����`�:�1Ӵg�z�ȽK����"������0��̪ϟ�{."�I���M��rtu��:N�E��\x�LK�����ɚ}Ԡm��YU����)�;�֖H\Y��q�z�x�rt��ʄ����6D�7n�L5�Twߎ������e���O���2	���M �����{��p6k}����sB�G�����Sb�!�0�,��ª�;���!?��2��([���k����"�ZM(�a��F�L"Q[�b��u8�!	ꐒ����h�4���L Wj���Qn�'�̙�h\Y�wW�	2#p\霢�ȉ�a�6�.�Qk0�[�ĉg0��ַ
����"�{_��Q�ΏK}���-ʪ���hG��X <W�Ϧ/E�;���"��]>���ςZ�_��q�߇S�~��6�ƀ�aّ�8�"e�Jҗ��J�6W�	�������;D@�vt~�io�\�AX��R!�d��=!|�Y�J(�2���wUQ[䥽��!e���(|R�^�4h�t�V�\[�̹�T��&c�8)�q�v�1��0����98>��<lx�⍥EOß�a[�/˶�豼��I�����7�4HE

67�'��=�e�1�BO�><xf�-�B���`�<�U��}�9���������V�~o��� �d�u~�l���Xx�b�@�R��!�D�&��m4t.�C�)s5q��3H���Ag��$�'Y�����q܇���APߧ�*O;2����Ś׫%l�P���f�8U>�4���j�e4�B|�cBDG'm�4)�%�v?M9KW�g����y�+NV�x#�F�� $��@�|��$:k���1�@_/#]��w�斥<K�Mӊ����ּ���|s��2�2m�Of��Jl�ė} �R6Q,:���`�R�v_M�F,�E!4�C(D+#=�p
�ǡ��}#��ET$_rq֦��rѩ4�t}}\��S��kWuj�Y�����$�N��{�>S��b���Ιc����;Ƅ�[v/w����߭fa����  H��bd�)J�V�Mu�hj.��Aq^�N*P?�7�|�=�d��P˘��^�i�t�Tc��0%��O�Z��� &�:D��������>R�c�4 3 ��c���5?�D���ay��]+z�衰x6`�����熍�ނ4�O��{��o�T�p�tj����V���z��[�!q�ic���ôЬM�͔qF��F�L��4��kDQ ��^^��3�����N�R�mRn��{n,x����\ڜ(�av<�������O���}�#�gs��f���Z2����l��=�ITl�����ӵq���#_�^8\�?:	��`-�ٔ�W���[�5-khᐼY�ϒ)��e�[���,&]W����H�䖍��.jhF�o�.ө���z����:���ۧ�ף��E���C>t��t}o=3��0�:M��ANT���6�lx� u��e��m9��'��r�}!��=�4���}��u���a�}��	�L&���r�Q$� %�<���hj0�-x_���$M:`f/�ѥ�y
]�6��וt�yik�[j�}�K�[�g|P�����36�OGCK����^@5��x麲�)�ڢ�a�S�(������"��6�#}f�w� ���EB�d1N���]���ی{�O�����i�d@�
�<^�x�+ߕ�}�T�M^��[�S��g�,0.� M��,�:<�sL��:z��@���ު��-�-������A�n�x�G��r�t��>��J����>�f�{�Xޗ��dg]w���%�-���>u�F�-��*4i�T�Ƀ_S��r�_�Υ��j>|g�����zU�>@)�_g��v5���Æ3�\aP����T|%��Ll���� `��i�-|�&�@�$U͗±F,�ɺ6��E��"��WeX�+C}aaʦ��-v�.�t�on�E�$[rd�̇߅��=N`9��R��} �N �V#� ��2O��Ɛ�E�׾v�ͤ؂�$s����ƌ'��w|�x*���D]������K-F,@�]����In��!hs���Ke
f'���,��YUm�t4;��t]�u���)i8?Ww_T�[I�����e�i	S?<�P+ s��r!Ai����ʧ��u�˓�]y�!�|��Ǖ1uw�I8�j�`N�-X�bE�7�۱G��V1�2=�ᆸ�s���_D�eiq4�6�9�w��dSÃ�B����y���L9��9!�B���j I�"�2�9���˿��ޘ"^e�^7$�*����'�=H�Ҹ㺺��]�E^���e�3��p�L#J��|��BJ캱����vD��D��`A�ť������X�3�1F)։B��4��h��w�w$�K���Q��`�	�W�%O'�e��xxj1�v�# 9N���X��>^�u��C�Y`�12
M�~Rl��h����W�a��ι^3zD���\�f��ŝg��Ц��t�Ͱ5���EM/�-�?�8/tXȿ�y������.�q֜l�Od�bz]G���.��<���)�'����j�N�ND �*O�|l��A���=���g��.���{C�P^�f�:V��1�AW�^�Ɉ���@��ŧ�cd$�+좀�@�Q6kX�g���Uɩ#��24C�/N.���ed$��$�[+¡�7a� �ؓ�{�̬mB#�^*Uyښ�k
��.��q;��4��q�L��tK�Dʁ ~�JL�3k���R�� �����	-����ήo�;h@�)�g�����H�SAA(V�Ŭ�A�0�?��wY����|���!w��,�|�l�l3!�*0�D�i����v�-���Ok��>��:�dy�4fDn1�R��3����Ty��}ς�ngI���B�Ff��ː�فG��ea�P��e�~���iT>ͅ�,��nd��fWJ�:H�b���E&����ƹ$�G��_�Ae�!��)�39%3 0��ض��m��VE+]�\I��uz%p�G����q��RQ9�uHOЃݥ���66�J���mb{��`��;���=�����	3N���6�@U�<�i=�w8��|`o��&�Ru빈YaA-�lQ���*KEƝWf)	��a ���3���@�\��!��$~˿C/�8�`��}v{MiS/F�6�m�NS�9bv_�:"P��E�&B\�ɼ�O�zC���j���Ug��[�"l^vL�v�r�i�VR���pKK��ͭ!+�����ɴ��b��r���,���@����$�:�j�ͣ2Ʌļ=o��c���pJ�H@t#�W�l�ɦLc�c���a~���[�vm^���
��!�B��6G#������I�Ѥ�;��2�w�w$���~�3�����X��j
'�5�*��z�{��I�:L�Y3�P�j`ET���2h��{`+>R�$c��L��C��_ե�l����i9�;�8[5o;�~�L�W\h36w���?\����{b�K�"���Ep_���b1(��ʸ^���:Z��Zw�kɱY%�H�1�d��O)a�$��a?yR�o���|㽍�����_3�#��D����r��,.����*���`����%����AQh)xp��L���Z�2���[�3kVŌfl�?�L�ޞ���X�oO2:�(!��=N��&�/ʄ���A߼��#[{+�/�w����hp��J<�۔8�_i�=4o��0����ep�v��o�o7n�AC��j�- :q�B����V��h���川 �H4.O�X�UM�tfJGa�������5��6�\��ԐG�e�M�ؠ�^���S��M9P�Q�;qҰ/?�r��t������I@��n�Q9��ҼU�E8lT�$Gx���Y����䰖�v�Z@�2���F�tƀbe#z�N8��<�G���q� d%�/�حmR��=2�UAH�����˴����I�Hv�&��p*{V�ѹ��F1�Hm�C�^�A�8�(ϿVg��[�[4��iMz9�-�V��t�_��j�\Kk	,e��%�c�F.������|�k�"c�����tՌ�HaZ�sE��v���D�;�1�>� �����%B$�o}���?�ĥʽ��C<%z��AK;��;©�F5���צ�'-�3%l�@���F�B���Z!�Lf�������ٞ��LÂ�c����*����f�8;�L����Tb�I}sT�p���n'A4$n4��"�db_]33�`%ݽ,{�8_n��ݾ]�����V����(;O�|���}�Z��^���yt�h���p͑��#0{Yu�at���aar4���'�W/�*Λ��|��2}L:�l�.Q�թi*�e�n!`z9�a��b:_���6���:.c�e��;{��pC?介_�w�Nقs��A��v�ÀUQ�y�!�F�ا&�j<Ѵ�_A��wM*���pO��n��,߷P%��_j@j/H:]b=�~{3�e�%�~�.n�4���P',Hx-��x���0*��z�q��62{�%򮫰�&;A��=,���Z0�f�k�U�h��㘾��Y1���y������T�W��t��v�vŹj1h���� R1P���Q�?�C�*�:�Yw�|E����z%�i��(���`5�&M�9�ٌ�1�O!�sw6b�^�e�F���ޤ�{w���6UHri�R���7�1���Z�ԛ�?�Y]/[��!��9I�� �+*k�>jS�,��E�b�jm�" �h�ir��*	Xj�g)��	&�ҍ���&%�����#�u{�U����|�gk)��%j�3���+-�Ģp`�c���KD�nn\Д�����;Tb�V'>�"{l���8�-��U��xD��B"aQ)�� ���=xۢ�X��/�`g�k��j��	4�¸�m.�{�L"֯��t=څd{�  R���z�`
Eh�^��!X����2�)�[D" 9d�BV�5�%c���s,!7���E����5Q~H�D�yY�tl$J��~����3�K.��N�,#�k���?���c�w	�-I���y��z���X
Ʌ�\���'Ec�t��@�����������rL�L e�a�P�����
Q�ry���E�o�";��z%���U����M?��t���J��f�Nd�r!�/�7ꍾ���X��k��93��"��{�	�"0�Sc��IO]��ghL�=dl�)������e->� �>���~x%+����h�l���ܥ�J �?����:�o����&��6jj�]IͭW֤�0���<�Q����;��w�D:��t�?�I�ǖ�o)�;sb��_"�5�ֈT��n<�Vg"��F	��7ѹ��n��c�}��,��@3��i�X,:fbә�
�ܯZ 汮ah�A�?�o�6�w���W�����t�O#���:�S�+ĥ
��J�	��BN���q��cߏ����)�а��J~���?�z���?���{�u��� 2a���O�m��>|��k��#r������c�����s.0$O�\P�D!��$�9��a1Nr�dךť�&�O��6fe���ŏ�j硙j*���W�nc� I��34��o��/���H����v���m���L�]�F���Q8j)n���oC���"�(��yA#����a��}b��Ah���CD�q��w������q#�f�kgi����Ao�c��w|S�|��8}+�J=��ϰP�����R�c%��_����V'�^��R��2A��]���^v�(:�����J>o�l����Ո�{�N?��_8�F����s��z�4�3J�1�JEw�A:��d�PwC�����f2��ؿ��Ͱ)@Vɂ�*����K���PK���݇z�(�V�YX��0�cˉͤ�d�rH�Mv�����fں�O�Y�r�� ��b��+큀��«ÍD6��v{]���֑����E{3FB41O�?w�b��z������/� z����Z���bpX����zK�{g?��x�9*��42��pӿ�'**#��&�)��Z��Ă�K���ܲՈɇ��fa��6��<�_��_���W���>�?��Qcp�z�FT7)lߧ!?NCLE�k��i7��%W�63�wȣ�FM@��h {P�0�6P�� $�t�ƚ�[�g'N��:"zq�� �/�@P��p`�K�YZrrHZ/T5<
��~�/�h��G�G3��=&H���['K�!�9]�x��zg���i��:_��%��8mZ��?g��s���wi���ǬC�[���w��w�9쫞�ߴ�^���m�ʿ�[�f��)�!W`39Z��T�����ʞ?��$�v׎eJZSsѧ����À�,x�6�3z0� Pu9-J�F7�q�����d���"Y=�/o��:�v;�~��2���'M��ڔ���S;�%Z>���I�.NV�\�, -)��� ޽X�[簒�����5t�\-;|`$n�/a�j1���n��,pP���(�vs�����_��[x�2H#S�l��*U����խ�<k�>�[6���ؗL/��8�C�,F4���
f�?��0@�/yP�W��(�/��c��z�{�}�/2�BǛ�B�nG���B�7�e0yM��6~���o�^�E@��r��.W�۵�����l���O�֋�6%v��@y"��r��4�XK]�
�e�7
��CD��{ֱ���a<���Qj]��$m��3�<�#� ɹ���Qi�C�Z�H�9Δ@�z�J煽�q�o~�l����Q�@��+$/��%GE��r�4�p�1@�
���ݡ�������2Z��8㨌�n����,� 3�\��;y�Kї��(����~�mT��:Q��|V�A�%��<H�Մ���Ԟ^���W3�PU��q���n�T�V$A�(GOE��y�u^A��Q���=޵���C�B1L� �1a��՛7e�f?1���kI�CaɖJ޷��n���u�K+�7P��ۺ�x� �8�V��һ�D��q;�#��k�0�s`�ߟz�I����f{Ĥm�j7��FA0���L��[B��$"��{����S zQ��o\]^,ɵ�Y��J�9V����EL�x��O�S�&J2�F����� '��$ҏq@�&ܟL��R-���vS�6(u�{��[�$y��5��
�%\p��̼�Xh���H�;{ĥ��<=��(��vb����\X��$3���-�}�W�d�;o0��]��]|#ŵF�	C�D�Q���K(��Q%�k"t]{j��Nd�#d���݄[���h�#���)d-�=w�Z�����&�T:���p�댶-7�S����@�v�T��D�/�ٰ�Z*�6S��(��9k"�ܶ�{�sD��(����7.�	<�EO��=C4w�����ړ"�L�?�^5�߶T\"?�y�ҔiI��t=�����hWo��H�?l���ac�9Y���h�x����h��"�������5�B���)��ib������'�[2���N�oR]�p��h;q͊�n����ိ�Xȋ��La�<碣�دHb�J�	d�˞�H��yn��su���߸���]#�����}�AR���|�+DS3�}ڼ���q1S� ��}G�և�$浙��Rm�S�!j#6��)��Ȅ��zQ��������� �����^Ji ��j�+і�ֈ���'����Y,b缋x۶)a`���,|A	5���`���Ж#�J�3�N�k�� Zj��ޖ����H�ᾲ��8��
���
��h�#�MD �w"_Y����]�xХt�I�%�~I��^�9��׋i��Rv<���H��ܰF���i�P{���2C��Yؐ�2�]��;��-�_>����L3��!�ԁT����O?E�X&y���_���'lVC�Y��Dc��~2kǠ |�C����"�.k\��G
�E��
R��el23�t�1S9mr]��˴�Y�a��#���r����J�?g�fmj8^�-U͙�C���������8��<�a��a�G|0������8�VrV[??e�:�z2�0�����/@�7_!��|��?��z����ZG:�H���v�.����{�ί�S�5V\���Z���ȏ�I �����B�T>+��A�p;LFfm�����qR����<r7��_�]��(��A�D��ր;%���u��3$pީ�9tz]ɼa�2`?ՙ`v�� �M3P��qs.���I�a9^�x1���$���jɭ^-�l:�6&�]Q>9�jz����cT��ZT�u�u��r��gE;���Q��W���������S��m��!�HK��} �yt\\�M&�e��`��Ϧܝ����My	6�G������4�Pc���Ͽ���-p~��Q����	-]FB ���j��<|n�c���� �`���qhj���z���Ax�=�<9���6�P��M �<׍�3�ƃ�2�Md���u~�c7[�ٗ�.D�J��>��x;�⠑`|@�ޱg#���(ҭ�E��EPv:�Z�Ҋ=�"����I�d��;��
�18�6V���
�vi�LJ��TkR�	iE���n�'�w���5�j1X5����*w����l	��K�2���&Q!��D%�,��l �:��Zm�y��Ω�	���Xȅ���b0-��ּ��E6E޳\o��l[��
>���S͔�N�z����+��,/v&���� c����p� ��#aↄ�K�c��|��W�A�tO��� P��[S Ɔ�m)���jG߸���n�q=���7�����br�e�q@֍3��^�^w��M\� :�$B!^�.,�<�ʷ:ļz�x{�*������/j�s�z�l/R��O�����.��5a�.X��S7��D<M�T ݥ3'N�y��y8�5��E.�?�ףZE��n��Pw?a�\	$-�$wh�I��q�D�	Հ8��k��AA$,����dg�k��z�ab��1�ɱG��[SÃ�ܨ���U��9�#"{��f�I����,�z$�)W�S��U�0&]�c��W"G��ʢ�V'�}�N*�D{��~W�Iv/Y�H�O���d (Q�\X��n*�MQÈ�+�@�Ls�����=|�Ra��;��?��l�}�*�BC�m`(!�$Ӈ'��@%@6��Z��ìG�z��yz'b5�w*���X88��ub���gϑ4�[K���0����۝�{ܲ��6�ñ��p+�W�/��6����{&Z&�F
�[ˮ�zd��� ��?tU���#��R�	h4n���/b��,6\ ?M+������꘣J]F�1��mԘ<�	!�c�����9Z Xm��1u���V�n�y�re�*�ߝf���0�BPi�c�F[f�F��®�f��.�;ߒ�GS�c��*�N��'+H�R�"�-2��ge-��nlr�0�}����kT�n�9plrH�&��
_�n!V�lO��qO�!�j�݋�z"�@�����.�,��(��X��[�����̶@���"j��,���]ؖ��ڰ�y'�ZpA�v�\m�H=<?��+]��.B�K�T��4�@��"�����B��m� "�Vp�C�.�E����
CBd��f���E��"�l ��柳~��V̒(k*�B��PS 7������Ţ��WV���Q��;	�"��+��E��Q';�Wq�Ɛ:��f�5��h��4nn�
��� ��V�].�q4�^���5ފhk�����
�ʡd�1$�����=���B�k��.�7�����kCi^�:��I�,R�~�m��ˈ[�a�Ӂy�q!���ӴDʠ���)0~�\�~�2�I���ӗ��G�C��Z�����,俊y.�3V��C�U��P�u�v� 8�j�i�����*Jo��T���ҟ�l<����B>=��Ee�x�I��	� T��N�4��M��l�G�vT��[���C��g�\bP���+�A�;�378��g7�|[aWi!r��O�ݧ7�����LY"�c��u�Y�u�(����ٵ�Fڻ��O;@+�6��,�6Q�9�Yo��/ZіQv|�Wj�i��il����ߛ��tQo��fJgŻ���c'j�&��w��O6�"�/10΁gD_c
�=�zW���+��s�2}X�J�}@�ރ\ۼL�_����g�(R?V�B(�7�á
-9g��;��B���,g������sf���K\o�-%������6����'�}���I�.�
H��?�r�2ʶ�#B�&��F���^�1�f"�Q<����'��G��52Z�X�T�՚����$O����Ӄ�T�S�c���F�K�c#��^4&cS�V-��;애ⰴ4DM����/�, �[���{�`^�4���݌!]Є�$o�U��gffk
�N�	y��t�l�t�im����R+�ӗ�f�W�_�e#�D(|RԱә�h�K���fG�n����KLH���	�G�.l�"���{�'�YG4�ǁf�G&j� 8����cm��&P˯��cGES������_�8���^���J�l�Y�\=6t�0�S���WwX裗��9M�
 �O�������8�5 ��w� Ag��W�E�X�7Իq��S�TJ!\�/��0�6�b�?'��q(򎩹60�o#W֒Y]1����ee�pI�6*��˞�����+��+�X�=�c+�[�G>���NK��SV
R�I����;Yq�x�Ty��%���B�(�	�jx@GT�A%WD�mL���w���e���F{�%0mI�acO6�q�A�:R#�W�Q;��3,8��AԆ�JnLJ����B�,��A��t�M��zO��N�� 8X���p��B��IL����) 0��
i�P�'���n9�Z�����'�NR枀��`��)//N>�͉:��ˠ�h3��p���c��q^�%��.�?����d���`chp�BȪ{����.�}~܃��=@@�!N�w��w4��RU`��� ���E�Nk�N�!A����9�X@�����P�P:1`��E��c��q�[BeA����i;������8����~B�jqޑ��u�i��q�J���R�F�\m�M���/Vĥw%u�>5	d�g�pS�WXdEW0��1�F�a}��ݿ�GpMmTI�L�W��P�Q<�_�Gl��F�L�0wɜ���K�A��m�QZ���CAF��
��?OS�S��(8]|��bw���F��!?#�2�(�X#s��A5W�(�'��k��
�w��Kg� �H�[Qp���'�x��;GZ�,�SZ�wi`n��������s����-eڕ h���v��sմ067Z7��
U(��]/��:%ScQ`��/���S�ELȱ?\[���f��5X��}�Ϟ��d�nb�W� 9MK�2��N����J��%���d���w_ꭸ�D�W��Y:,ݺ��h��>�p���ë��O��!>�Y٦����{���!iD^a�ą�G���E�����L�u�ֳ?��L�uL�w<����R,�E�wcPlt��y7'��;��mc�Z�(��Y펜�k"L�ؤ��BV�Jb��������4�06�Q{O<�y^8�A
^S��o���tVI6��3駐el���n��e�W\�?�Lm�~�@O�9jg�
�h��6;.q���w^�{J�d!ա���JW}C��k�$�k�opCB�M�e�k���WL򠰿gd�,e�*��[�CY�[j=����L�M�.��� ۾����6s�Г��"���k�n���cŬ�$�*n����@�T�1�o� 3������OZ��X`�g��jSh�`���A>���隐fu����B�@y�a-?��Ѹ"�}�-�O�ݍD0}���nYܦMi����M��)�[�e�E1�:j�>]Ŀd�(�dh�&5������Ŧ{h��lj�a3q��pgn�b,�=m���"ߠ�\eZ��	7����Jj�X��D�㼫���)��u�q�=�z2r�x�VJ��S���E/�@}J�uqg��So�i�F�<�|��5 J��#v`液�JG'�ُ��/.�'s��K�4!Gse��y����d�@꧱�NY���yG\6�~ѡ�5�I��"
�d�-��r_r���Eؼ$o_}l���W(��G��5]�b���7����ܗ���m�*!n%T��}r���cIt�p�T-��Q�]����<�y��-��p����Y�+��%/F��p5k^�问�rfg
g9�r�4r���Zv�p��˃�Dה�tV�)r����BL�τI/Scb:!JLW˟�h�;�^x�R�.T�+��W��"�`9�U�^<�ޠ��E�~DZ�[wu��|�qF։-�!��Ct����O���'�ND��)^�t	E�+��5�U|���qx1�7����}wQ/r9Zd�V1ԕ�g�u��}q�+��J����\+��~�N��Hh�A�i�e�&P,�R/ ��;�s�=�b1�9}s�x$����J>'��U����/jU][��*�Z|�Ya>G�	E损���#M���L
�`�*�һ�9в@�$�ZϮ�7�H���W��5Jb�-LE�x�^�hlv7@^� قLA>(7|f;#�9�C��nU'�$"���sH�(�vR+�����~lWH���_���ɓ�>���ڎ������T0��5�Ĵ�'�VR�4D��\27[�{p�X�0�J�B�� ���6��a���Ki~�(y,	yN��`C�P;�8����j�n�!���o\-���$�Qh�B�uu?]hY;$8|��~��րej�8-����s��: �m�b��w�6�f��q������f�iױUb׏�xi��@]f�h��[.f9�Ԛ�B�0��o�~Uq�!H�q�%C��6�8���)��0��Yo{ӓ�j��.�����[Qf��A����ϝ7P�+O�wjݹ-c��T�(=m�1��Қ^�A!]:�ػҜX�d2��T���vvNB��\b��Ǳ u��r����YW��]Q/]����G��4���uI��'�G����z�r��V ��y�t�*�J-�z���H��u/B��mx�N�G�d� =L��A�Xj)M}�lE���r��0�|:ա������P�YH45����k�\����E^:F)�JM�~�!*[i��v�O�%>Pfw*�X�F��+u$F�ە`���'�ܟ��G��M{!!ſ�Jr��L�������E�f+�Y��O	��Tl�]�r������Up�5�� P�]�<ޑ�F-�H�����&6�NV���"1C} �R]nA���vQl�N�SAΚ2�{/GZɞ�9$ w�8�T\V�B�L��s��VkA���{9�$+�R�}�� �"���a���Ѯf�Dwä��g'���0���hԂ�]`}��?a�M[�_���j
c��Ԋ��+�BrE2�#��tEB�dD @����qO�o���=�p5^{�t�Lg���}
2F�B�8�oɧ��7���Ph����w/�%X��p�AKau�a,DD�x H�T���}�t]��Z�A|��JJ��@j�e�R	ݳ<O��gz�;ې��a�7z�#"�(\�Y�9��n�1�VK^��*E<e�Y�G;�^z�̦:y$���,o'�*�C�vXa�)�R���\��PM�,�ؐ$�=�6n�|i�A�`��-h���m�Jїga��a���"4~ͱ>KU=���Ҫ5�/
�o?b�e����{��2��_��t@���(���@��q����,��<el��Z�h�,L��YTs!�9�_ �;ۉ�0�ֲ�y�<��@S��?�M�6�h�}p'����%(�m'�Ś2K��t
�q�����d^��Bx��@$���jO���["��2�jE�&�!Ԛ����� �-�K��A}����xH��$�X'����~�3� >��KI���P6Z[R�}zߺq��c�t&��!=�3ý�1�r�0�D7�ug`=O��k��Z��%�S�S�*�k�$������U<�ѐ�����@��pצj �8�G[d�����А3��<�W�1�n�iiO)h�֞@~R��ՈW
)�8�*+CU��������1ɚ�ͥJ%�ث��i�s������K����o�K�ފY�:�g�����}�yNu�W�`�B����s�]����p9�S�ۛ���@؁Ef���`n�SO�ٚ�ݘ��-����8��"��j1)�����������&�ۏ��g�|������ V��!E5��������j8�&(��I��i���Q�!C{O�G���84֡0KI/�Td��*.q��R����9� W��-�c����DLd����)��-w�K��_��$B*;�qv�O�&��ԁ��.�4�����]�u���u~��� �K��5��B�}6f��.�^��E�BGd\^U�
Gd�X�fh&�0,�y-��ArQ�OI��\���������jӣJ���./�t�C>#�	�(��`�J���f�$���A�h��e(Ԙ�i[Ƣx#��:(_�-��:t!���LD�w�v ������}�X=$@��q�ޑ2�f��p�(�q@�	�>�����nԡ�����qR�0����=��7;�
 �����abch�����%��4C߆,\¶�;Q<��K���d��+�W��:��W����������‬�bR�o.I��`d�j��O��-�ҕ{a"QW����2T` �K�0�P���xI�����KDH~�U�������*��eR�Qh��7�g3����E7L�(�j���&3AC���voR_�Q�����%�
ۭL�Q��#҄��Y;a"uN���M����	���9�e^	�����d=�hav	�sk𞰐�� a?r����1e���Yr\��Zs4+��^��ɱ�:��m�8�Y�{�i�֑�����_�$=�
��S�	�2 z��EA�x��i��z�E���Eos�� �� �����),(�-z<_5^4=/�%��{������� b����	\3T�-0�*W����C���"�:0�!x���(�R_���ޓ�L��.�āX�q��m�i��~a�*nO�?n�[Ru�}��L��Q"�5DF�'Z�׆��*чݟtY�y�z� 4���^�CNx�6X	Y�I�\J��a�"�A�H�. ll��/�LZC0h/Zf��f}�e���f�3��B�k���:���W�\�wH8�a�y&Y��Ͽ��!gU����x��%��9n�S���bRj{ (�1�)8y�7�n^�W��T|���ݯ�fnx�Xq��]��v����e�	������F�������t�$���ŋ���X6��a��Rl,B��:S�d��r�L}��d�ؑ�x_b{qt��SY:�J�>��Ă���/`ŽD2t�Ě�����"T:#��o�7|_Z�1"����N�L�?W��޳��.6(嬒=�O��q�I��Wi��V��|���3��;��F��b;���j�2����}�$���0�>��=g
G����ɌH�6�'V�_侜q�GI2��Hs�>�@���zl��G�D)�0!�B�WwA�.�-�R��G�?za۱�P�Ŀ�pHߐ���JX�o��=�ߎa�6/e����'>q�0�{{�'�N�)�-$�����W�^�������o��޷ ��^��=L�+�&��RR�տ��š��;��ک:�s��ӯ�i���)pX#}�A������B!B8	�c̶��]$�}Xf5ko��,!\U�E���wYDLm6&�9���X����l-8��u%Q뀱��Rj������y,R�&��#|
��ɶU�"@�a�JB�A�'�@�~/��?X��,=�q���X��	!1��p!�Ӷ���	Nn+�	�.�7+�	=1��RJ|�&�.�MW�aX����I�G�_��;�Wu�E)����!�[��koF�u��`^�b�?tuN�G����
���,hL�~Mv��gR!Q�x1���^�H�o;���OT|��7�ec����FP'���Մ�+��+�b�Q%X���_[�<���d�H�q5�a<�`�Rd�j��A�1��W$���bTQ��;�֚7��L����xZ� �tԇ;Mu��Ԭr�v�6��g����>p��H��X���H5��]���t��}R��-nuIk	�:���d&ZrE\�G1}~�S���;�f���?ԙ_��P�F�U6�a;7b$1�u*n��^�1��~���D�ZZ����},l���sw�Ŷ9%^rxpi��t�T�6���kN�Jp1A.0��hƊ�x�����H�� O���֓ǲ�t]�>��>/<�����D9�Y7�wݸ���V�s5w�Y�tcy�|~ř�T�(S?�� ��8L�m��bB[�=+a��(ɾ��P����H@�Iσ�V�2.~����ÝZ��v��2��ٻ�?���3&Mc{�8܌?{���8c�)��/ފ�2wRx�n!�#o��`�+���*:yo������g��\��+�(֗d����T�����k2X�W0)�����%(+L�q|"�+���i�_4eC}�������eS#��*O?��u���f�Ü�Y�|\�L<�,�ana���C��;��2{�O���9:�����қ䫠�+���4�Ί����mi��|gj!<����;L ��g[��$�I]��xI`�zD�h&�H*�4�� 0�!`hR��3���Z~*�{K�K	��"f��i�°�_�ڲP:�D&S#'�,;ู�}��e���[l��dCd�pa��&�8�dX&+��s5R���(�]M��7҃��x��蟳��L�x�O���b�U����j������e�2nN�}���>h�UeJ�����P��Aך&%�wn���B ���������X]�@KMh�� �T�T�[�N-q������U�=��2O��cO\T�(3{�p���4?jM ,+���
��j�u)ѷ�m&��2k�j�C{jd�%]�3�W5������+�B���9d��q�q\�R�qk���@l�g�pŝ5�q���b';z���������9��5�~r��|���q�D)��4������|�$����%=!������7�gy�@� LEG��o�/��/�Б�|fu�����V��� �������>�S��\]�(\����mF�`���x�e�L��(�}�	]%�@�<n�⨲�����B���>T�w�Z��h���g�2z���yo�ع�3
�}X����������H1Z�[ �1�_na3�]H����<�C���z��5�&~yW��y��f���
�cjOw"�k�UW�9��T͈Cj�=+)�`~b��lh�ƉN�<h���_t�@�G���� ���V�I��/T&:��������7�_X��p�v�~@p�C��O`�(�,���28�ze.�bU�ܼ8�:3�NᯅSd�I�Pup���F"Ià�~3���F��{��WނX���_�_��>4��A�iw�h#�,)�7��zXO�xIJ�) ���I��t0#g0��WW����Yڞ��W��ߒ3�
Q�D�ʷjO��Z�8���UaK1��?��9z�y�1\{/��gP�;�� M����3`��I���K��iT_�P�G��]=������ Q�01O2�F��-���Io籖�N�m�������̘�S��4XTշ��`!�#�b���n�
� ���gM��x�ݏY6���6���ʭ���ɉȥ=��bYY���:�r�<Ho '������>wT��h���ހ}�h)��3�*ֺD΍VC!}�����C��<x�Eq1D���T�1�ĥO�Jq(�P;��rr鼇�
?��}g�\�f�͎��,r�Ig/��Ѳ�"��E�x�^i�X]ާT�u��,��x���nx��Z=m0�ALk�C������4Ca!9޷����/�%�ˋR@���Gb����� 
�j��[��tw4�"��{��B]5�¤BK ���0�7]�7EK����AsĮ�d��lN|�(<ц�/���Ϗ���H?���g�>�*L��#8*��|ED�+:��i�M�<-P7a˂~M��t^����y�u�W�(N�mI�K�7��8�Z�h�?�E�?Bm�!4 r;��V=&�Wu�����u���^�@}�`'���/�#���Q[ڳU^�V��<0.�ۜűM�^�����P(��t��7�ȥ��+4�ʬ'$�����������}�J�;ҠF�¨N(�]u���"��Ć�������Q~)�>d⸼�G�>M-!�/0�4��C��f0:��F�	�k�u^���G��z�~^'VЙE͢k�i����'%��7_���W����:8���x��'
�c�%y� ��Ä`2�%�'}�!��؅����)��a�Ռ7���n��g�|P��A4W�4�@�#���t-�����J��6��6�������1��aG���2��ϸ--A�WKa��G�yR$V�T��i�5�Tќ�S�R7�t�S�X�r�p�/J�WH�^	;�d�HU���Ǜjp	݃�O�@K��-��'f���^� :���Y�}���ߵxS�..o�-��� 1Hyk��a��U<U���7������{�U}�%nG�6RYJ��tW�������m̆.y>�-�CH�E�˕o�,��>&#�j�T� ��*$9.����G�&)({��%!�Xя���@��<
��rq�ݷM���]�8�Oa�-�Γ�Ib��l�=RhQ��N&����k_Ι�6D��nKt�h���
�ryZ���j��m@��ٝ�)Փ ��RT�/��T�rǡ	����KP���?-
~�B]QIY�T��'p�v��ڔ�%��l�r��ɫ�y���#U+��۷@��B�vFzP�"��3��k#��y�Ao��v������J"�=�9d<Lk��mnʱ�G �2J�<l7�T��_S��}��.(<����ԓ#�9(%�d�NJ/>�U�B!��?�&� �A����N���:���ѽ�a��̗��F�3ᮙ���$lܟ[x�a� ��J�%���k̷�Q����L��`���a���F=[p����N(��|�c���m?ɿ!�k">/�Do�p�=+�*�щ�a!�S��U{��� VE�T7���X�+Z����0T
�S[3��U^JsZ�*�3�%$����i�`�f� b��mq�%�>�d�)�*�
��Z &�!L�Rtyµ�ɒЙ%uy��E��s���ec��[B�w��ѧ�o_���I�|>���Xl���~*QL�/�h�|����ͪ^^���
�_���|�U|/�,��p��M�ïР��\�ܮ���X!�1�� d e�����.���/�Gy�0�[*�1rb-@��&��b�$M�OX�t�I�\z]	�������k �}�����)��-�ĸ��~u��v%E��_���f7����x�2��ۣэ�Ȭ���@���~��Y-J������8@�`_y܀/�[~~�&����$����W�ͧuMppzY[U4$Ct��`*B�u��C�b�Y��[��!��0�����\J��):�����uL�'��K���n|�-���Ԓo$/�d��Ju$���EY�-첱�d�W��ש�T
PYSNRf�L#nR���i��cx�^R����ͬ�qj�D8�{+�J�h���<Ӛ�����Pb���M7����
1�\�j�f��s(�%�BCa�?�� P�ƉԤ�X*P��_c�밺u�Q� �e 3\��F?Rw@�B4�C��}2$���Z��MZV��.��{%��ǹ�%:D�������n2G��[���_���	��$^or��j �����3��P�$0x׻�>�������9�?1�9~h��3/�B"l&x����I�_E�p���r���<�Ȉ�
�>��ߞ�.���zl^�@�(���a����{VB�l�U���o*�A]V/�:%?��6��  �H}�����T\��0t��7-ٰ<�V�H�>җf{$�vd펶U�1z��mx)��b㦝�%���N��8� �}�vJ*������7�T`�X4���8���nmra��]ri7/� �Њq�xv�.vT�]dssJ��s�k�%�����v�~#n�GRBJ�*��l�m혾��0�2�a��y�˿�)��Z�_7�7��n�~%������^�I�XO��(l𗨥��ǀ>PAq$:�_�&�U���W"�u2V�yaF?�L&Se�(�K��^��ph���A�1V�]_�s��������YI@�?��>��2j\Hs,���
qjk/@��Q51�/�a1'��d� �Gz���z��D@g[�ۦF����+U�|�mLŠl����d'���t�^�7�r���J E(�ə��7})�Jۀo �e:,�D�\qP櫻�{��A.Z.j7��/�t�c�ƈ�T�91:��*d�h"ċ�W�p����~u��Y	L#�	&�| Wݎ�Έ���㿖> ���J�x�DJ�M�R5�)=eJy���J�/Á�i[�Tؖ*�>qc-K&��l��$@��]��W]->)�l���y��w��Y���� ���0��&��V������&`G�ؖ��ĳzl?:�R3��U�.�i�a��);���h�BroӘw�[>��_o;!2ܰ4>C�3{
�;3��\������q�֓e���Hu��h,E�v �ר �0t�g&z�R�M�
�_4�-h��/;�,m�ޓ~�
���n�Pt���`�M���/�Cg�_����Oe�f��sy�`�����}񙥵��?�u�BbĿ.���f��4��:�Q࿰���l�@��e��B��)���!��k�iFg��wE���S�w�֔�g릜��̶��\���G�Mv_լ�� w�!��Ƌ�lz�bVF�v)��5�	������֭C�|�L���H�	����\\�.8AS����ԉ���h�+삎	��ۜ��0��F��n�o�����dp�&ǚm�=/�'�C�o�䃓�0�x�J�����M��]�$��l���T��:��"P�5=g�2D:a�FՏ/�i�AbGR��r9�E��2�yIJ���c��˭|����"���jƟ@���Q��w��~ޕ恨�I����X�Ż��xto��w����H�O�Y�Vf$y07��,�W��)!<�@�����{>s��5���JRq=&�Ȯ O~�t7g���Hkh����U)�$�MSTZcgm1Ϗ�E8�0~n�p�ik��:�\H]G��8�C�9��`�7yPǝ���R�I�����U�%�����XTћ��we���?�wH�-$w8��R�#� T<��y׼E5M��O7.CE�������fBsLM�8����ٰ��O`R���3�_�=-j*[̨��̻���&����C�.r|�1 bD��Б�e,$pG`��Z�B5Ri�ޮ���pA���ԗ�r\L��<@����Va@���2e��X�j�Z�?B�~��R5�1N��s	O*eE3}��9�MJu7P��ě]�� ����P��W��Z�$�:x�-Z/���7/>��#�^�Ds������>Z u���6Oܞ��?�/���8�c!	���B8W�+���q8��>]����j�e)ղ����ཫ�!o��8�S�D�F�q�tEC�C�xA���'	�݊&nV<8�aX��8����Տ��
b�/���6e����9?A��+;���&_3���h���_c.�
T��������._Z�
��$*hS�������y�)�K S���T.�Dt����	O�W�����������Fj�ظ��e�D��A��fq������3H�G�����(/�����
�r��2�s%�:d�Đ��|R���!��8���6���E�$���#|��U��t(��2�G�ȋ��yH� �%8��FC��y~�w����}m��o�g���j!�w����T�G��6*�͡��ݓ�S:�2}AE�G����T[&=��TNl(=uu�|�#<�E\�Y����j�P�z�'Bo'pz_.H������2���).��Ȅ�h��0�k���)�e2]ӏQ�ں�۽V�W���ٚ�6�'E� ����M��ʁ�\6D�Ο��'D��	%�������E�o]j��G;��8�-5=?�@NH퍃�b0�P��	�P��L��H>`�U��u�W��������g�A`�[`rH�K����Ma�UJ�f�"
��?�(CV�!|�����Nl�I��i)
�hq�]$���Z����x�W��#FH��σa��s�og���@���Ef/���r�¥FL 
���yyR�Ʒ ��&�/ !���dg��j
o�"�A�Ҙ���=/֔����Bq$.�A�0�@G]`
m��f`�(Q�cK�?+�8]�M,�mD��E����L�r9�1�j"�����X(ցm2���ǖ��nD�}�{'��,��Osш~�z앮�J�Np��j�f�e����@&�jm������M���Y��^���V�/�;s�(�/��p�{#xJ�Jm5X��ȼ1���QƔ�9N��E+
��њ�P��i�/��X�
)7XGJ����6���7��#g���z����Z�t�S�<��3/����l=l@�۔`�~����.�ˌvHqs�/DPM�-D�u1G����LExܬ�MRGZ<��ۡ�v����<���͐e�j��W��MUD1�n�L�[��P�h�܌(]����[�~1�2 -VRK %d2y�]*���3��Ą�,Eַ3S;��'w���o)���3�W�,V���	&�.��L
@�B�9�C̳��`�,֝�����k���<��$P��%���a- �!L�KTסD�,��S���(T '$�$M�-ed�Q�-��Z9�?���9�C��2W/�e?}�]����D�	�v&�.�`�q ocNQ����i|�7�<�H�=�~��\T��5`�$���D�t�O�Z<���W�b�"�(>�e�����,�Q�Q
[��֍D#<�\	D����aL,���������@�l��T����yf#wc|��2�rV�,��L[jI�Ā������꒴�ܭJK`��1=ߓ��+!-�߷ݳWں�'�"Mʙ�.���ǒ�ÆgF��6�R�H7	J�\4e��聿h}��{�Y%����qLy�b|_���JgA�ݯ�iĜ���9�Ӗ���z���T�$�\U�1{�~����n8�tᮨ)3]U��*�	�3Q��5mNU�nO����>�ŭ�_u��U��kH�V�Ѿ������C��JveI�+��+&��8NnX�w�F	���<-V����VY�y��R���su��!�u�(t:N'�<ͩ/`\�.�o��i(XC|��o.yVI�<b�Yu�;�)UѢ뚸h4�C*��-P��"�Z{֌m6H�&_H�~����\/����ϸ�qш������N��c���y���=S"�~r�0���Ab�a���o�A!�cy�g�[t����_V5,Q���<�6��=�a�����n�����U��>LiQV_Qx���&hqs�!k���3�����X	)j�G)�,He4á^J�\<Ǿ���|ʪ�l`��$�炑2�zu���aB�����zՀ��;u�@�6{��΂�i9vt<@ٽ��U����cvx�q�> J­����W �d��Y*g�j)J'��1<�b���؇���v��BF)*�wJN,�	!�ف��t�;�@)�;g�w;۫����֛��g�U��[�b����W�ug��D���4yR�0�+)s�;8�.�������J;?�v+B�e�J,����+���P�D{��P��!@����C�,	Q��!�Ho.�a�����*�|�j83W  {�#�W��Wژ��������fJ�� �3n��V�����1�*'W5 �cW�(RDp7k!�[�]��}�Y�5��~p�i6�*¸�=�h�J�M��cO����:4?c���K�*���@9���%
\+��L�o�/_��6c���6ȋh|����q"���,l��q��|��*����^��c����ߥ���ʽ��kL���~��ʰDU�iE�����*��U��o��WAޒWM>�}w�r�J��
�knJk͝����>T5vyZ�����%�埀�*�:�����u��H-��꯼�:��!���`1Ӄ>O�}0��3��7�ǭo�ؘH�K��\��^�^b<9K%�XG9i�+�X �~�܀Y`RU+�]$��a6�Vh�%h{�l7���a���u�|�u���Ӣ ��G�g�;���9�;����>	aa!d���}!1�Ș���t.� uU3kR���?֥��b@N�P�9KH��Ƃ߶f�O�I�5�����9�J-��ׅ��Vy�S�q^j��j%?�F@�M'���%��	?���(�^wLB!?���'o��>���\���oPW���+Yp{2�Y�'�\K���x�T�Y�ۚZ85�j0�)�!�p�k�P��oS�!lnN� �&u�3ȣh�ͧ�k�EmJIC	��T�)E"�^���C��ßB�D+�5ċs~�sg���&c�,��
����=��G�+������ yBJD��a���[�F�O�Cg�Py7�Ka�򾩌ރ~@�;?�β���	6��EM^k��sk�æ∭�rx�e�ҡ����IT`=�����>�ey�/>g3�Q=;�X��I�5Қ��R�+hs�_N���z�0�3�?��^�?��э��8J=���@��Bcc�]�ӤA�·,1����;\��:��B2�����\i�_��^����(`j+9�7�}7���u��j2֎�1 �5���-�a��چB�M���HM��UvV��Q)鞛�R��4��2*iw~�<� ���)?��ZѺyl}i��[��CcAQy�К��z6B�坴�Y��@!(aJ���Ry�w��t}g�\Gb���V�=����� �%%�:����T�
��eɅ�f�f�1?�p�F��{�S�R6x�E�Gt�kI	��3嫲���3��1?ԤvgJv���jS�r��z�M{�'ҹ	�eY>���
�i�ET�u@�4/�Ѓ \S�/�����莘K~0v�^� y��(�{]�	�1;l�y�R#WU��4�;c'���D66�;���~Z���uV��L�p�L{u}��ݩ�Tݕ�p�EdnWMQj��=w�������=�U9|uWv�;'#�56��9Ӹۦ�
��
��(������.��5I+W=�����+�
��	CT	A��%����̹�0�l��W���ʵ�ޖ����B�,f�e���=��RgT�B�"3޴�`�l}Y��lv+k�܉8)���2�x�	*��O�A���P[���̃����!�5����!�᮷�r0�:I� �V����M4_�Or�����0:W!��^���h�|�a>Hm2'���e��DgYa~�>�B�qU.���<���� ��N�xɌ��GRY\j yh����߿q���L�%WF�i9�$l�����PZA�cc~��n�Wa�^�cE��N�UiA�H�ߎٻZ������"��s8�r��F ���/}�l�Jf��+m��!��}��:⚹��D
��<Z���>�Z� 56ڷ�X!�a��NԪ�>,zʨW60Bدٙ`��%^i0R��H=���p��_��ݰnW��Vv�Q��w�f;�+.`��@N��;��t�w��ᱰX|������S&����wX�[-&��Ά���Z�b��ߪWPJ p��~X��>YM�Z'W[�Q�?���R�1׌ϙE-��=o���o��4�qn�#�'N��qå'���x��.ꢇ�oI��n�6�flP�I:��T\�F�jlJO���Q���esH?�f�jV���7Q�XȎ |���:p����n�Ĩ��XPE�n٤�� �:#8�v��x��D�)-~	6d{����'O��w½�f�X�✍��A!��Nz��;�rA��Q������y�� c����l?ri`�VD��#�A�w5ܷ�V�`�Q�^ATܱ�Fs���P�ڮ0i[^����7��u8��	6&;�y��z=��u���1�?��J�z�9o�o�H�W~䕛���/곸^j ն۬#h��U�g�#u9��x�
3���CΔ2�xޤS�w��~��22���S"��ғMۨy(d�d8$�Jau����=9�C��߲耞�r2��-��*�7��~'6�� ���� +���R�%ژ�h �:Cf{P�)T�[���% ���4���^dZݤ�Tt8={8hI[����‑׾e��%a� +c�r�N�N�E�?��h�ƛ�EOb�T<o��ԣ)�ゔ-�����u���4�2��m���"|ب��G�)./F.z��s�C�o�Z&7<��_H-�J�$JȬ�:��<׬���U �2��Z���/�5li�M����US���5'W�q��T�$�%�XA�6���ww���nE0�f��~M�o�T��r�<σ���Ml_�6d��ܫ���l.g�/I�G�!D0l�Υx���Bc���}pȍ-Zϓ�9zsL�`�z���k0=q�aߵ�!@h�:��x���������(�����xP�S��؄ذ��)A:]uN�|]c������g�Dxá���ާFJ%�}F���_)�45�������=|����+�4�zE�M�]��9�4r��K~�	6F�h
VoL��s�7a���;+�(#�d97"�)�q�D�.�7(����o.�څ�;�0�)E�C�1=��h�t�H�8aÕ-�>YFK�������Q9E�z�gFx�Dea>a6�����XB�&ϑ�M�)�-�B:��+4�-�_+\*�/.�q�����=��uIF4��Y�AjZ�+`�J��d�̀���`�Qz���� ���%������HMB�ՙ��!Q�3��d_��֫�Z�Ju���U>V���$S���b�/.DYw�������RcD���̪ji a���|���T"(!ݏRn�+���w���kg���o���$z5w�/F���1Z�h�Kx��u�t&�"�����Y �-2��֎YN��U�f���)>&u_�@e0�D �wII/�p� ��RF���n
e'Y��\��\E���RF��!�%�۴v���r�RBG���Sl9�F	+�fo��IN��s��<�&\Ǵ�N��(.Z�9�g �> ��=�[�0��Ձ�͸3b���X�k��4���(B��N�MG".����(�������YH1`��X���ra<�; �
 �y.��z��l:�[����V��]��I��1\��.��Ɔ��ϸ�j�����k0)�?�&VT�"����񣗸���u�9AZ�S"������Q����e\�9��-��������ܨ�W��[}�a��#{ë�9F32�f�b
L����x7Ԏ��6&ǐ
����Hعj�E��(� E�׌9�0M'(%��	Ua���4v�K(�1ʤ:���'g�-��b���o����/�������\6-�ti�K���d���M`�.=,9�dw#������6��D�I�j+λ�Z��q�C�1m��p����eX�,Cf;�rl��9����D���̬�,���M^b�u4����w\༶i<��h��D�Q��l�|&H�xt��Z�q`�7��(�}kD�����?L��з8��V9I����=����lc��c=>'&K&��%���_������Hg'n+���9��΍w^���&ҺP����5R�����v�Z7d3���σ�7�g��v�X\��%�iږ�ސQ *��-�DڦJ{�g���^9���z1�3z�n���x�ߪ�P
O�7;�p@�.�!�<�Om�_Y>�<�%CE�������'�yd�1�;@w��ȥ߈��a	WP��F�L�@b��@ͧ�'W�;��ob��Q�P��c`�4�A�q��05�@�P�_R�(t�������P �gV��Ahpl��`Nr���"
��`پ�5��9Fs�dY��M���N���{��E����l-#��z�Y�e�!B7@ ��Oð�A������S�!C	�G���ִhA����vt��V�nu�NO���D�[ RڛD>{�V��=-�����c4*Uށ�
2e�R0EFr�!���Mp����5��;>�}ள/���퍦���U���zp������Mx�w@<Gc�N��T�0D�dp���3U�d���K������_k��Y����b>��f�.��=�,��1�j(Jf�>O	�<*5��Mh�y�qg8�1;<�@��N����^��~�+p{4�|�t��!z�����$�E�έ������!Zτ�~��	�;�)���T�X'I���arm)�	�A��F��������Kz��Q�Fx�5�h�秕����gzUr�.����F!9�}F�I
/��O@&���1�d(#�YR+�������Wy��a>
��|/U�y��@W�lx7���GÂ��/zH��V���(<4^�(�c�4��_�@�93�-�CWp��Y�B���̊�P�qU�=2���=�X
��+	��n����^(G[���	�x퉎q����т�^f��,ʉ��j�R׽�<ܑ�B�5�<M�8D.�
j�&����{X~C�T�v34$m1ܵ�bWJf4r�Щ j��#�����	6�X��V
����;�Df� ��[h�:��C�7�:=�5���,��^��>��;s���5��(�V���s=��+Wb�@<�B��&jI,kT���3���:��˚fE��X������g+�?^�:Z9=��� lW�Ћu�x:��iu#x&�߼�g����M���l��[o����g����/7(��R�%��g<�y+��pGa��CDC���[��@��U��������� ��!��*���-y'ʬN���`�CZ�
� q�jI^�k��>Gn��_��7/i�h�x��)���jS�R/�=��\�R����&�B�BaM�dn�������G�gX��$W�V!_>�Ű"R�c%5��� �k��Q�b���B�O�?�0}��R^候�BP(4@O����m��ݝ�]��V�Q0s�\i����;'���v�ӌU}4Tqg_�pR��wiys�� '8�ǆ��.HH��k&�Vc�g^�-*ة`2 ?|�.��A z�Eq����^��ԏ	Nb`Aq�\Hh�11/�|B#OK�^�z���߯�Wt)yQE� �qi�O�=D��:3�ރ�����V	<l��m�Y>�N}^h����n���_*a�3�$<��,��o��2�*p�_:=
t��1�	=]��c�P�^D��[����$m?�%U�˻
vp��Pa
��`�3���#I��'�m�kr��;���u�<���:���x,�g^�Z"0];R_m�͌]�����}!��-��C�^���Ա���j�:�o�]�h��X�u�w�IG ��:�`��B�2�0�b퍾[���	��	��<��G��ņ�]֟y���%K�CD�/Jj�%�!��cl�z��JeI���3�:P����歯V�U2S���{�bh��k�ą�>�|΁y)�1�X��6��ni��X(����*m�����׸����	F��J�@�)�i���~Ȩ,&:cldO����ܧn9-�#4	dibv���7�ԏ^A^��2�~�:)˾��}Yo��'W�<hr�d�.ڔO�v�#�l��0kG*�|�]N�ܭ×?�j�+H�"a4��ڹ�gfB��a�}H��<jv���N�Z\3�E�J��e�E�����m=��S�<�?S�����0��E�̫�h�X�����*����0
b"��^U�������(w��~a)���m4BG�%�y�h"��(�Y��w��|3��qe�@BU
��V��7҉�^���b3��%A�[�j�<�a�_�H�]P0UbD!T|���D��n͝2Ϡ� #
��/�+�4����7�N���om"��5�S�
Y%��5W������"�{�+ j�"��p��ױO�7����S��,��;�G-b1��q��t�����u�u�iK�ѕ�M�"�����/�c:�&��{�be$6��!`ǵ=�s�A�FYSި��/{�{��(G��{ �E�u
��".�r�%��F�6*[KQ=jd;�(�=�@� T�c0:؇WȄ�F�����`q�f�t��~�Fe��� ��e6�Ȋg ^+���xk1 �ogm|��Ю���8����a�N�(X>Y��ꯩ��Z��)�����7����J�%��.��\n+Ry ���p�P����v'���>L���B��Z/{:���M����`��(G��z�'i��ohpɊ�5�&�"�P$�&I��<�^��/�����ۤ]eJ�7ᑃlM��~Ƞ�$+��H������>��D&��y�� l�2e#|!�ֿUg�C����f����*Q��1k,��d�-Ⱦ����ˑg滂��f�
���kO�F�lD�X�!�l�J��GGw��;4l�=?I�W�v=�=Ab޽�~=�������vdq<m�rU�\�X��(77�G����4Ω��ݾ�o��e<��<8��
���Ά6}:d�T���T�ȤP��@!٧R`������$;�����zI4tI��XW"Œv�kN�L�Ҕ����[u�:MQ��{PLT��A�������\�T�O.r�d7�6���bV�iX�mf<֕�e`�6:l��_�2J�ȋAb�]3�L�v�쫎3Gu=B�]��\�Wix
�����ٮԒ�z�a]�"�C���㣕�UL77��������9��pb��, ט�Ģ���`~{����Ȥ����1enNZ��ʂ��E2I� e�!�\vs��%ހ�4ŝ�����I,y#�3Da�&��&f�%����QXQ�Ś@V�C,�Q����t���[yE��6Q�"����Y ��,�`+�\���4zY���Cڀ����_�O��+ �kr�&��]ܰp0�����ER��ڮ'0!V��]co�O�5Zu!��X�H&WRkz��Ur�W.>V�CJnj� �r/�*�𺷈��nsE�Ɍ1)�
��oj�^��ɯ��7�1Q���'�}�Z�jp� ߢ���y�h�GZt��_�&�'>j(�b�'���1|�R�5�:���-y�:"r��^|������XC�A:��i X�����^Pr���t�R��O�{E	p����[������<�fYO���=����a�Lp��w�f�E'�e��\Lw�Q��-�Ş27W>u3� �ǵp��A�?`�J�W|k�� �E�>:�[��z�By�}-#�]�1˻D��+��%&�pãVKp�@��N6����3��^�b����t^�TҲ;��.ҡD�j��67oe�U>P��|ߤ���A-�s��Xx�2c�����y���;�* �/=���8X��}ހcQ��D�E�X[�*�������.�˒}�j72���z��F=�;�I=f�R/v�$�2�أ̈́�VF�����\x.��Swp�{�5)���2?K"ݷ��ZM�-E){�WB�$�]s�
�&��BUg�gv�[�2 R����Ϟ�'�ֲ-~��{QΌ1�Kᆈ�]�/w��G���u'�'�♤4e{E�gy�����2+U�W^�F���&�i�}����s�Ŏ0V���l�0��!J�i<R���il"�wMqW����8�i��"`�f���=����!?�g�-&HB16�8�n�Q�n�D�.�#|D�ayN�x\�F�m��;veC<���oZ$����\��J��������/�^w�ײ�qv6�Mz���O�xt����0p��O�-K�?������tZ�nI������+;�"퇂`8��20��E.2�])��7�����'&��ww��;3��S���f!b�GE���`ĺ� c-2��5�k�L,��(da:�ٕ\�����9|L𑟉m1�7��n��P��[��-F*�=EݵXD4�$���fe�3��\9� *N���iwڰ�(�����*d*O���/��E��inQ˧!�ffp���MkF��u��!2ح��>���Ǉ��`�b����(�ٟ����+�<��O�b�z,2��Dޝyd���ů�+�C~�~,�&/���m	��rj�P�WT>�H�+:���e��ⴔ�g��=}Kf� �<�x#Bn�ii�:���]i�{�b��8>�;�V����7��?��@�.�� �O�F��{O��2!��q�7�v���V�(��N��i>7a�Z�y���o��v|�gp�mh��~��@ݾ_'8�~��	Z�i�.W������.�EI�Y�!�����I���L�\�,�2���	=4���{)K��$��D�Â5�_Ô�|{�	���.w@�	x��������Z�Б�cD�;,��E"��ss+Uq|6g\���ѡ���@���R ,=*�K �����{.�T)�U��܁���N��ʩP5���LHR��+�I�,�o��bE��b���+�i��m@�c��E�|b�	u�x��AӀ=��Ά�텘���Č���cm�x���
���rc�W���4y��h�����_��k�`^�M�!/��j��'���ʦ�E���j9E/\)^P��u�#�/f�#����}2+�n�QQ�"~yJ=�7����%[�v���8W�z�]	Io�9
n;D���g`����9ʫ���N�ϴ.���;��R�5��;���*��ua��ԇ���hW�r��?:��\�����Qo6͢)Sze�A{�"�k�Լ��ux.v~~j�8������K���[���n�����h��$�P�*����V�}$�^%@u#�V���-Ԗl�ʱb��~X��^m����3�:���i�B�$��x���ўLr�\6���}*��#�̑�XB8sǺZ��<��c�\�e��9F��z���Yw�5�nO�:#oz�w���8�t��ˮ'+�M���Y3�2uUGx��w�<nbݓ��̒����k�K����|4og��x��1�Y����P�f;KX�[ߝ��l�NA��7�i�����{�5 `�;��Y#�I��j�������Iٺ>�D��`��J7^Y7,�vYz�	j[��[�fS�;p�v1���s�d(p�a,}V����N���ݻ�n�!7�9�Y,k�Wfr>�up��j
U_�w�Vc��1�{Y�F�����,��S6�Ixuu��zɑg�l�t��Ko���i'��/{n&�{И��7��}g��e��?�~�;����*� p��a�lT��3��ׂ�aRJ�|��A�m:��Ʈ�%����ώ���/����3ʬq�}�[Z+n��hM�m�]���d|=�'�f���%q��_k#ԔʳZ����a���8����q=ֽL"*�� *U���mYU\Y|3h_�m���H��|ԏ�"�S k� ��ӳ������c�<eho<[�H0i.�W=��:F��ҊR�5	����-�@�c�B0L2��2�C��D�J2>�p�N�9���zM�p�_X��E�~8LX��nz�WG�-]�y�F�-	��T������heI�!���uddkM��WL,��`F}��h�����W��Ϻ�ӡ�X�<�N�S�iojWkY��BN:M�h�:�vd��O� +�v��_��[abM��z�6��� �"#����l���f ���Sdу.�-m
YH]g�ZQ�)І�(�ZF�1�d�)���׃LIc�GG#��r�\�� Uv����uH�fQ�r�;��,gZAV咚�y�*v߃O�C�mƶ�R�8�o��^�b[�N����<*\�3w,/]�J��G	��y��6��>��QFo��-��.a.��4�1��{��
!��˧n�z;�����p<q��o�ZP����o�J�?�N9�7e�~���-U0��y�:��,R=MO�,�=� �7 t)�n0�іz���w�(�
�^�>�q��zu�]O�:���Y�.�Q_�c�?��%�D��>�/�)�7���R�D�l?i��dpG���x�г����0�<�1��x�T�^'^F%>�6�5|J�qez��*��t����lO�w��~.pŜ#)�G�bd�(쐣�QQ�k�gP��������{d�|�H��6XI��ڰu�,j���,�&i�'U b���oc����B`_�#1ǆ��߇�����?�Հ�?�W�E4Va���Z}�\�7��'�Gv�xX\{��?h�� _��X�O���X� �~L�F��L���zm=�:�[�gg��BXT�Z�U0�����/�Q��j`- �V���J��o�32���&DV{�$�/��]�?�I���׈�ᶁ1/u`c�<���O휻�ծ��~�"������T�u�b<kTvnRUlS�:��eI�OLq�Ʊu���v��#ߘR��Z��ps�)��[I��@�����L�-�(<��?�J>�FU�;�6ʵ�(�4���[h�@?�uw�	�S�䉖BA��Q80��3zIݩ��-cޤ��zn��l��߀V+qO�B����*�u����/��@���I/*g��G�+�꼁�=H6����u���
" a��eޭ�c@,b��N�7��8V|RQ�ް�"-(B�s��-[:j[r�^��ZD�ϟ� )���N #�?�����Z����H�B
���e�������6�a��o-���}�։"����2�[PaYͦ�3�%װNf�{������˺�u���]�r5&����A!ߗE	fL�L8�khiF;o��tO%��w��o�8�F����f�G�=����W/�?�<R��qViPI0��:�ʁ�����2*��^�A���"g�)�����Ũ!����C��Z�B�DC�ߘuN�#y�����@�4��ֿՠ(�<��|P�WE�N�5�@�7�����X�f�`�;�"�r���L߄��DD�^��ZZC�m4ޤZ�&�iJę )1��n�J��e�oC.����ly|3��J�A�\���/�h���g�g��	�w�(t	W�
M�I u��Su��������x�΢V~g�!��+Ap�@(��`�9>�nq"wPf4ň��/�{Ɠ�s����?)MJs���O&ר��������č�$�p�>��~X���=��E˂s�u�3���L"�V��.�>��i�K���_uM�C����u8~-���4"���aI8T\�� ���Y���M?���7ydya��bך�/f��N"]�5#&&�$9p��H�8"��[l37
�g��Z�+�Q�|����CA���k��c~E��&�).?ӗ�t��	�p�? ��[�� (�+!�]��$=��V�U��<��<�*���;�!O����L���y��X&��p+s���?�)���I?X��u.9\���24��
>r5�A�X+��CERv��[�6̵��+1��:#���ߊ�h �.���!TR-w�g��2�'���:�#�r�+IY(�J�����8�{i�=2����b��!��$z�͇y�yGlcl�OV2qŏ$q����|�Q[_]�_
�3L�0���k�i�i[��T�w��\�cS��R��i���u��"{J+�Y��q����4G���w�j�s94J}�dc��ݻ�qګ;�D�\�?_��S�(�Ol\�x��1cFG�IjR�3��ZW�U����D��5ƯȽ��kӁ"oy�+%���P�)����iٗހ�����\����tM,`7yU2u�%����7�}xQ�Ǘ�������q��츀bDRyƄ��9X)^�XB�ȱ��S+���Y,����_���1=�|����*Q�y#d\�F��֭'�Z�6U��:����c �����:�P���c�;S��F &y�^Y��o{���)P�Q ����� zL��zb�K�V{�����k�LP�������BE��5J
�f�6��O}�g�|��j�p�W��}�m$�����l梟T	��a
�	K�-�q0nѴ���^������h���i�-vY�b��D��~�F;�Y��n��^���I#�MfVf� �7O6��s�;�A|3��|����|I�FW�d��kB(:��M!�i~0LK�K���X4�ONˇ�>\�P��zd��⒜����%E �t�)ΜG�ʙA8�9S�u�/���bDquNܞY�R�F&���ʗ�K=c�5��otV��J�c��.�Ϳ��XK�YCN�q�/u'3�3�z����u?n?��
)ݯg���������|�"�E�D��Bw��()�q��p�׮+F�S,����FR?����^&Uz�y_F�OR�pJ��2�l	�ʧ�0ަ������85��� �\Ħ���P�OZ�3���_�o��q|��I���	O��v�ޑ�G����k@4�:��|$U��& ��gZ���̎����3�<�a�#�+��!���ۙ�*�����u^i|�ӄ��M��V#��"y��6��q��!�L�o���&c� �D5��	�j� w��k�w�(4%�5�-�Z��;+��!����U'���V�=6��-.#��)�� �e��}�g&>E�_"f��}�9�ԯ4dy!�^Y�z\���dF������Ϭ�q�����wm���֏���X����ȼ�ۛ��Kݲ@��!�j�d7�%qM�|1��.�����"���]g��� ��In���n��Ȗ��D�̆)�#rV��[N����֘G���CF�R�Y�90��I��+f�w[���Gs��2n�QO}P�E��jU<k�� 6P���K�]���-	g
�DL�qzЬ�����+3���֒�x����	�Bد�]~0�����r��3i���<'�5�xj%5�aF�H��	���m�<pW���Z��b�A+��w謒%���ڭ��@�3H-)!��8��榎��9!m�`S�����-��(�q�U�G ]H�)�]U����()ߊ'v�0�Z�����]��>%���	:Q^�2��h+�e���k��,_�N*
�&�/��t��s�1a�f��������ϒ:�C��\��A�~�v][���:}�����D�->9�'vA�Nwt�],y�Q�w =OG�dG�ڕQ�O㦎��H�]����R�k,Ʌ�AS���� 2x՚�3�-�l�#xdJ۴ĽiV�{�\Hݚ��x8K���;��*��ϣ�U�"�Q��`��1�cɩJX\������\��e8�X���@l��){e}��N���}�8oH�l� ���2M�CE86<�=�%�+���lI�/}�s��
���f��W�}�D\o�s8d�QG�w��rt2�sh��G�4}K�a N��-1mq�tʈ�h����(��A�������n,DwZ-�ʝW����/*�y��l����"�[��'�<Xӡ�q�WWÖ�|h�vKv���y�z���+#�l�Q��-BJ��r���F��)j
��Q�B�m�(&�s���"�&���!���:U�E��F�L�4���p���@E�������BY�푂�� ��Z4���`�s��/T��U�р�#��Cj�ЗM��#�g��k���H@��h"�{�C)?fۼ�$��Z��g�+N���_fe,p ���#%z�}�Q]�u�:�3o�VlJ}2Z����G�w��N8�,����_|���q���=�`٦2�Wv���4�H*E2�w��͗��O۝=j�
�q��p�M���7���fi��<_�Cl����/��ut+n���q�d�ǉL�}!P�Sh��\�,>í ��� �_҉�\0�W:z���o�Zb5SI�}6�[�����S���b��]�(�fC&_���mV���v��L^}m&�3؁+lO�}�tk�+	id.6T6�sx�D���a*l`$�s���������2�ycQ<�M+�jz�a��*�o�pD@��_�*3�:?���ְ��Ԃ��a�����Z��%""rW��P�[�֥I�?3U)�jLڑ�B:50O�@����5���m9H��++y��G�YX�'��8$'�F�M%��߀h7y�`i	�`�u�������[��F�,j|�4��GY����(�j����6�*K���]���s�q#�>퓩�&�)d��d*�!�����pdŵEX
P�2湱�D�u�$r!���^t���7pNLX6|��EM ZC���n��W+TN�6w�"��v�r�T��E�A>u4%6���c�!�j�����Mk�K�l��y�QauV� \�{e�|���z�	X��ɽIǱ�vJ/���5S|��?��c�Y&�ȝ�9LH�A��CF���Mrf�T"�J=�fJ^u�2�+Ϫ�)=�ϷL&Z��($�/V���&f:5H`��O~����>+�w�$px�iQ;Ȇ��jH�5����(�D���r�8��\F?/�(q��!1d5#�u����|T��,W���T���e�UF�y[SYx��0H�n���'�gh3O���z��01. �ؙ/K��f/�#�����'�Hd�{c��F"��Ԑ��Y7fG��gS�0��/`*��:?E�mEC��ˏG� !L��ȱ.u��k6�^�U*��6�t,���(�95Q���o܃��ϣ�}��w�;�3t���%�x\�����S�*ַa$�P(gd(��c��ԭ�_�0�����/��ZA��r��Q�
�A,ׁ�B�p*��H�1�t�4@?o��m�N����$�}���5zP�pd^Þ�h��iK�]� ����B�j�5J�|��#'":�,�"��O�	*�G�)�IrPdAS�)�0��T�Xv�@��Y�Hr�}�L��鹣A���O��XO/��X�PT�Y
��z�N>q�-��)�pG�]-������~�u�w�]:-beK�C�P�E�s�˃�nlP���L��jn�
��H�55���䙉q[��F��վ��HG��<Թ��Ύbn�&ֱ�"8~r<v�K��G�RW)���<��NA��N�\�Gr��������䖪�c�Z\ �M���: QVօCJ�.�+�ގfv!�m|������ۼb�;�2\���k"�Q�AK$��$`n	�[.��k�$ 5މ&��t��_��l�����a�;���_��Lu���p��r)�)��*�Y��M݊�<��4�#�/�����^��l^U�n��5Bu;�Pb֥"�����-�4��lx(����Q!Z�GS�AS��WPk�2Q�6����9��dӆG�t�^

��3cm�����g^��5Q�<kbi����U�<C/�{�z�]��V�W#��A�N#��a2�1�xeQ?�z^��l�[U,d2����2����� }\9Cp=g���s���cF}���Z��IH��$�=s�q��� ��֣w�1�k�c{�JUBr�~�Y����Y��~aJ7&��g�~��F�9��m�FD�Q�d:l���z=0=�A]s~��
XJ��5����P���#`$�x�_2�]�ⓡ;�TVol8b&)�wa��j�-=��hxG'��sz=��� .|ŏd�D��I���;Z@b�j�A�a-\��\)Qeq���t��٬�Ij�ی���\�4��}�a:���6�c�Z���]#޿g��i�
J�@bc-=�+&͞�n���X�ho�"K~���y��پ�4�k�)�S	t�)k�@"T�nZ��U�8�@`Ɠ�3P�c̛MsnN��EG�[C��&�R�?gT�ϴS�]��*��S������#��v�:�v �5L�LҐ�Qѽ!��ǰw%٢D���C��=ձ��"��d���&X��3D�>�s������gErˣ�ܬ(EiQCLnb
I�3����9�@O~�`�{};���,�#�ъ)DF�I���S���i���A#)d
�+��ԥF����%��v7M�[X� ��P��E�2=2�Ė\�����z�L��hm�HW�������/�$���`Q3��"%+o��l%���y�p���55:�������@�gUd<���~�zA�@����]�¿�i���-Rh2�P��_�'N��&\i`��:F�&(l5������S���[�����fA�� �e�9��W�NA��_�y PL��OoЬm�@[ްJOt���[����h���1��r�a�!�����Q��Ci�������w��*f��<��9d������g\4M�:/�=��)t%�g��+��x���ʭ\�F�d�$\�mAQ��������I�+�O3�M��ƋR���Z9������i@�&��$q>HQ��~Ƅ��$8�E�P�a�nM���x��zz
Yn0��9*�����@�<�M��f���?��]�����<��L�>4�DA���N���<v%-ƌ�AER�$v}@��[Y���"ٌ���=�����������F�SdG���!Hs�Y��16o��>"[J@x���Zh.�7 g��l��O6y�/m�=�qJ��J�1~^��O��Kv@C�.�dBH8�/,M����ɉ��[[����P�([#%6�$"pY}���8O�<E��v�����(��� 
������=����#{ ��[��b��t��Jr�xu&ʅ�p]&��,���>w����Zy���B|�4�L��h9��ņ�ENL\��uF�C���IkG�&�\�Cu�?�<4��Gâ"��������8�H.|���\��:�l��$��8�_��.Vu�<B�E#0�E�֑f����ZA��������y_�y�X@F8�^<�_��;��u��o�0�{�đd�e�a��os�FÚ�����!�[5���`@\3����H�i��>����@M��
.���*&ߔY�~�t7cE~?@Z� W"t���aC|X �w�+m�Z�$F��k+ػ�pw�ۇT/���K��s�R�����%�%��Z���0g�;C�I����#�gf룶�(��M 1*3�xU�э:=^�d�Rmʵ�1-�^cn��XK��^@l�L���笝��5���j��;|%�%��"�%���Ep�����4�40oAȄ\D��cNU[~:���8+����<�O�RO�Q����VyMBM��������<f
E�Χ�f���I�<���#"Ygj;ǭ&u+k=��c
��ȣ��)����i����X�ۖ��H-��H�!���L���	���e��1Y�Ѭ�[�-	N�.�1S���|���z*���UH�������4>@�2��_�y�a~�ia�2u��46�G��,3�q��$K�UCY�Պ7q:D�i};�{�uDka������c� Ҟ���
>���v����w�v',*�w��M�R?7��"�w�<�~M���K��Z�%�)*|�y���@Vn3�O�ʈk���7jBU���7�q����H�YH^6�<+<���0iE���<	vj*�[k�8I|#ϛ �<�W������	j������=���-*�>n9��l�D��)��s��㼅�����ҧ�=m!KM�{<*�h�EKS�h�@��!띰��L��U�O����#�|4��Eቬ��H-ٻ|�$���@�q�������G~�PƵFe�T�VN~�~[^Ħ���8p}�k����nV²\�>�x|���
6C
p�̯]��8T��S�^ݥ��(��k``c:l� ���Քw������(<#�UB-�r$c�X�'	r����~�׸��v̝x������5�ĭB���ui��vߣ�'���Y2c�
}۪�-aI�bV���w~������2O,��xdODH�$�l�I� ���dBޭ��D;X�N�h���$Uف'�s�o�����rC<b��i���t*��H�x-�����߫����a�Y�|���B���!�p�̝p�W�ӑfډFޮ���ƫ��A�1�@0������1��}��)�*�����5�쨥��Ձu��:��.x�T�����	�����	<��Zˢ���2c�x�*�[9�NA��Y��;��%/��=�q'��|�B��J�t��54,�i��������#o�� ��M�ٛ��V�;?�kw��[mf���k����I@ �>A��`>-�?o$b��9�lF��dӬ�"]8 �d��'�'/?�Ð
�d�u99�ŁH,,gcc�_�Cy����\���� �}U�y5+L�����9��Q���K���]k��j�+Vn�
�U/!%��G��Ep�d���y-�H�|_J1��G�8��c��|����T�ehV���-'��V�Oy��yQ�	� ��3�W��p}��)6+�z�]���R����|Y��)$S*�IXf��-<�$L��	�4��j�\͑��%e[8k�<���Qv�lգ-�ؚ���s���杺K�+�	ӟrC�P�"�m=�%����&��4���z/����1*�O�x�ylYgB�'ϴ���a'�7�'�CW���/
b��&���"��U�����_U�P#Kͩ��?�?���9>"�|�#}"G��N��h�'ϵd�6�H	�P^<�9P����3L9��_{��%s��2z��(��ѣ��5ڰ'�&F��N��N����P�Lk���Mt4��8c���b�֋�,˾���?�M�����@u�q�xs羦�D"�z�=��%Mm9k����/�<�����"v�
���8c��0&p�dz�ð�x��*���9�{�Xz�Ǒ����n:%������YD=^Q��k���Hƫ�ۛ��:��|�Pt�a������ ��p���(�`��Z�tdCNfA,*��@�����==��� {]����~@�::? ��_�㖂A����úGK�2��a�Msp]��BN�����4�-�@�tؒ�c�:�u��_DxZOW�86\#��}��\�a7�X�cA_!�Ly�5B��'B�ۀd���a}��0&����Zo%�VL� p�1D��?x�zs��X���C�Ͻ�(^�y��P���zFw>ڑ�y���E�W��H�X�y�leI�w��pZ7-�f���k�99s��k�W����o���:�juz�m��g�$��\����d������c`�����%E�b�<�NѝLM��5ֿ,@���}��&�FSO~1�M��
)�=����ݨ��qI� ��ť��Z�߅?�Db�8��]�6�s� ��h��L)|.p�J�4���*8¼�ڋ��NՄҚ�*�W9���Uk�n;{�H(%���M�o6�w���)�i�O��(]UJ�7��E�EcU�䠨*���g(5<>�&�T1�-�d�h!,P�-���N���^?C����Ř�lS~�j����ȯ�֯����gr
f<�2Vz���E���#�lJ:��c�Չx�/�i� 
q�^F�m�w�Bpf��7l�(u�ۇ9����~+v~�9�LFU6�k�5hx�|8О;�-�jC�,�{S�t�)������B�N��?ʎ Z$�O�L����L����4$�;8��ٖ ݵg�h�Є!6h��>U��r�l�5%��o85�"X2Xo��Q��{�䱶�<Z�tτ�kB��Gq�f���ض	�X�󂏌�'����I9���³�lL|9�>ҩ�-S�>`�+l���t��19	���ļu�Ϯ�pA;��l*�?���j�JZb��9�a�f�z�r�����/Bl{5�@p���*x4NIw�y7�pI 6�ךa���|$���2�����ȏ���h���{��H���'�b44)'���@��J��-/s�U��G�ַ}�)7��
�)��#f
-6���4�~���gxj0�Z_���;�vX�m��/|�+D7$W�4��g���Ōw�W�JB&�H�L݄�kr��@�d^G˓���%��5���:�M)@l	�c�LYA�6���`,@�<�
~�C� <}ps�)� �_����CŘf~J%`�@B�\��F�����Iu��j��#���^ҥ=����-ݸh���bx8�u�O��(���J�
|B�"����P� G�b��y1�W�B%�ʧ�iq�*�F��.Ϙ�'�(����D�� ���x��Q�e�!su��/��v�?� �^�(�ŋh)�N2r服灋I��l���c�9?��o;ub�"5Y~W��f!�0Q`�H�N�������"]�z5�{�9�e�)��-ncxY��[W�yn�nE�PA�$�(�1����}�P�����I�1C���T͌�Ha��~š��p@y0C��52r������vPӒϼLd�Gݦ���$���du�F���@<Q'
2@?�$��L6di� �E�5�A	��3�Ds_�;����J4�e�5;�+�KR$> h��_������i�G؅9��*�-7A�kg62�kO��w��k�!.W�~�^ƪ��ҋR3Σ\�j�e��vN<������D&���'���.OG�����[n3ߛ��>�jsH�#Q���o|wngLZ�?��� �+{�C�f[�P�թ�����g}T��t^�
 � �*��Tr\���1f'CTwE	��r����( 9xf��YV�0�T["<��{6��t�i�X��\�=
��"g�����VS��X�n<t��9�[�|������CC��7_�����2��:FNL�?��q�s����q0���1�Q�T��@����*Zu�q��j�(1cUPUI�ͤC�I��M}��.��m7DwR<��ڀ�|��_0҈��;o��^m�B�J5Ҵ�5@�4ho`�gU�ɰ��:�b2�[5&��G���AeQ�A2jo�sYQׇ^���h0�� �A��w+��[O�;0���Y��j�O5�h�j53b�6}��N�3�݁��'�9�v֤z�kP�4�,u��j�Cv�>�y����ZB���%���sX<�̣�3h&p�g$�lw8!"h�ʬ�a��ɂ$���7=����H>�yF5Z�@��JLYC;��iO�/4"�`��r[6(#�����-��O�vv�!/�z���*v@�NX��s�6�&;^�&�諶�5lu��;�Xb�P�|(h�L��}�:4��|`�g��a��@�,�� 8���M��ĖTj[`����1�=ް������ѭo:��8��8�Κ��f{n�BH����Mv�,�6i���=�o0�`��b���"�K� ����]�/8���t{�;�f��hk��3l�Ѵ��TSGF		ꅙ��LM;_e�l�AD(>�`7�"p���}��$g�H�$�%LǬO�*����3A�;���F5���(/謜{���>P/Y�w���/��a���gAa�j.M��Ѯa�K0�9�"LpRa��X(�o߹tB-	� �bdh�<��tYmE���|\M�*���E#Q�g/R���]�j��8[a��r ���ؿ��I'P;Eٟ��g:"B�Q#��
H�3V��@M=��X��$��򁢶�a��/���dW���� >WGe �͔��Q7H������KHS��sB���)��0���ݠ��Uy��@�h�h�;�/����l�W�f0ZY˜��By�7�4��%:�gg����i�$5r.��ʳ�����F��{�F����t1��Q���"�0��<�Q��ʱ��u���My�7`�����H�ҚP���|���7ω|.$� ��ЂC�-�]��@d�v`�<eF���ke�4�_c\b���s����#�fM�
ӝY�M�����v�+t�u��hg�"G�2�'S��z�>�z%�%ǓDPm��M��b���5���p(B�Raݑȯ��`���q��(	NB���3�����|��O�:�f�������lC���oe9�>��`��&�/hy��V�ҟ�i�
�R�\�8��G�Y�����a�ųHr�o�o]N/�y6�P����jŌ[ ��<S���ýn��S�x�֡/J�F�]���ϔ������	dED��*���g_��w[�~\
�,�Qt3pϔ
�u	��I�f|�▅ɐ�X�v���
��қ�����n�P��?��G�����O���%���#�gmE�}�^D8��w:]!k����f4T%Y�I!��]���PF�^�(�晛����j~�Bt@���gT �B��XL��n�]�@b'��	������`�J
��RZH��b�G�5ڳ~,��Y�5�p�Bm��d�QYF�2�~�;��1Eg�8CB�:�5��3L���P�x���������AI�gi���E �������I��/B�Yx�i+!`)�(%���b�����4ӥ��|3��M�'a6@晲��#�;,E�S�&K/�+?�,^��mt���x^�t��i!�ьW��0_���0P�|�y㆚
2�z�
gp�5���C�X�����W��d��'U�uτ"�����9V�n�]\rO�a��;��/���V�T��vf����ޥP���:;_�����w����$䥬�����a��?�ѲRK�F��
q���؊W���e�z+	baݢ+pB(���8a���9�@IԦ��2p���f{�P{d�te��pų�\�RS�׃L�)�pƧ��ٔ�G��ihm�f4�7�م�$�Үl�q�>f��Q�x:Z�2��s�D�M�WT!伅fX]o�]4A�$�;�~�W�C x��C�s�ὲ�pMՖ �/8��[��t��n�;)7��?UG ��~�3(x��b������8�4��+������\��U�=
���~�V��*]!��Űo���BSk)2��oCq�3R��bD�:��WdI/pHE!�3��]a�ǜfFM�X��8�߈�Օ��὆��ۈ	�!>z�ڙ�-��O Pm ܃����O��C��3��"��{����Kپ�X�efW<�xSؼ<��B�\��!ц���I.��R��95�$PY���Y�p�+N؃ԗ���ҁ${صԔ�����`��ÚYwO��5����s���KPu��lʿh
�υ��C4F��˛��f��0��$6���K��e7q0п�b����e9�(��x��z�;&�љOzP�E^��>����'�x���2�.ֈi��,ڧ�1�"X�2ۦ׊��J�����Z&�@c�@$�ys�[�E�����;)8=�y}��D
_��l�l��H֬�3o�2��������G�lM����|f�s�u��"R�En->���Y]�����~�P/K��9�y臥��	]��*EXt7D�/��c���!��N5��q]��a�����x�����P�S����4-u�Ǔ����0�(.I�![���ǔn��3�ʀ|�]�Ћ���J�t�9�iۗ���Ϋ)e����n��
�=�d=ɚ���(��=]���J�
#QE��&��Lt�۾��Sf�JR�0���@)���՚���:��X����V����3�����f�ѝ{��p\)��=�
Iަ�@U���=H�������A #�\Ot)r��} �� �w�v���=���BI�VGԣ��T�t���`~q̣ė"v��8-� ��k�}�����͆��[IܛB~˸�'AX�P�BzfԽi�//3������Ed���"�x[W���4B����(�(�,�Щ|=����n��2���/�~��DҦM���x=�(ET������T�����(N�졇f�ş*��:���1@�F&%�q3x�*��jdY��3��`F�%z��ϴx:(��B��>��m���Z����?����c.T���m����\�3 {�#i]�?L]b�V�s���J`p�k��욵�t(Ո�梨�
�;��Z���or:�Q9�㳟�e��#9�D+nfHP2��O ���sSQB����F�K�gv���_)�TP���'cl�+I�pD�*���{��Xg�ow>��m�����M=������P�"�CF��Bp���/qOe�^�`�Y����J��_��C�]y�-tz:]-NR�# �1�ձ�,MG5� w4�@����+k�w���a_������L
h
&�M#r��4���_�?]�'��wbĬ*yv�^[(�	���r���dШ�Z�"UM���0��7D�uv༖oK�Z!�Y �����8�w�V���Z�z�MSU�X�F������	|d	n�QQt""v�mr�q��K������X��ٗ�����;�Нb���hz�C��X�xJ�<��ORԙ[�0c��ѓL>��>�y�kz�E+�w��xͨo��V���阱p�zs��#��89���7��7����Y[�CF*EI����H~�f���4�6-�ڔEd"�R��qH��߻������N}D�D���8��\ejQtP�of�Ǣ�ԯ��0Z��W�*ɣ�g����A
��&+���U�D����5�m�#n�9ג��ej�CC�����7�c�'���	g6�G}XO�r�o�(nD7=x���o�oZ�����Q�0�x{� ��&Vj�7��A�EVC�Um�M������!��N�'d�����i20� ����(v��n'Or4��'CPT�>w��%�Tm���]�DJ�jQ�G�����ϱ����v��!�u�@|5��������|�7_�8��B\:��ZߥѾu�i�T��]-�<R��IAF�IZ5��} �����:����B�a��<�+�&�-�Ϸ�n�m���ރ�BC��8��E���d��<&��T���̃.�� ����D�Ѵ�� ����<RcAU%8��._�2�~��K�[7peŽޝ� iy�h��.��k�WMk�^�~��zS��G�x� � ��M7Aw������Es����+D��0������\��֧OC��#;��t�}�ʳ�IxSFMNc���# 9CWI�ͦY�]{��I�n=T����c
�
q�&�ܳ`���q���4��K �����" j�ܥ��IBIv�"�7���z����8E��ÿK5�rDt[g3r#����=,�o8fB�>�7%�Ě�ü������I.v ��A�.�L�ٟ�K��[S�s�$��A�r*aA�>�9��zJ�n��]H�D��f?ӣ|����	��#�����br[K�}wB�fu���~?8��fc��j�c�Vz���O�NП�tX;`<!�����^����c6���:¤`��ʛ�%����%&K���r$��U'�!�V[����-�>)�� �&Xݜ~Ó��LcK��Vx&Џ������.�Aw�q����"�S뷣0�ޘ��U�}3;bd/����J��c,���Y~K�)�0�����y�A}J���?!V&�X[u�=ә�5�v�>�y��X#>n*ʩ7?S���z?e4YAX笓���*{��<p���e_��2�����Ђ��id3��?0	L2�P+�A����(���wW%B{�=u1�j/B�++�1�.�h���=���@����U�������E6+���o�U�y����݄W������[��1U���M"�f���P{ FڶN7M��a�hh�����}e�(v|-b;D7-|?�F����n�aX9Q$��Hi���OR\L���I�++O,�����E� 7�B����(�}�=��^7�:#����*�yIX='6ɩ˦d�W��+o��^��BU�X��[`�B��e�U�/<��pԩ�ڔ`WQ����w�5˅��ɹ��5oY-Mx�c���JWԌ��]�@eX������S w͊O�dmk�k'��+�Vw#�f�BM�0r��c1[����?$t�#���I1=̓<�)D	�F�|5YN�p/���
&ײ�ڏ���b����+M�U�Tk��-[mq�YG�c�]=��:�Jz�`��lj��XP�����k>m��&{~��ږ�A/���?��M���wl���8E��w(��%Y��ׅjs
柍��+�`~$n�+�;�#����'���"�S�uC���W���+d��<^FT;yw��>�� _��Gm�!un�=P51�?hs���gW��v�N��-
n��C�å�
�m�,�.�}�I1����yZ�/��i����?��}
]"��7$퉵Ik]%V���N��k���rAh�u�*d{w����-/.��*8 <�{�)Hw��ʖ{��r��Z�7U�7��v:,=+�������+���Ѷ�ٌқ�~f�52d"kWu�
v�����R�)��r��4�;{�^t�B����'I��WI���b# �~g����'����6���-R9�Di2'���l�$%{��x[�X�Ј&\�$��qۨs1ǦdK��=�\��%oj]E�����e&D�{2Uk%�{&�<O�,6�l.��"��(���D���z%H�~'�)��:g}' ,6n}P]���Z�����߮�b��Ċ�D-� K��X��g	��R΁�\%�67��G����l��(W�S:����;���ǲQe�^V�'}�bvoRN:{��4^SXT��i?�r�<�Ĺ��΀buQ^Ȣ��Ը��G�6j��zMI�r��u�DD�5�.+��o;;+MPS��89=���n��m�+�(ʄ��<�ĕo4E���?4�H�H��1�f-�Uww�������]��3Y'@�|ֳ� \(:bH]cN�pd�|�u��^�;�Q����H&1Ƴ�ju���&����2��v�T�V��xsu��<��ya�(��F�|t�04v�ՍUuR��qV�C��q>�b��o�g���х&����Du�I������u��XB���aV�|�g�Ip�a���KKz�`�&X��V�A���\����Y��Kػ��=����+��7RH���h�v4�9Z��ޤ����K�9文�D8�4���)�i���)�q��Ռ�,d<���z�bHe�Wyc��
]�I��t�M�����+~v���P���@Z2�����G�NB(��+<KV$�L�#��Y�(�0�/x
�a��l�(�����mi�q�XԎYǎ�skd��%v��j��,�����A� Ӗ��q��:�%��*Ϭ��<��l�6��J���[�*|�f<<���V�?:�=��ʍQ6M7��9���ytIy��3Y���V���Mũ��eg4B���q-��]puQ6C}�fG��&�Kl��bƺ��v�5�*�D�v���m'C� )/<˻h�w�����k§hː$�T��#�o-� Y���8R��ǐ�;"?�%�ӗV�J�G9t]P�ئ(���n_{��#X��W/��l:(��`���~��"\�X	�gk�^(��Em��c�s��v�pt���213�
0�v�vf�7\ﲷ�8��+�헆<�Cz`-6�ق(.�R8;����B��.��I� )E9���n�N	`�=I�2'|7�L_&�Sz|^Ŀ��A��4^ծ�Ղ&``A�R�h��A��=&?'O�4o�7�j�}��iz0?<��b�aXͫu�%\��	��q@@EϘ��~�����]`���L���cĕ�[Ľ;M��/��揁�>UO+� #0*���P~QQ�A�6����LG�<���t뽠2�nc��?�3��`S�L�&�ە
|e�5�C�5���m�۵��d��/n$�ؖ���٨�?kB��E�0����fO��?��^C\�#�1Z�{�tJ�I+�)�iI`T6��Y$�f_$y{u� ���խ�p����A�;v�@�Jĳ�yr6f׊��KKϿJF	�O�N\.�B����B�	���F����$S��Q�yt
 u1���ՐK�{�#V��$�,)�c�@�M��+�ߎn=���8��2�dW�����T�jw�;�^����(�	���6bY��S�}��N��f �Z�`�$q�r#���f{�f��1�J��q��SX�u���Z��(���L٣G���nQ�s��sV�i���~[m[�|kz������	ɚ�� b~%��(i�:��G:�������1�M�q܄�oGD�-��=c��
!��#x�E3�������əir[ܿ� 83�UJvTA�d@aJ,j�u V"�����Dw���"y@�q�?"�`7�L����X���%��cs��j@5p� ���&v����@��-��`���rl8I���}�� ��L#��'���E0z0l?">���T��1���v5w7�=�}������p�ͭ�UPU�a8(q&�>?��ad������/8����COkL�i	��B`-���^2������\6��� �����9P.`8�.9�yaβ�Ğ���Xb	
yz�ROKY#^"A�β�d9�	f%%�q�m��]8����嵤�Qvѵ��Ɋ�8"�@�pn���w���^�ؘIɤ$��|��x�\�r�Y�5ݞt#On���c)�;�@�u��J�9�ˆ4ߢ��,Pl���`��t�����7	m�`Z&��Lq	���Kmp�A�"���C�������ug���L���Cڍ�^�';����t�Ҟ.�?�Ĉ��z�r���@�2��� ��iר8�^��ʰ��2�l'Ԙ������5�+��6\9��D0�$p�dzv>��+�p��X�'���V�j���TŌV��DH�_�jk�`v�s�[�C9�n�����D��(����C i�՜�iq�\����T�T
C��qF��u�7m������U4Y��J���i������k�J}�'��ˉ$F��c�_<�@�c���1��"$�-���D߀�E����H��^gW~Q�kCW��R[�-�x���}��&��`�gj���Y�f�dqT��`%��b�*z(���K�ERO�禾����(�bt��	��"Q�;��3�IK�� ȇwA}Hc$c��WIQ��4)d�F�'�%�1�0����R�w�D
�c�fMR��^�f�M�=AY	�y¡��u��ph���tH�X悩[Mb/�n�c<ia^�h�j-<�����IWa�P����*���s�c#��`y��?���"*�]此c@�}�F�7ӡ��GWr�ׄ�8�lU8��4�žJ���8�����ۇ�H���6U���16?&
-sfU�6誊g��G��� �&�~����c\���/�[
����PZ��c����u�y6�#ڣ�:ẏ�x�ˮ�,,*���F	��9�2w�[�A'|��g/D�ak"��^x R!߱@#A����/�_�����C�X�.;1�Ak�J��RfDr��w�@R��T����O\��fS�ld��1D�72���`��A�G�"��S0�
�pI�uO��f �8UW�ɯ>���~.�	��+�Ps)�3;���r�
_^ikd������M1�5sUDs�k�颂#
���c�/��2�*+�
s\�~�A"����H��iN���w����н���(e�������Ѿ��hvU��Y��pt��	�ꛢ6V�MeSj2�Z�y*�
��ʭ<��(e�J����-�;Q�LC���>�J0�R=�b�I1c4�Rw�-���~u�0�����k�%v�`��+����WW��QfaC$��1ɥ��I�-�r��㟢=��en����עA�ߜu�tR�����{���fق���RS��M� U+�w}<���]�
`C�o���$f����\�ܿY�|)!@X1�g�1z*�u��sE��l�IQ��>�Tb�L��oO��iL@��BƄ:�0�^��s F�����PGe��\e��	t�u;� ����I�����t՚��b��3�O�U4�i�
����%��E�ӳhXZ�.�T�1�m�7��wwE^0��N�5��d=J�d�O�y��:��<<�p�$��f�(��+ �~�]f(Ee�$�z�9���\����~.}Ƌ\���9iݎځ5��}|��U�ї�|X�ņ�i.vd �
Z��=_�gku�/c����w_�r/�g}<mHS��6���SI�*vR����%�����(�د�q����/I9��g� ȗLTx,AA��/���۱\�_2]�xL�u�mAͭ�U �*F	n}��.��-��#��I�����!��\���|0���@	��t�c�l٠
�F�1��d|yH������џl��,�EР,�%�v�X ��1��	 �{6�'�ּ�~�4�� ,��.ꧭ�\�{R.�H�y����΍���l�ZLO}Ӡk^q��*דO� a>I��I{��@�1�ƁHP���9��^�M33z=� ��MO��պ��iO
xÑ��+S-�c�H������a�ށ���E��d�Hhh�*���0}��hp���)���Ch������ξ��	���~�SL�o��}���,���;[p'�g�؈�����+�ыq{f�˲�(�)q}Y6��_�l���q�V�W"��!Ŀ'�1��u���9����U�?�u�z�B$R���U�$S ��QN���gdֽ:�]��j���t_���K08軔�^�b�3_GX��E��Z�!��%�G�O�8&�Pp������v���6�o�]�;#ݶ����/#�A�i��1��b���/��Pv�p�s�Cvz��4HV���ɖ��&���$<%�+�RS� X�wחn]s��'?�=����6��g�� 3�ˮ`@b]�v��`��U[� ���~
��ډ�i�Ml����+�KF3�&�}�ß[ĭ�nI?�q��.�递c�eP�ż�V��N
��4m�'rM�4�w�FHaډ�K#���� �΋�\��*�i��L'��Tܿ�M��S�s�߷-�<呐p��k�N�U���*Cք�)����3�B�?����K�d�z��@mv9\�p ��=w�^�S&����eXD�~��?N�G[OA����%�p�2�>TDA7��݅,��jN��k*C#�����ag���9ϟ�J'���~��ܝ�w���aq.X����\͗u8���=Z�O�VB�`V�U�!��3���%	�	��(`�$i����%�.���WP������<B�e�A:�oW���8E�G�ͮ��B�5�	���K@�Nm�uW�x=f!ߑ�0�X~#�-�RB�(�O/kk]Q�,��If��:P���&���z�X6�T9���5�`�z��-b�cE�LtZ�D3m�Zv� �&��H�H�`��F�SA��CmM%��/C�6��{��ܜ~i���Y��YdZj�^�v��!�((���\x�����Ux=�O����Td���N�St�}��é�ϻ!���pk
�D,���K��sT~ϥU��x^��l���T�ñZL>��1�5ɘ�2S�U�W�u@� ��Ka/���҈�3`��X&�J��^��证�x�ǎlS]u3���by�CȘ�p�ȼ�3�]Opx��P�������7��@�(���Uac/�i9���U~^�Po$y��OM�G����q��q�s�會�cx�Hۀt�g�TP`
Fm <����nL�`���)k�iʷ#��P�e���4���2�Wu]�xW�@�����(Q}�
����טsi�w����$����ˑf��
�up��� 8>�#�c�o'$<�l֞��N���tOW�B!���7�g�8�%��4�S�$'�}�~�R-&�3�U�����÷�d0(���E�[�e>�^�曖�W��	u�*�N��3+����ݏ�b�V[�t��i�E��TB~����W��阆���Ĺ��a�[�-8&kR3�m�!B�/qV����gs7��.HR0#���u�/u�H��51�p��ZF�(�3��?ߠ����E/2�٠E'�����U�!;i`��yg6�.��E�t�M�b�C���o�"j��[�]'p�K��l�o�b�p�	��m��h�
�.R�qÙ)��*������c@	t�X���2s;㧉*`}]�Ht*Ox����x�	���f�jL+ugđ�d;R9"ݪ�x��:çʒ�,�K�����<
-1f���g��GI���@¨nr�`تu��,=,�>j7�'�j��(
��? $����nۉ7��&ȕ�dz'����le�S�^1����DӋՅ��-�k ��bP2��"������s6(�Wgn�k��-�{$,�C|87��Z�7��l�{��\G��fQ��~<��Ձ��B���=�����F��h��*?Y�jRϣ�h!����$2G��@PU����Y�X��&d��Ej�ƚ�:���ٜU��M�/���v���z���+��[n�	�ũ;7�7p�H�y.$���"zMg�|؏9�z�/�!��k��G@��!d�G�T�Eh5�)~�~�y��	�u)yK��wk���Bkܗ��;�e�\(p�5ٍ;j�� �$���)ī!�;wÌP*DCo��D�z5Z &,��u��kX+�g��q(yt�c {��a�`�oŝu�x�ArlTD@RF�~G�4˲8�@be�G�cKH &t�i���f�	�n?��Qۣ����&�K">��C��n�8\�x9��r)�O*Q�-���6��26W��n��Ü����+2�T��X䏴j
x:�{f�V�MP�UK�d�Ϻ�t���ś�{�~����k��:
ֹ
1�^%a���l��eH�*�E��`j�ID���J�-)�l}�N@ɧ$J�׽ge��rA��Pz W�?[�+$^"-�XƬ��yK��H��7	<��Nr`o+�h�H������.�V�&�Qcǳ�dp\��#�^���h����8v�j�^õl'�!]��4�_~!��V���Z��o��[m=c�����;�p| ?���/�b-�oE�����^�,�Hq���9%y��b�@Sӱ�y[�������e6�.a���=�#����c)Ϩ��j�;�FǪ�s�ʩ{�X��\�oQ�:{
҈Q�%5�ؒRC�[r�Nd�-o��+�,����s+o�p��*�i;D#�s��E��]�L��9h��%��#��{<�����(���{Us����ĺ�Ga"������q�V:{](��h�xd��&f,"��d�4���N�}�P����5��&q�iWI������AN�5J�J� S��g�Q�t���Avbi��Mְ!�\�/z~�q����z<��T��HI�Oչ#���܀ݨ����qSȀ�v?�Hؔ�PU�C�߈�nD����i3L�u) ʰ\�2�Y���r:��p�T���yTr#��;a��>�W������(�6�Rs���/�<C:.�r��﬛jF<y2nE)���x21���9�\�E��^&4/.+.OX\F�U-�üp���@7����x*���Dc�X��D�tOjǬ�6`[_;�4�(����ʃ����)�I�:"|>m��恻�e[kL�qږ�S�� �O�>�nϿc�~�B��r�Kd�ސ�-�����	��P��pcv��_$�g�����Y5��%�Z���U��{Ʃ+��IG�9Y%+���p�З� X�4��X���x?��\�~'bw
4�<_ُs1�J��P���զ�n�Q#Â�`�)M�AZ�fH}��ۏ����>��Ϩ���]��r�����_]`���qs2�kW�R��qŜ ���B�Q���̘+k�/�O�֋���c@���ER�ظW8��~R����dCF!֛3��1"k��>�_v扵f�!����}�$x���t>\4��a��!=����/׽�:�7ML���ڇ�1ӝ
V,�H �"�b&�W��g�8�.庣?4W��CX��gW�ޏ��WFMi��O��-f����[��(�TYd\�6���]�E�����{GD�g����+��F7����*����g���ы�F)� �m�����G�D Ǎ{����ڝ:M3A�
�U%���~0ɟI��M�%��!�����8���Sr�����k��>i��H��1Ff��<�RE�8�������nO׎�[�xry�X�Y��DW�N���:�ܙ��&�nc��3Kj����`��	W�������-oA����d���S6JG��4����õ@���u�^�aB`p�������KNP9�%��G�a{d2�3zn�qU�P���c<�Ͳa���j!/m̗Ӣ�c�L�9عt��|\e`0��^���[����% 9�XI�%8Ƙ�}�����p�UJ~K7-Oԉ�^�=S.�� �V	�ǝ��[���N��;&9��d5��-�D�EˊD���piz�7Hu�@�@^�"�y5jmՇZ)o���ڪ��${�3�V�$'$}�x5� Z�G^ڞ�e��*Fb݅f˩��Xߜ�?��z*��m�%������:2i��oO��
f;$��f�W;W��]�.&㄂�p��6���3�c<݋֔��q��֏m)4�	@XzV�NB�.�p��=�f�j�s��������"�M�A��:���0�!��V��6�y���BƄ�0�LM�c��v�E��#��S�̢��H��eLcAZ�Se�
���X�'�ve�(:0�µg̭��$����G;G��Z�a�5�-�iER�d�L�L���i���^F��ćE��8�I�� ����+(���0������Z+�����x%c)�h�EGn�Q�T�zč�7�Ԟ��]l�ژFi30�"�A��D���V�77�>֍��Ӊ>�3e���Xo<��d��FjҚ�̄�lhH;��S�3M�Zu a��M�Trn�b����W��K�
�$q�D�5`7 �_���=i�j�d�݇aZ�x�{�3�'�c�j�lo@jX���:f�DA$�������WD0h�	��(���j��ΌR6��1�6Y�>��jc�[�x(�;RXXM��X@^G��m��������iX��[���(Yc��;/�"�������a!��>T�2T1�����nd���f:Y��aG�����Z~��<��2�W�ks2�H�-�Mz1"\���RTv�^(�[��J!�����\Y?�_�9�ʳI4?�?(*��}���@({��� -���V�����T�I|�S��?=����}(y���*�M*�*%�m�sv���&h� ��jSBB���U��h���=��E{v��計�a�D��T=�v�G�T��og	��F��2;IV��" j���p�Эn�u���ŭ��$��xm�� �r/w�4LܷN���XJ0gNZ�7�̲����pzF5k�LH@�ޙ~�ۥA�p�Բ���w5ψ�/l�N�b���T�غ+5�j[�hP�Hk�Q�f)���U���If�bdz�
�c�-��h�� UL��� ���*�]�C���G��v�(b��z�xfa��.���:����n:*g}�a��]��T��}���:�w��0t'�y|���*uy�#������{�o�jamu���iWp���6�-�o�"��P��&��mf
@�&��S�_�8�M&���0<&*�
Z��n�Wcb-��I������kcB}պѧ4 8�m[�R#WN}���(W���@�_WO�I�"��.���ບ*O��0��VT�$��>�+��i�+���_S�ˇ�d�gN���'.��sS3�ıb`'2n����������pX�C/�M��]��l�`�qsSm
L�q�jX���`�\��7�\�z_+���WG��'0��,�qF��$�ODr��{`ˍ��`4���*���-KO#��-��a���Y�r�������|h�OV�j����Բ~4k7
�I���Dq���>�_��{4��ÅvY�Jr�<��6GV�jn.���ba��ʧ���m��Y����x��
�u�IMg�-;�q8Y�)�����# �냏��tM�5�Rj�F�ʃ8��2��T��/=J�W�����$��݂Q�`�OR}i�WS|m��fќ�>E�����8�t+#b`����װ[���QUwy��^	��I$�I�������K�[2}1O��h�@s����w��a��_;���"Ւ�3\�	m��M��fǋ3lKS'�|��Nvә-��oE�����ݟ��*>��C��5ܚ�Qd�[)��(������3=sH�,�(uljF�9�#%1����=C�B���a2)%	A!`E�:�O�k:I�^��o$9T�`:BW!D)���#�I��E����Y�9 e�A
zj�i�ӂP+���_η{�<���oj!�c�W��tr������J�c�]��t� G�F_a
l+���x��/Yٚ�v.�x3�U]v:sD��#~�./b�?҆���yGkxR'��o�[ќ;��[��	8h�K3!�M�ғf1@7�?�a�<��l�	f�fʟ��W+���C�	{b�߅�f۝������s�2~NKR81 ާ�}�]���΢V�,�����r���]�+�x7���qj��.WH��M�1�GG����y�O��tՀv_t������) �1�ղ;#�����V����5n�~�л�N�(_ndݳ��n5J�����a��8�2���
Q�K�V����8wo`rS���;������$)(U �ëxB��6�s��]mtmp�!����~w��4�Hx�5�ڎz��s��sW�ӕ>u�G̼^L"����Ԍ#I�֩�n��G:���D[�+�Vܔ�ɡ��q�b���j����DTS̅�E%d��r4ύܧT��7ƚ�<D���C��s��_���4�>���/��*m�� +���?�4���7�5��;�����{�Ɯ)s��b	>2�Y��3��)oK��Z_T]Uwh�W^�Ds�&�)�^g�M���S ���!Hl�̵>RU�#b�g�䀣���|e�����	�;iKz7�y%�M�	Yy���6\�F&��B@���������������G�秭��i�V����T͉�M��cZs�G�OXEǧ�a�j��6q��&T�$��hː�si}��gB���hkh���}��zC����Kq��P�N�΃r�<W�4#h+77L9�:g"W��/�:�G���>��������0m|/�0�1�A����Ǿ>��7Gs�c�����mm���-����,����-=�3u���?f��y��q'����,W���g1~_�^V��`O��4gO�7��-�|��IMJ���}`v����<�����~����������,��jU��њ� �vd�(�����BGrY-��+򕀥�:o]H�"kaH�Bg�V�H�^i6y��~�n��#�*��R8�4|,�`|	[������7�xQ3�9�#�$� ��� �ۿ8���
�\�?�n<��Q��1��a_��g��'�z^�aݦ���fslʈ����H���0i&%y�HF��I�Z�G����|�qz�ή�Wp�u7�2������/��1X�YP�y��_�0�����FA� 1�`�8��۫"�b4�l�R�v�&���@.�^��:��&����o �ٝ�¯�8�B�0Z�U[���*삕�3�G��9�=��Pe�9��=*��6��z���1�5aK3S�֮:��if��mK�4|�"�U�������b�/�_��?F�*��0ַǁn��݁�(Y�4��ctji�����7<5G6�;��S���ۑ8�Q^��vLE96���p�}�Iu�VW�܂�zKmi��xs`��&��7�X��ZR*H�i��(P��XIL��Lqį����P(��ZR �jܶ�P_Я��$�Y�\�˛%"���pʿS�T='�%���!cdl�D�`C�Q�(�`�Y���G)��l�|P]��W�� ������Z�uhM�n�wU������Z��72s�ʄ�i�ê��ڮ�}.��}.����vL/,������ ���1�J\��A�?3�U�=�)�A��\1s'�Le�M>�̮�N��魳y�����O�o��5
I꿿%l^�`���,��LE�.X5s��`�7(Z� sWZ򳧏ݞN��m�`�{8�VKk��y���b�f�m�� ��\���ԍ���Ķ�2��(�{xJ,�Q�A�Iv�H�	:>,���8�aĥ��r���:@�׮(���T��7nx����I�]�����>=e�\<iG�e\�u��=A8p�.��O
��1�O�p�E2������Jt�.�Ӭ�O���V@:��<�������F�yO�����H�e�
=P
���b���^#�$�l �Ov��t�����$P�D`��A����F@aኦ�	 �RM}sR�<9Ok�����2_��A[���A���f����߫�ZGS1�M�����h�_;��m�Fޙ=2|�W��}<h����J��F�*Xe�/�.��Dp7���U��4!Ԇcv|��hٵtv�?���Yؠ:�W{��B����^7#,>�r9kɐ�
oD��B��1j�C��0ny\��u6^q�A��ݳ8cr9�Wȶ	�O�Y��ܧL�տ\A�_�Rs��T�6�1e��T^�ќ�`�|��	;�DO3��|�ɶ�Dv0�jJ���^u~��=JC�,�!�[g��(w����ٹ�At���DOL��z#p�X��@���	֙S��h��嘶*�pǿE	gF��k��� ��3�s  �P�u9D>�E|s�ˉ�^�� 5ȓ���V'��{�V"��>�~��/W�n�e����#êB���P��8锖3�2.�R��x�n�
����N4��\�֤�o5?t�.�;�@U�Y��Ө��#�"�Ƿ%~^�j%ݛR���*9���Ib}�"ɮ�.���������"ΥG3?B�t��I���vn�| pU�=�Ph!g\_�g*Y��7���Wc��;��W�I*�*w͝�2nf���B�>����Iހkl�U0��Cs�.��:,��bb<�!`G�m������$��/\OB�*B{nxfI��:}��"$��Y�g�=z"��'�ں?�)��'?�sG�'y��ۀ(�DSږq�.���ة�����(>9͖�ʸ	tr}W���u��HmH���3�#TyX^�%!�$�7B���!t���3}R��A��\6)&g�:3�n8I�ΝY�k�Rx,��]�M�>���]L�;z�j���i7di��J�$ޙ@�l,26�Ϸ㱟S�Df_��Dw�쫅�G���ⷵ*ehc�)��^&k���g���ݟ�!��:������{�t,W��� G4�޼Z�3X<v[Vb��j'�t����{�G+�4 Z���|�RQ��ҕ��Bn� D�H����Bwq�a�W[N�>n����Ϸ1��-��
�1��#�
�a��R�q����tTh\x�()D��*���LC5����2��h_�5��ډ<�c\
?�ޓ�k�7����fX�)2./,Oq��{��ͼ�N�Ǵ�Պ!�I�n�*�c��58fD{�@sl@%���Y�_��&�����:��}�m�=z�M����0~%1��
�bmF���t[�Q��������a"�,���q(����P���v#b �l־kl�0e��k���7j��pԥ����F�>M,��Z[6mۈ�'�t"�$�\�
�	�M(�Az�L���� 	�8AJ㤃���Mn�Oş;k�@�!���f��hU���>?x@Z����?,=�E[]����OqΖ�	�D$x3 ��a�C��P��@Cn�t�md�J�ڠ>���#SfA�'�d��@_��#�SU !��A-h��8.��\\�rc��؍	��c�"#����$%�n�e�+d�x�����v�uў�+~�4M$��$��2IM�p+�����O�������쌛���g������Q�	9�O�%Id��\=��a9���C7�U��b}$*��d��ފ��	���c��-4^������:�qL�kpEh�1�sx���6����hC=�yݲ�\��z�5�}'���#N�ҝ�ؘ-"?�(�@�6�ҩ�mTR4:�Qޱ��9\t��������Ҧ	�������.h6��X�Rm��W�C���Iw�z55-�jT^�9C�I�<�E��Wq�z�����RK������r��e�(/�v��	���.`4�� $GǡB$�h(�bi��pN˭Q���,f,Ʋ�jd(ϝ�5�~���)�����g�G�f�� ��oJ�-\�0�^���1�<q�x��m���C��������=���ě��QH˄��
>��<O�ޓI����8P��P�)5,|�=^�m��L�\�x���u�G�IU0|cΘ���Zl,���АY�B����((���HРsF8��+�vr�
���*>X���zt���`60��~ �N�L�0ͽ�(�@sI0F�q�&�V����c"��c,/�h{L?��2V]��}�&���E)���P-8ˌ:�=Rl�'|�҈C�t�鴼UI��D�%F;�#�]z\P�����^�D1qL���<�J�z�L����ݴ�ڜ��[ʬ��ƻ~���^��Q%��>V�е�1ޟw�^>�6��D�Z�G�k�w�d���$�5R4 7_�Bb�QX?�6\��H�_�:~�W`��8; ��<h`���E�M��aM?7�[3i/���/`~7����T�a8���1׶�?F�п��u�E���Er��ñ@�3��i��uw��Dz1�{c�+��IL�^��P��8V,I*�=n
��U�!��/�b`��X19eݡ���o�$P��!���ߪ=D&}U�D�|�!-?X�|2�iy׸�WFDI�q 
�!���m��:e��Q�� 4��a氱���Wr��5A}u F�W���"9ʏ��h!#����J�xWI�%��6-8H��3c�gb�/ҿ�-�3ſ��<�o�M3�/�m�`�)؎�r<0�Ν�C��O�f���w#E�p�����d C[�=�Ue���|f�k�<�e�Q9�l����f`�ڼòs���z�W{ڄ��4{nO�Q?h}�`�P�-�������X��$�㥺I���{cn��sTp��έs͏��H���\���H��FĊ�<�q��R�J莹W��{D�>:�zsp�08�!@�MT�&��D��h��^�yۅ���0 �iZ����.���}��lnrMC�k2��Ӛr��VqUZ]E��sxď����y<��o�@�	���\��4�y��'lcK� �+פa�o�ײcSx��9]�`Ǒ����՗���I���L߽q�Y]���A���T�w�F���\ʈ�k*����k'+�=c�Z�p7��w11YU�G�ΚP�p-Ё\c�%�JU�Yy�T�m�S#�C�'��z�w4:\[
,��ȗb��R1��A!����	�M���_7)�&<z���V���:�%N�*����MK�>�$�gt�z�X_p��i������� Ksd��O+�=�Z|�𷂛�D��ϛ
N��x�&��*�ۣ�dx!�t��
�Q��z�A�����1��\�ҽ��,&�X�z��07��a�!(�r��#5ϸu���,�����i;�$�'�=�L,>��ڜA��S�gt��_����2ko���.�r<�A��ɬ��k����x��U���F{�B(�� �E=*.��7�1C��`�ָ�*x!�q�v��9t�X
�]:Q�o�����8������MY.�~-B6+-�]B؉�R/?7���Р3b:ĭ�(߇��*���Po�}o	W;�F����Q�rccA^��ldA��-~�I�gߕ�I�§���;^�W#�q:�/k��(R���Zk)^���+���(y�mTa�~��\O��~��ex��5�$�;rt���<�:�Z_~1v~C�kp���d�l����=���� 
�F��M��@���J��n��O�Yy����KH�2���*U-U#�I���JDuH�����=�J�O~�>�rB]�x*�# wja8\U�7����\z]�F��0i�V���"t!a~��_h���>$?����%nf-lY���l)ȶ,�?@��"2T�-r���=ݛ�K���y5߇��8uf(��śR�Ӗ���}5�1�K�a����4ʉ:	n���0U?�5�-k���o�p�����
+�䳎'��@kƈID�\�>���E�9f>R����N��пz���#i��5���ǈ;�� <��	�&��r��)�ŁM���^�{�b+�Zs~Aڼ������0��~m��~թ��|�s�sb������^�����َ'��ciLox���6�^u9tw帾������ ��#�;>j��t��b8@�!��Z��=�R��E=_�n�kɖ�lC�4��U��*����(<�o�Ԓ;y��b(/��&1�$�n��>���a�ٚ3��κN������7�Ԫ� �!�_�%�B�/h��x� �*UB; ��ƥ��P�l$�Q�(�`�L��'��?���`����&���+z�2k�`�3J�]�]��؎���`�|�àa�iNf6���|�#�=��GQ�j6@�N�h�h1��h|�=��5����L�p��N5fl|!~"�n�TJ��,��f���^,�U�^O2�B(�G]�.,��)�Q�d���W�ר\$vs�;�PC9�}o�gG�g:LՏ���Iַ���t~���4�����q��ĉae������i�C�쿓f �;Y aW6E�@L��cm���� ��j��S�q�,�BLg5����b�7Vr�2:��an�=��J�\m�-�,��.�p\��$XtW0>Sƞ3_�[k����>��[��G���A_kK7D��&�ʯg�)>��ǒ!{5��P�as���!�~�8�s�2q0y�\]/��;i�}V�X��xIf��~qW��j��>��w�J���?7���-�ѓh),�h�;�1	�� )����`T�)���kO�g�C���}4�3��O
�'�<��,�2�: �_]6Ǒ;�߇�=�%�e�a[�����&�YU&c��	t�T�Pϑ�ŕ��&���h�X��2�<��X��R�vD쉂���r�Ś�=�R�bQ�^A�u�����J�]��s)�n�M�Ld#^��"FC�5T^���۟��Z��Ă�W�Z�Ԑ� ^L3t�֘nv5r�K_Z�ׄ5���
�(�ϒ����Zc�����:�J-�ͬ}ή���#ws�������`!���}�|�4[�X�����9���Y�k^	唖�w�"@�r��_��Y}��F�]r��*���5 G���Q���	Z�ҹ���0��S�Zs	WT]+%\�y�Ww%�[����sU���e��N����F|�g��� WO��qa�����jc@�?6/R�N]��CK���;������F��/p�X��	��Ŝ�΁�%�(���FO�}��!�_�,�[P�b���60�*4߉���;��F<Fs+>�>o�-�5p�8���(xgR��-�j�Xc����������L��+S�l���4UL���vr?ȕ��Y�w�=�*�0Uh��)q�!S�;"	?����=\9����!�$v�pO�-($�V�s^ �}�rc��1��z:N9�q@`��u�U~�F����]8�O(�PP3�y��RoN"/.��N���ha���2=��m�� I�J~ �=y��\�"� �M�N���J4�XN�D��ZB5������l}8P�9���'�+����W�K<��vw�h�
Zh��>���X���;��V����_���gm{#�t ЕZf�s#��lK��P�%(�B�0�e�í:/^x���G�uK����W�K
ؑj��'��\��r�:J��!��L0���'L��L����&�X�t�z{���H ���8�%��@h�L�{.f@�>�� =H�Ұ/�~u!
q�h�սi�>y#�N���a������-�I������ ��bV֍�F����&z�?Xg���jC������V���2����TČ�Yfa�a�T�����	x����+�C?���4�`�rk ��$���6n��e�{���8�إ\�|�p	���(enݦ[DuT瘧rK����E�a�p��4�rGn�Z1%dJ�_(g�Z��:��+���k��?^W�Z�d$�ު/���-:ٺo�!&D��ӆ��Z�c��J���i}j���6&��j���+�"�NL�(-�@,L���~���Q�~�|_Z"��ku��7����N�=oxJŉR��GNjD�f&T�L����ޮ�-Uao�ӕu=�F�^>7i���H-��� D�i�Q��sT�x������V(�=�$zmdM��JG�9��>���>b�Y����F�18����-Lc���z�:)�k+UUE٤H�t:�C�p��N�>^���˒�lF�Ã9�R.�%��2[,Y@[��$���1�������^T�H�(vM#+K]�*d�Yᒾ�hhS����C�FgL��Q&y	h��V��Lv�]G���nپ��)�%����Q$�7 >F����`�����'�5��Ed��Aˢg��0��{ҧã��I��8������64a᧙�eT��B'�: �,��bj۳��)���&������l����\U��PB)��6�d����5��rD�/G��u�n�	sor�"��5A[/ͣO;�w�ն5�L��4כlox���������Hܡ���y��"�	"#V��B}���8�f��c�M512U0ʘ���Fo"o����.�A����	�uU+���i��6ǩN.b��`�nw� �ь�FC�+�x�����[UoQ,K����q%��G���si���.�釥������p���G,g	����O�"�%%��U���FQ����}S�90�k����~7�x����1\c����UD4z�p��LP��@e׽��ֹ ��T��ĸ�����C�xP��H�,i�-7��-��p�'��w�g��ÎK̀�z��n��N��g�4�6ݨd�ㅣnd��Z�(�;��D\"o��ߚ�X�-o3�Q��e���j��>dq��Z;jgW�S��;����7d����s|��v�Ԣ'	ޯF�(�3M�B�;�\�B�Z՟>�TdW���Pn��jۿ�k���e�x��)�˖6Ѵ)#�������:��7k.�@ܧ�8�玭�(,�kxgu8�s�H=d�F��o'����I<p�Ш�\T{;Y�Qy��x�An3 )� �����~a�e��A*]��]��)^'��-�Z�� ,���#+ �d=�~��PǸ!���Q�SE��#�|OK�_������	��(d���#&I P?�<����q�p��S�~�L �� "�N�>�V��=:�<�C`���`�-�=b-���B)�3��]�p�еD�E+�t�F?��U���Ydɡۖ��ʑ��j�c���x�$���0Rh����T%��������쳥(�}#���5�;�c� |�OC�#Ā�����2��j�P����L!0�+tL��%�9�Ԑ9mZ{��&ib�:�-o�b�X�G��t�����D\9 b8���T�mܗ�>`Y�a�F��tfh�xd@�$	�~���<[}�]jc.���3�Bo��,~�3������b�)b]dS��à({���w�-$�@�$����bf ������3q+�hՕ$h�q}m���P�_��[\�~��~�[JK�m�1�,d
e�Z���$��Cw�����_T��bH0��e؄ݵ��tܑ�>�6<�2hNe��Z�j�$�!���q���7���  	��d��)N��z�"B��KK��̚	E^�ٔk�Q�X���q`����B_���,��H��wѨ��=��X~�Wh�!I�G�������8m<���f��o����2k�eW����D��"��<t�!p?ϔ:�q�t9�½�����~�	��4q���]��d�Q.ĭ��� /���q;�� K���cw��T\
��X��).�`���t��5�C��R�
�Ճ�0�Z?�H"�9#@��:B�Hob0Pw��C� y[�my���g�B��t䝣8}��5�@}�:㬬F�{�u�F�L��Qzi�|��9w�Q��{f*�ب�R7f�(�5;�,��*{*�x�����&�=\�qdl|�,3@N��V��͍�L��b�I�����L�ߏI(ki�Sx��6DHiEo.M�/��g&���x����+��X������	�~빰��c�C�:���}RG��7��׋�~�[���B��اϫ��pʨ}'�۵��W����!~�Ga%��立r4�%�F��K����	˰N)�sļi��.�RQ�N��L�<

��6��j�u�Z-:0Y���������k��CP���*���
̪1g�m�T�H��&�����T���)�D�C	��ؽ�^�4����m�5�����8e�8�Ez`
d�Tp+�,���e ��)YK��v�E�~T�֕6��^�2mW=?�+-�O��h=b��?	(��2�����:vl+�μ�,9����+"�0�����zS6օn3�3�؜�]k�3I���1*���V��R�7@�R8�˫H1��U��q�1	�^�����">=�w\�peC�n��%�؊��\P��"�]�p����k q�A;{bQ�!4!�	r���y�3H��u�k�և�E%=��@�����R Wm]Q7)drx�~J�^S��J�ܞ	�tI>�y��9z�M�}>'tP�v�9���-Axu��5|�ik6�բ�����o��,�R❵�V��t��rm4��:ia�m�z���:a�(��� 0�sJ��P8C\> �]�W")��g̈c�?T'MtW߾������ᡯ�-������ع�P���$<��j`-<[{�O�僋(?�,���`	|]V4@iE���v�輸�MXK~��pB�y�섀%q8�Bgn��7&�ݕYD����`���U�<��H��pl���c]D��1��}i���VL2IMTI���M��� �}��~�]�-�s��� Zpӷ��ؘ�ƉL޵�n�(�:�n�;EM�R�� #\�z������jpU{����]�2��t�#�����(,�%��s'�MwK��GA=B��|}b6�
��y.L��e������%�Hl��񤧄�{(�g�ʑ�4������ܩ"�r�p�w��u�;�',��u�"��d����T�y�������P-��n�ja ���/����*����d��85~�����k��K�3��$�o����o4��o <�M"�P�H� �+Fq	<D��!<7i�������/I�T#3����(]E)�)��â�Mt��� y�3�r�*�@��L3v~ј B��L��z{	�=�KsW�l�!>�D[�ڢm{��rwvH�Ӂ����ψ�1�k��C�z���?�������1L���T���#>3�'�!B��i����Ɛ�ya��1o�]e9ȵ����)�u4��0xg ��F0|2�>�$�a?=j�Q"�
`���k�=ț�#i���ϑp˻3��zW���~WL���1�_�^����'�Y�{� _nV� ��!�����o8L������$W\L�����_�ÏY Dh�9J{�IX���Oi�z� *�ZcY���M�d�!�7Iyr0�Ty���C�|%(��0�*��xERS��O�e9����އ�Q�nt!������qd�:�܏���#��,�x?]K���w��w^����^���u����5�C5y%d��� �1�
0x�:c� ��Zk�vO��
��D�N�
s:�	L�+L����Nz�(�n���}�3���21�:�#�x�)ۧY�6@RE+$�9�Y�/$٦cv�B��%x��}�KI�7�[����`L���� �Z���Y�� �k����7S�4����D�=v7~��\_z��v�[X�"�t��e����S~�J��ԇ�O�s�wJ�k����|�6��$�n�M��}o*/C#�!���%T��5��� �!��k%C[V����ʾ��Ó���xH<�����,�܁���猧M��W'N�H�(��m.�Ê�#+��(K�XRв��-]a�l���)ZO�#��0#�F�����N��4�re�_��)�Z9��ِ6�Ý{έ%h�Q��$��]�+W��CS��Fȏ�5�M���h�_��[�h�(Je���޹�I�!Pe���0�v��@?)���hB��fV�z����^T͗�Z�*\�}�����:ߨ{t�Af>T��y�ܹ�Y������j��j�3r2�h!�k~^��\T(�[p2�l�w�{�6��#�����C�W�/Uuu�=W�8S�]�V�l��W�\Uq$��6~.��~�iը8����K}�)�a���^��W?g�^�}E�~#0�?�yK��B3T����b�+�⺰Ŀ����PEB�����SicV��3���U��RӶ��x	���&�2XΒ]�D�;�����(�B��0�=-��~�ؘe���.���sU�uNBWѽȨ�I���?�`�iM/ �^��}�``eu�[&�bU�k|���4Fqeӭ�/��TD��;+y�H��j�I�&��̬���р�ѯ�j���1si�W4�>6-|B��Y�<c"i�G�#k�=��[�je<�L-�_��K �2H��9����^{[T�B8Z�h�ѱFFY�ӛ�6*�^ˮ����2x����]�g��ܨ(�T��0��Z/�XJ�;?HoÒ��D�)BX������f�ʊ���j�"(8�Y6V�����:���k��BBU�b����l�(��Ų�.�T���S�qb����V�3��m�(!�z.PgLH^�������;�O�s��CL|�*o����m�7��z��S�5�2����<�a������)��F�P�S�6��MC5�7Dv�d#���-\��tU�Y5�&P�	��zń��e��|�9���se1.�W���}Ĭ��g��y
S,l���"�/������$Zy����ߤ�E$>�$j�)��n2�&ρXk�;�}�&�b�h���ae����f����XRٴ�I�49����t:�q��j�ao���#�kB�� '���u�L.�ҧ�`+�N�A����\hSyb�ּ&�����:���Q�1�ZolzԾu���"a�=�>�B-�ho��� 7�c�v�	9�S���j<�����U��k�D�ցH6�<���@<����}u���g�;�+�&�)�`nӾӰ���N.k�&��gu�_�]�~	���Z�^o7��n]�;��$y�G�\|"Ic���?��� �?H)[(K��a��PY.F��%�-����k�(O��A2��J�s�>��h3�#kG��6d-�A�.��C	p
���==�첍f�9!]�F��v}*V.�*Y���t	ւ�GwXal�scb�2�a��YH�Z��� n\��0j��b^�^.�݈7����������F
u5H� ��[�i�M3�kڅ�m�;�ĝ�mKUYi���f� �^-��	��7�s������.���Od���W1���>��a1��]8��
�O���n3y`Fpr�w�a��k����Z�r�����U�طr-�}�-zG��_���k�= �:�1�)	�H4��ը��?�m�d!�p��?�^��u��Fxo�|:��=���T�����Ԗ�ɺ��s��nz��F7~�!e�ڴ����6 ғo��$�#�`�<���n^ �ե�o r�.�_�E�y b�`�L��(�ѱگT�)���d�N��
0�cׯ����O�"�������"�bEDsi��s#�l_E�)#�"�;�%�^)��f(�J�&P� �@�99�;��:Z=��éx/D�ȓ��ܲ���)��I:@>MO�Rr��6�l~�>t��������+?��(Íɾ"�珯JGr�nY���p�:��|�ě����.�8DE��JŲ���p�J����Hɡ�f���c����6�8M����$f�F�����q��kZME��d�yV�2 8�a;�flC���
Mjy�߽V8 2��1���@$�ۨj/+ͪ�������9N�.1�BpbI���	GpEj?��`RZW���PZ�n�������z���F�����u���ʡw��~s�Y�N���5Ɓߗ(Of�)��j{����p�P��1$���W����MH�9����"֨���q�� �e&J��-1��8Yw��a�"ľ��{�T~*k����j��ƺ����х	r�1��ŗ�M�iY+���}��$��=������$�R��x	�.\���l:#0%��υ��ۧZ���������i.�x�a
�⚿/�A�ٖH�I,�Y)�����0 �/%z�=L�'����f2��~�J�}�10M�Q��z��u��I�>ݥ"��U��7}KVx�0ے���+�z}�<�Qt���_�v&����'}˘���h$1��-�.w����v���/������"/��s�?��L�����Aa`���R���v���1�������hG��v�U���r�|��\����qi3�.7�?���%p�����m&r�*[D�� ��ͭ����ON-B�J�]R�[��=�s%3T�O0������t�0���'��+N�f�O��MjM�Y���iY-���7���v%A�xןQ����4^�/��O�hN��"g-ҩô��`;F���NL(S��z�s�a>u���xO=������k�Eca���?�;k�7�<
b�.�)�i��ԻO�vy�EG��g�lെ�-B�� D��3��ܙ~�ͻ���ڜ}@�<8�O7��rʉIe�OGEE%J�x]~��|�QցAtQ98�7����?����/����ԯ�!B�֠�ե3�zQ��g�I|�i7�^na��d� YՍ�*J��§�P�ʓ;��i�]���썣��5�p��F��m�fD;�~�[ִ���Nl#��F�+���{i�	O�м�Z8n��{�9�o#��r��4pLt�����FA��#� ��Tf�g&$Y	^ag1�=����f�h��/�5%�Q�6�,���R����`��X�+I�ѽ{yHCV8�B�B]qo��	�j���Wߞ��g�'��Bh�L�4��_�����3���"�E`#o��w�#[|U��1[�f��
O�!��.����b�g%m��l� ��M�7���%�\�oh�6f���O��4��E�^�� j$r����J�_+�v�&wj�{N��R�0��ȱG� C���/��o�{1	�٤U8	�*hټϡ���4�./.ZD���|\b�A�*��_`Jq�p�ӣ�+�s���\GIp�#>�k��zd���;&�	չo�\2�?��L4�ہ��G�#�"�0:�JD��S�G����f�(�0H��� r����Neh/��*8���]�*+V���;�:��`B���n����v��P.�P�m�f�u���D@f �Lþ��� ��|�Dw߸�U����i�L�|�XG��Ckp
(�$�P��n����S�:�,�N��ؽj;^�"Q����[7��͜��m�u��a��2"�U���f&`�D�Ǹ�_��'i,X�F���x�9���j2�f6�[@E2o�#�:�ퟏQF"
%�P4�t�/c�=�5qB�X1��Yl-���0��@�	m�Zn�)�G��=,����I
�Ru��!>�&��$�K��D���]N�ٵdB� =]��e��c���gVf��{s��nn�VYG��ʹ�������[Ј���M{f8���q������bK{(.b=��d��]�ڟ��Հj]�uV ��Y-��%f9�o�B@6�7Xۦ ��8�oI�IȮ�x���eJ�qi�%t��0�\���lԕD/ɺ�FR9,P#F�Mϡa�$��`o���L��J�wݓ�	Jc惠�.7��4MN!N,S�)V|����n�W��^*���~_xNҳ�l�	H�A������mo��_���U�X��Jz?��W��|��]:k~�C[�	U������{��I~7v��A�PU������T@5��f�h��/�jj2п(-񧅒aM��c�_*Ég<b|ۘz���EC��A�O�Mm����}�	��Fa��O�?���]hٷ*��2�'��\��Ý�b�3��a�.��ȵ4�'�.�21���R(G"��-$d7� �k!n�-�L,O���Iwý��-lc�R
c/�܅����}m����2�Z��p$Yf����h|��z|�LR��M�!�v�1����T�ڽ�>̹�(�a����L�y(�Mw/vƯ�j����Y���~B �?���Ӓ�q"���X�y3񱙴S�=3�;r�s�"J�C��M^bQ�K`?)~R7\�v���Y��3����@�,��qt��ƴ�C��i��÷�7��gr>�gʵ��h�����`��z�0~/@05�/;[`�
S�^s�D�J�����5y�p���X �o߆���F�Ԁ�%�tÔ����q'.����_Z�M����V�>������ߺ�Y��;T�!�}<�7<8��`j`�H�a�Y��t1�*8�t���7�۹��[��7G3��u��,�� *z�tqY���zb0��`~�!1Qxu��ݨ7��D9L:8a�n�K�D�U_���^�(�@���c�o��'핰��9�^���Mm�z�S=2���4�f:�fHA�#��Me���pϾ���!	��$�S[������Z�:�z���ƛY��bp��ơ_JA��.�U��8 ��#�>SÔ��j'52L�9)@�`&P��Rʧ�Լ���`Y	&�P �N#u��2�H��1�ʶ4��ˮN�x�sob0Dox-V�A�ѫ�n�A�R<�A4��3���i�G����%�&���lR��|h�P��(�T.����Y�ud>=_����=4���3n�?6s`]3�N��NK*A�}{kDmqi�����s'�K&	��uX2�<�Ǫ\�����n�»"W#�"�����4�ުX�o�e����L�hoc
�9�"轚!�k&�����q2�y"���0�vRw@#���|*v�S"����1˵��� ����� ���g5�w�*�ET.�U�JX�G��
��ƚ���A�P'\d�	ж$����4�ַ�J�n0Uʅ'�L���M�7���w=�'��)zӴ
�^��zߤ^]Յ�I/��c���՟@���F�|K�&k[i>�#ЂB�?�f��/dc��'�q��=	�깖�x7%q�E 
��+����o���Ԁ����C;����WO�KK�݋|�fB	�2͑���=;�to3� �rV��|�OLf#T�J��x�>-ȬaKmn��Ռnc��	&��+1r��L�ߢ���\��s�?�<�A"�W}�?7�A,�5���ic7��&��/�i��9kR�g�Ywk<�io̰U��y�� L镗���:>+�X��1�C�h��s܈<n��,�Ρ`(ShI��Qt���*ͪ���U���\>�*"�8}@��z�
�4n]����sJ�W���upA�H�!��r�v��JԴ�Us(u�r�+[y�ۉ�|���aJ����=���ٚ`O�d��s���l�����0��?G���=��Y����L_��w�u&�X���������d�Ӄ�ґ�����w��b=*������L[.����>��o�  �:-)�tb3��ur�U�7�| T�_�9�eH%�z��h�p`�}ρ��h�%A� P�X�4�YL�[�x���0;�з�V�uo}���)L�d�4!
{�m2��bJ-9��5��#�`��?$���5�����Qy]��gSUϚ��� �˹�6EtHƀ)~�ׯ������s�h��T��Zgi=�O�
C1�[�K���d�W���	6�˽��h�;�Y�&�h	�I� �U�(-�0B2��ƹ�V"c�J��q5{��1Q�?]B���\/ggw-7.N#γ�2�-E�1�_g���^aVa/ĥ�<X���v���p�_2[����l�/O$\�'
�X|�ͱe)��3�绗�c=X��֞��|wKz���5/�ڙ������Ǖ���w�����UI~��q�8Q���Y�zfA�
-ԕ�3t m5ٕNG=7?R�5�J6)�$�,�)��HWe8�����q��)�Gyp��S���ˠ���c^k�7*����i�h�W��sJ�fN/Jز9�o��,-l�!?�� =~pA�})�zH��SJWo�+M�F O�q�/NYץ],�ڽKG̑'���A.P�N�h`$qu�F�=��ᶈq�Y&e��)�;����H�z��y^f�6��ҿ�. i�+�No&�=�
�ub��هڸ�?�����^Py�]������&���0;7��=A��/$5j�i����W��RrO���ו�3D?�]R&ᢿ���˯��?��/t%�I$��d#�i�`�=��߭n��*�Ҫd6�7[��G��h:
S��l���h�e�U�i��/�'{e��`ᗖJKU�A_ĭ��~���j56�^H'�,�'�\f0i_4�p8~!<��;�1���I�K���HT�V\�A�]�b�H�fn�6�+��3E�YG��#J�R(A(>?"��F�rI�j>�߲�RSy��Z&����6���]-,����ZOu��5�|q���̂q8A�����j�z�a���ҩ}��gS~���j��o��q�ֻ{Cz\�e��=��=�����[+e2�W��t�8��lqҜ���4�筲5����WxR$�uȐ�@S�.��̃f�U�1ҽb:ʧ����L��Z
��Oq?�Q~d�F���6���LKͥ��jZ��� �.�J)���29;�볒���C ����,;��GĊN��NE���4�&��&�d�ޭ�d!R`|�8�N(	�I��G��5�E�0?R�v��D�O��,���\�ȩe?hV���xBbQ���T+�qN�av��ڑ�Ƽ�c`pQh�ێjB&j�(�\t��;��Ѯ�Ɯ��=@���v�/�?û�K��܏7��t�\x��#n.OL+b05�ßȆl�%<���H2Z��&[%��)��\1du���>��`��L�f�P�\o���	��~ٺ��F�w�Woo���X�26P'g���x��4$��=j$�P�,�9��r"�מzr鄣��Dex7���<�&e@�]����� ������݅f�J��:sL;A�U\��ǝ�DX�N}>H@�� ��j��� ���c9󱪌UM�;�A�h4}�J��4��y�Ĝ��-�s�����Օ�YWc�N��V�\������u�w7��WZ�ɔ_�98viϝ��1$����e@h����_#T5Pa+�2��Ɣzw<͕�e���U�ӱey�u��|c�K
�n�y�	!���Р�] K�#X�
�д.�M����`<��\��,�=ԐU�ѳ������t�:C�t�ޡ!�9CJ��5L�g��%IX޳9>d+g�tSe�j8��&�f�͢�����I����QDJ�I,�=}�|�"LU3�t����ӝ9�sW�O�*${Ea�5B���j-��2{<� Ӿ��IEg6���� �n�1F%e��"H���|�1����Vfl�kL�Xc�-��'�Z�ǝ:�XH����L-ݢMϲ�r�k0�����X�<���_�&���%�B��'I�Аː�C�P�����Ȋd��
'�'^\���m��Az�<T�Â���;"�����.�B/�l�&�9oH�gXSiQ���D1�P$0�:
�"_�.��:�B�*��s�����`&޺�|{�����f��c�X䂜l�H�ƹ.����S�����i1�E���{I�$X$��$�9�,����=�v������mon9��8Gi����x�IE�z��[K�9���Tڸ/t�|�l��ӾF���eU+M�;��(�2P1/њ�k�sˆ�Q�;�x��p�"P�b2jȁ(^�I���YR��ڪG�#�߂�6�y�L�xղҘ�0۩6��]hW_�<�OW�Ͻɛ��gP�O�=��ҩ���/:�D���]8�,&<�Ff;��flȤ�gW�)�Lac�C��U���i�1�;}]PAO�!�B���\OL�#�3_�s���d�ߴA�⾦�b�7 
K8:8���C�\���Q�D��M���ڡF���� )c
3���""Gӕ#����Z�^Z��<��$�|))�s�����L�K�hL�N�;U[V(d�w�W�?dT"�-���}�M�Z�����
%lp�
����,�&2�f�'�/ss^��)m�گ�2���FB�灶�S]�����w?����\=��6���՟sI����L�E~r��m��J�C������>t\�׎���^�F������:ٔ�6�K(7�㠃Z��Ѧ~	UI�cv��j�׌����øW�J���]�u�^�[���O����~6�K��B��
a�^�F:����/��S��/+��3R:��E��1zZҗ�}� Έ��˒�bD�;*�7�M�Qpٽ�1>�f�7�̑������!
�~��%�&��sB�&��w<�5֕յ�(��+�O���ȯD�U��ڪ�Y�	 ��hL�lYCl��������� ����_}`�.Fm���0��;��y�6�ʜ�%���rZ���Cu�/�^���±�����g��Z&�b�$.d�	�_���s�I����z��}ö�A%�ԃ�pV�1�D���ybb���"�%4�EK�����5��NҾ�a���:V�$��;����O��ox�rT4�9���8'F�utԾv6
rd�Ϋ���EFU�����E���G7�Ph�fu���&f���"���T[��-U~�Z��;5]�:9��*������cVP �� �/6ט���	���/�-~*�X	}�*m��x�&gez�3�z�u�t�Wa��?� i�>q^�
\$������]���y�ɾ�� ~�ʭoA��;1Β��'ec�3�g*��LUǏ�zō
Ⱥ	݂�����]W>�ˁ�)9��z����Ȣ�	���bHk�4��p=���`�i
�5��z��O�]���l�5y�����l���4;}%�:D���o���p7ﺽO����(�[�!cq1�B�é�yK݆^Њ��R��9��=3(�J���ōѪ�	*�r�C^�Y ���ŕ���y��w�k��|�|]�V��1����{�
����f��b���q�C��'�]�Z
��-gpਧJ�g�&C���Y�jz���"�[�ֻ'��MR��	�wYmR��_<���3�M��v=(|��`���չ��l��;!�
����{�S[�N8`S�ht�D��'0X+�њ��S�ʧ{Ɗ*q~H����Df��쿧-�XP��K3�:��/IKv��I�20�۵�/n�|�*�>�Ӏ���[���ʋ���f�v��;��G�Rx3@ɇX��?���j��������ZR��4�[���?���9�*��Z�HvJ�H�O9:�Щ&��;VB�X� ��(DR�LiA8z+��x��~ֈ់���W���p�:�֢Π�=;����M\ˠ�1w֌tcL����3��}Ǵ�u`���S�T@!ߚ�.�"��0�|S���W���_]bRZF-S�(��K9=�iؔ�N���rLWmm�>��Yv��%{��9�:��k(n+������ �qD�/�5H.X�\}�����"~���"�g��O�A�wRqhE�lp�����&o�Cb7���ufL;�y��D�[(o�c)EEl(o��7y�%t*���� �h JF~�@�)Q�cwӤ`��-�#�O..��R����;y��Gգ�9t<��	h��@I�F�^/!L/7:c�v��7^�K@���6�^���X�LJ���7�`��b�%ý�E�:JW��T���L����i~��ֺ�d�Gi�E~���w�Y���L���JK�~2J�
]�c��q~�X�pFo����8*E�bF�>{n��2ѧ��u[��d{�e*U��gCG��ee	@za�t����:bfa��G�+��XE��Zm��}.�".QXQh��v��4�լ�9e����D1H�AڏlR�("���EV�A��pa`�v��A��w���d�q���L�X3�M�B����*�L<�k^M�Su�۪���M�)��0�٫�ǟTU�_��\Zt3��Xn�*q2��/~A)qRs��tC(��x6w�.rF2dީ���{�A!�3ڶ;M�5�s�3N�e���o��`D��5:��%�Q8�+�=��N+g7)^x�X��L�[��^YVwP׬vh�Ė�Xѥ�Ņ�	lbL�Z��*es�B��%
)�;O{�m;�wjN��&u�jk!66�����4��� �b28ĝ���S�ѱ9܁�&�&Ղ�0�}bh��A���miiȭΙ�(�>֎��u�j�nӜ/�N�0OC�ۦ������7�'pP�_tq��1���ph%5PZ�U�k<A���$@���P>"AT�d�}��*v�^�R:�l�s [^��[�_�9�*q@mR�����[	7W4�"�VFq�1��~�����|�%�T��	��/��|����2�n���F�oG$��C�pS�J���C%��ԧ@��?�MrD(v�L|{����������=i�?X�҃
.�8��g�z���>?GF&������j��ֲ��8[=�M�+��f��ƿIb�WV<��M�J�:V,��:g�8طp�#P31��*��$�ky5����3㡛�2��p�U��7~e��>���ݞ�Eͨa��
dZ�~DE/L�X�VԼ1�FI��GՅ�%����,�&��F_:��n�۬ڍ`h�d��E�P`-a�>�ϗ:�]��a������t�p1�n+��/ea�����%Cg�U-� �5tc���%�5���B](�7�_F��|���}<��0��Ӥ���O��ϙܜ���̶XM/=RόY/��R���3Y���Puu�HJ�?}QЌ��	�L�Q����Sa~��6}���xfc��Q�^��ҿ�txL7�Z��H7��C�2��ۉ{���OW�p.��c�)N��T5@�U"����@'͇J���	w�u�><��]Z	���c�]�b�J��j �������羱�+�?s�7�r��L����s�9FЂ�.�����/�b�1�3��#t]������tq͵"��:AfR��P�4�hn���0X`�����yaӑd:���̰rX�V�������N�����{q~@�*2�~����ّu�G�6�*�H�~ˡ��� ��JJ�Y�-3/O����{�ї�m�Q=�v5�� ϓ�s`�+C_�Vh%:�܄*�:�G�?U�`+ߣ�VK�XFe�Rr�)��$�{~�dz�c�&`ܹ�pV���V�L~i<�R�l�%�C��^�4��GSI�f�?��
W&���2	#�����V���J�~.���P'|Z������.~�;}r%�8��-U$��a^��I_�ONoQ��WwF���E��c[�!�l!�kdT�^�>�k�9����bA~`I���.����Ʌ\p���`�Rv�|�(�����h˴��q�5#�u����<:��wTu�z+ "٦/A�(�4�R�/7������e?Zh�aX���>*�����W>�<���AǼrS���:OI��P�̐��р~�"���{�q:�� �X�Kk<O=�R��Nc}���!RE8b����@��#�({+�:Ѩb�U�c���]�Nk������Z���Ku��/��L���c�8��$��T��H�s�k��q��k|f��ʑ��u��o���/�>���r�\��C
6�O��8��#d�B	Lrv��&�A+3�QJ-G7ٚ"�"�̸��=�\i
0>i��4�z�/v�����9�N���x&?a��cI��>F�;�"^��S�pͻ��6ۛ���aE����W���R�}����
����qg��Jc_������q^���8�\ۡ�Qxj��K�pÙ K0c�B *b���6���vĨ��v�������X�i�_�`&h�N@9J�t����~���b�:���}2�q�x�ۦ_վ���S}hR����* �/g�n�G6�Y�����>��bӭM�dC��q�����"����|97��qc$��~3�{�_)�<F�&�/;�<��f��}��g�.�����>����9w�fB:-7���s���Ge�)ѩ���؟}过��C���,r�B^�R�k�(�\��@F_2�8��&�� �A�|SmU;�5��3i
���a���.ʑ�,Q4�TtR� �S���_�UZ{Z�5a?r��d�i��~�ֲuN��GS5T���/�*��Ju�|��{8�7a�}ن�,�d;-��`!�=ݍ����01���C�t�0���BH�Q��Nl�����j@� l����i�<��wE�/̎m4��gou�+gy>F��5r?�v���_�3��u�ڒN��DCŰ7���T�-whW�SȦ�TA�J�5���4.����О���c��$���^���l_��Y'�ؿ���3ʇ��a�����{SUoY�"߳e�NCM}�X~w��C��&A��.!˭ɥU�4��ua�3��������i��������BL85�1d��hgQ���V����C����.98]+Xa�v�h3c�H�a���O\v���Ŵ�4��\�=�)�:�P�9K���p��n�夵�a�=�&o�ݪ�{=�����XB���=�Pm���D-eK~otY,�#Eb��U���y�R���%IE�(�#7��{�� ����Z8���
rQ����v��ä�}N^��ަ��E��&��kޕ�R�a��+�po����Q�5pF���7�?}�
~G��(��N��cBꂗS��s�L��SG�h�� ��w�U�@�_d�*�^\ǣ+�^ f��4��^����!3�m��8��fs�`����E=�a���������A�`��pI�^ܘl�t�1�tPU&_���2tZ�f�^uv|��^X��H)F҄�*�m�ĥ����I��RF`��?$�����ɧ
��Ԯ�4�f�;E�7���D��f}�9{=�'�Y�U���:?�k�2邜w�cMc�>l��`���U�֞M�9BF�o9Ѵ�vx@�X!�Ly������q2�Ll��>��ݛSh\��+)e����#���	���f�y�:�U�o�X��S�q��a�.�gߡ��
�*٫&m�28��'�ɱB0�!a�/�Ls�>0V�]�4�/�*�1=R�G�Jʴv�zK7�XmM���O�D[�����M'�;�f �j�H0�?}�j�ß����d�A��`#��QR:5���� 7�v÷2`��rǰUa���gvai�
]7����LԳ'=΄V3Vх�h���\Ɠ�{�q��_�k!�q��m�F���n�tX��c�9�<��)��uc
QU��Cz��"�g��ҭ��� )5lr[O7$���nx)�	1H�4���Ԇ�B-�j�B�9U�T�����	Bb�-0G؋�j�UMxV�/ҩ��Q�0WX�׎�d��|�Xp��#���h�!/�u�w����҃�؛ǟ��|be6����l&��L�9���I�t8W�8��ΫRS�$�S�r�䁿��͊Fr���&>T�B�S�%��I�y���;�5�X�!WW��{�w�C7dJElG������9b(J!����x��߷�Չm��f�a���-Tx���v�t�\�!t�X�g�"����Yu��CT .ǭ8UAu<��ءK�w�>l����#�̽���/��((:lSq��'Q�:�L�~H�ܾ�2�z�i�>+q"��!�+�9�F��zΙ*�� .�g-^�l����#�C@�jٯ�1s��=4`�t�����f Z�k�x� �#`�g=�^'[<�%��	O���&��C�zI�U� 4G�?�k�+��u\��
�jC���f��7�=��=��C�?����g�p�:�����d��P��{@��E.E�/B2��Wr�h���0	����$6`�1�HJó��?Uf�؀��_!���/K�"qQ�D>���#m�2d�ԋ��?B�e�GD#A��fm����fF���:ބIٙФsl\�m�'�s�t4����w�*����!uy #�	w�`����9X�ѩk �Uu�;�� ��G�1���q��w�,\κ2��.����``T�A��㻚_~;~��O��3y��q؏�@��Ι�*"�K:n�v�X�� �г����n��C��Rx6$���:m�HKj?q}
��`��@YCN9��T��Х�^���T�[���96PF�0),�����"x _8����U�id��E��in�	�фュ��>�6����i|~4��뒂
�F4��A?�##�G	<ٸZU�]r;�]�)!���&��o�V�T˓͛b��z���J�a�i�g>\��Ȓ�1H�m$,*��ԟ�T�0n�f��Y�C(�?	�
ϭ�=��v��\cx���w1�ٓܣ�ҍ�,�<�"D�GB�)a��;jZ�����1�O��Ĉde�p���/*^v��#^�����1G$!
1ac�B��c`&>�t'tD�4�?>=�mK�{���ʄ�o���q�4�F�Z��ʞĐ�)$)$�W��Ð�l����a�ʋ2�7��V�d�x{穤H�ӆ�,�3�s��]ޥr�byt��i���zr��O��E/���I��"�s��}��8[tWw�?�{g������|�{Qp�łeĠ? 	���_�ƻ��B��>����&NmT����i�|<�h�oN73��V�ِ]������r��	51��-���w���T>�)�0�S5\�����{
;\l�م��xҡ)��S���ū���R�d_�7M�P5X�%��5��	^7�ӰrP]؀<t�r3&p���&ǖ��v��� �B���C��W'@ϜO��=~�LC�Aw�Fz�\�����h-���#pO��_��INT��ã��2q�	����e�����LMr1V}O���Jx�C���$��T�V�!w�jS�lP�95��a�2o\V��'������R����;5H ��j ��~���'2���⮹�Y,;��ߡt�5�o.�|&�BrH���mT�lE[�������	�ݵ~� 8p�w#�-�G3���l`,m��C0VGQ>*�9	�ɪ	}t�cuV�F�'�>�ka?��Ys�����Ws ��S�R�E%�6Sp�h��b�"RC6��o	�>W!��_]D2����s0S^sD�HjG��	�z��D�"�QB�k�鬜��4<���'��wP�/�3r���}�JZ}!�	�*��-[vI���y�ǹ"�㺊$&�7B��w��:�TZ`�r�Q����ۉ���H�K�BB�?�	H�� h��=����$��`�z_XA��W'�h��{�#e��5#��"�;	�~�^�/����$�I�R���DP�	a�Z��rPz��אd�e~/y�gv��S�I��X���Yi�����F���J-=D &�n�^�\�=�Xq�蘆���0�lgڎң�J?:S�2Pf�U�\�b���2���<{'��.=_J\5W�;��Z���'�h�ՠ5�V$�S�����;h3�Yyv�"�GnH���=�fs��ƃR���t%��%V%wDȲ����,=���8b�UF��F���wr�!>~gB��E;�b��);u���A@o(T�xx���U����Vseg�Tg�X�ř&I�ؑ�kk�_&9�S����(�)�K1*���$c����{��L/��A�C�D�ұ�V�P��2�8���)z�W�	�����M߷�J�_�%0��j�oզ�C�]Ѕ�R7��<r]�.,v�#�5�֣#Uf�����,6�nC�I`�~q#�xԀˢ��~����5Ʌ0;$�;$��R�|���^{N{�C���[�N@I7���n���# ���^�6J+s{�Wi}~L�� �������y�[.��E�?$U��fW&�ў=�6�瀤�@���GB��l?v��{���X�X1F�\���̿F��'�6��;���7g4�!�|�������)���:?rl�gY� ��D&_�����#��� !���R��,�Ԧ��|Du��e+���<|�W8�#���M�N%ET�Ǘ�2�>1��ÿ�cvh���z�����S_�9��k\hM��Q�p[�3��*�����X���Fl��{��g����n�A��+s~�R��n�t�I��c�bE!|����L��yu]��iAk��©2]�~���ޢ����4�pF���
��j�v�{��C"h����%�s ��2���v���G<�ז5��WҩHco#+�5|������m�W��
q~.Cp�>�(���I=<���@�%|���bS�)q�pY��&x�~��ߕ�& X7m)o�W��8��)�ͼ6O|[7=�ʸ?�~]/���zs?���e�o��Q�k},dW �܂�S�A:�����	����V<������f��!�f+����u��������%O���i?�<ᔤk��t�b��v��*�E�B��@�I.aC���r�����w�x}�`&3�1|���uq��hM|o�����n��y�?7�Sx�A~K.+�KR�$�ZL��s�.R��F���� �����(-�f��u���שQ&H��%Yѱ�wNг�b;��*|sT	E�f}���"��O�u�����✨u#�Aô0��b@�9��Ug7l�(��0�E�V�K��A4�$���t��YHzH�'��˰��.wL^��ѓ:�P,�W�|ۨ��E
�k����5�����,�`7蒘�}��T�$t��E���%OՇ�r�>�T��Y��IR3s�V�feh���f��wk��v��Q@_n��C����z�!�`��./�Y��=�;��w�Q.<���������ۧ�����{�x�9�G�=$&%�e�$A�M=6����d<�u}RR���<����P��O/&+T��ԑ�'у�b98�E�8XJ��2�� A�+G��Պ���� �>:�a2k�fͨ+*���D���@����>��~��P�c�P��W��v �(�I����A��)+�Hq�]�렝x�H6ް���TZ�\�� ��爎����ᔌ*}�g�{y���&��L�i����g��Q�AL/��>I�b봱�A��qZp�w�@mg�_u�q�D��!ȹ�UQN7�洏��N˹���d�p ��}�k�,��8�˷����_~M��O�qxP�s��<f��˽��� ��@l���w�h��Q�\4�|R�$r���Z�0p/s��YFսk\Z]��zD��^uU��E�F�� �7b���b����f���M����j�ob���$݉�4���Ց��O���k=�ǘ<���X�?����[�"�2����l�����Q
<(�����*��a�x��vD������n^~-7C"�;�z� ��Ԉ���P�bCI�' =����F+! P���eF^��`3�>ebX��a�o�U�T�=���ۀ|�-ض0�O��c���.�wM�E�ڈ�9l��V#�0]�Co����z�4�A}�J��H�I���V"=9�.QW��|�@/W�0,��:I^:6��sI��ў�b�+����9�������T~`���&�c�<�=����w��
��=B2��L��nN-%*�bKr�ƨ�!�����J=�����@�=��>��/6��r�Cw  ���P���E�̀���,L��D�b.0 ���Heʪ%�+{$�O)?�,~�(IFr�Ȓ��2�,�/���/����D����;�4E,����?��#���ߩs��.g>!�M9mc����%���ʾ�'�o^s�� �ey��bxҧ�'qB�d"
��j(1n|3�Y��:P�n!�����=�Hj�/�u��Bg�g_�S#�Ĭ�ت��.���a��t��9�V������9���rrB����
�x17
r0-e����\KE���#t�N����� #W��(}�>�J����T1=TV�g�|��PN�w���d����5詍s�{�.J6r98U0��V�j"�����ƠXbt��l%�] Rb_3_�]�I+�F�,,���:axI[�Y�g���*��+@?zI}`y<�37ۄĚ�e�;3H%O������2��Jo8��}�!2)�V�,���«&���K�W���5|���W��\I��"\���_�dur�z����bߦ��sD���fM�2���'�ˣ��p�6�H�Ժsqƀ)�s�	f� �MT�݈͇�Tr&yG+O�0��=�V�0aX����
22�
ݗ,\����)o~��v.��A���u����4��N������r�!t���U��UƸf�L�%��
��tR�w~�	{��1��N(�e/�;Jp��YE;k�?���C�9;B7&.��.�f!�k����I���Pz�ݚ�ݦ�J	��D�QK�?�hʲ^��Y�[��^��n�]�ŘM='����}nH/����-�x�s5m�])W��7�,G��1иOϋ[�,?��cZ���Ss��#��m�#m��s��*Ц@�P���o���D�d<�E���P�"e���.J�W�q��|U �x�p���V�7�x�|h��LY5���6_#�9�Z��uŜ�����V��(A��p��i������ˏ%�zR�IÝ�`��7���b��ݴ��L;�깲� If *V�' �V�	�iݠ{Y�j�k'Tޣ���9�m��n�%W���Z� 5��A�ciYTQ`�j�I2�Zȉ�j��b�p{�{0_����`o7׺#Y�.E�d��c��Ԙh�����n���xH)l����;���c���^�:��i�z�x�5�T��q�#* Aa�"�^�q}jj��9[��rw��8�#��U������֚�D�v��V*v|h�h9�c�C�W`LI����N%�#�0h偸�S��������yD3W��}��8`��+��p�A�J�f;wEd�I n��l$c�1��vk�
�o�8���-��1E	�n�y��	�\����kbڳl�����n�q�2��O`b�3^�o��c��$�I�d�3&:�k���M[��vـk����Jr��Z�jL��GɯǑ�����Q�Y�F6�:�1��w���܈��:��3��ȨP�=��ڜϡA�j-"��k &�l���3t�͙�tx'����A�Jd��>��A�@Y����k��*�� ~=�n6���mx(檑�W�1�עk}A���)�	8E\��sߢ~R��1Q���d�ҋ���5��ʻ��w{�*�$_ �oX:dl2���m��*(�㥚X*{�r�� K�V��Ne�x1��b8li�עr�@|W6��)y�$kz�d,��6O�5�8���'H��3k�:�-�3S���pspn|�H���ּ&�-�ĵ�
q}�}:a�&�Φ�nG� �'t��vU�^B,��zC��
�w؃K����3>��;i�4R��V���[��2�9�t �̴f9�x diw����� a���6�:���Xx<dv5�☹���N@w����1 |��U����W��U�o�u�S^lZ6�}�R�J}��By���`��ϲ�9�F%���,fE�f�D�`�T�]hB�e��H%�Z�v,%y�lT���T��ޗ��Q�����~���"��mD����U�FtA�X��?���bm1AC�$�3�_ݐ�����Iu��E`�� ���|��
�|Ė��?y!�h2Ίǘ&����$ORK�S��
_��MEVw�k�7Xز����X����HP]�i<�~�j��K����C�nL���d~��.�<���/I+��Hu[ �K�vL��ƅ�"Pk0�!�S���W��sT�`g��~F�����'#�p���R�e�v�F�쨻ђ��S� ��VT�:�	$���r�3�.
�m�7�b<���S��^��*�ƻ����NY����h|qW�0�S������L��#�Ȅ�+�+5'�s�wb�Aד�j�dhA���ȍ�7B��Hv����Kv�"���}2�sB���R����I��&j�_&�:�g˄(0�$&�zfN�;*�۠k^��ڡl4�C9���m�<���Zznzi��X���[��qb�]Wvi��s@�P�R^��z�f�3?W!�ja&5��#@��fX���H�����9�a�5�1�F�閆0m
��
c�������?�R�圙':��c�6��c#�az9oG��$��d�h:>\�(қm��s6��j��K�l�͓���X�e�|�⟊�ո��u���m��BJ4��꛽�P��0ؠ�k���(c�
�Nʋny�pM��� ���� 2��̠�'�Y^���rX/�I�-���>�Z��!}PGMs�����q�ۊ�����8SJ9���?W]�΃~^���
�+,d�`~Z�ƕ�Zo�j�D�W�����75�1n��@�!AH0<�I����!�}� >�P��j\�#��0���ș�V�Ӏ��w��.Aglr�
������{n��5M�o"�+��qqk�Z9�֙�9	c��9u���`�ь>-���nJ$��g�=�,�z���~�n�>��=q#N�~&T}�Y���|x�HN���Hխ�#&�	��IPӏX��(�+�Fa�0(ޫ�Mէ�E�[õI;e�P4����[�=�H��e[wyz#�R��m��P���.�)�]�F�I�5;0���RN��%~�kއ��5l��f��l����E�_�Q��	�6r�u(z��/{ꨘ
5Gi��$�2�3\`��G.=l��b� ]��f��fl%p��+�i���q������2/~�5��A��S����"x�jي�Yo����d�N��0H�a:��χ�~��8�PĴ�/���U�<�E���s)rz?H��j*� e4�/LK%���'S؁[,f�c�c���j�>��4<#4�(`���6�3�@��I����BB��UY���:�ɛ���4� <���P�.�,1����������~QZ�.XިWIy70,�p���:���1�x
��(�VW��S�s���34UD<��b�B-�u�
^������CI?߽��Y��]� ��,[Xl���l�Ҧ�PTT��PZ�z���	q����`��0)"���Q]m}|�>�n�MH���-*T�K/o�G9X�r'�D���Sc�jC�@�ҕ������g`#�qꖰ��v���T/��m@Ya4�e���݉�؈i�ŏ\ֺ�b���%�o�R�P��eS^���t_OW`߬m���I�0�!�ڒODpu���@���\�Ԯ�fE��ЭsqV�2@�^d�����uT28 {�+�J��Dk{ΕO��#{� ��5,����z�wo�ؕ��Y�M��P0�
eN_��߈<�\]u�ɞ���$\����w�Br+)aj-ł�	�
r!i��'�zs�����K��ş�\����|� <A��Ê��W)4��9i���.��H���]��q�z��^4Ep�Lo�Xo������/p��%ʪ�.l�LzP�0�R���)I�3;i���,�G�Տ�c��cn��[K����T�<�s�Y��@�h�_��b�!M�>�����e�����U�{�m�R�UxH��_�*tR8Ifm���M�iq�w2��&����b(R4L�[�.���&j����P�Ӑ�V�!����n�X�����]�h+snm�����F��A���-Ӎ랗�bv����''�;������|`�	ʛ�c)Hإ3}fD@�D����1Kշ&��}�4��sʃy��Y�,����������G�$_�Z4v�)�=��j�nX��B�k'����e�<���MJɾ۩y-�p���(���v�{>z�}�{%p��DE�����8R�Y�}~����I&;wg�� o�*���dH��_��D�~L���i�^�hdm�q1ƞy,��=�ˍQ ��g�ĩ�"������d!l.�^e��7��ďd7F��$����dlO'������u%���ً���{���IS�����Zvц�A+b�oP�"�χ<��\� �,�y
f������' �B\#��i�M�<�K�qL�Bp�J���lX�a�cC��Vn��j�o|h�@��G�e�6�8�LqU��;�z�Ê�Jg��#���@LE�"*	U�'��%X�`��'��⑺�۟��N��t%���;��=�3�(�60�)�@ej���S	��]����� o�@ K��z���|�~������R-�Se����>B�&|�B�����
)�,"��d8e��^ǀX�bR��Ai��N7gm;�L��+��C+�y����H��'�c��;|4&30C�4ԹW�<���4�Z�h&~���m��2:{�i��u�Wz�;��"�'��:a����+�{�m)�����^��E��Ǌ�7� ����ܒN�:	��G���>�Cj9 p~,�©���e�����(!;�~LR��m=?Ѯ'��1���L�`��dUƟ�!ffl�������<̾�;
&�fS�hν���\���Őʽ)�\� �.�J)��s:BaNȢ��p�:uX�D�"�ϑ~!�c3YT�e�������w����BH�1܆�~!	r�c���D��+���O(h(��b'�e�����H�o�ת6GK��c*p*��,Z�� �����j�<^�(�9~u�5���/I�;��m���Я�6w�c!��=U��*�5%lҁnh� S�|����6XX�`��o�qlp'��[���[X�j�D��§��X|<����������<����X�v�a3��^i���(W�)��҉�CK��p;���Hנ ���K�e���,��n[�Iw%�0Z��ޝ�d�"��l>°�D�d���Ar��epY�u����j���KpNOɣ��R>M�#\?n��c���@6��}�04jV] 1Ϲ�����1� #p���z�]��%7�r���ZF��xD�_�~V�>:nC}��[GՆc���jJd]!��Gn�O36�,AH��Q�;K;�V���dX��jo�ZD��ǫ�Omׅ����J4������:��fWP��Ք��0���ydf���١:�zUN�����'2I�P����E���Z�<0��zxG[�w��L�C�����n��	�$Ŕ�<�0}��l96�s1_'��g�6R��I��>H݄^P�g���;���pޣ�ok�ǅ�^��C��7yF�u��^ܒ��8S�k,�*�tr
K��~:��AH�I�)�|�/����BM>	a~f��7��2��!v�����=�֋#�5��P���v*G|V` ��g��fZ���ŝ�k�k�K#S>',� �-Y�{9n�g��2����x�ms�wWT�9�P��RF�9/l� b2�$���p�wn�K�Mm��X�2}+����.��Nٌ�年BtBḜ�l] ��Kl��đ�m2�������*ϗI"��҉��U��C+�N�A�-`��k4���a۲�!Ӈ�#՚��u�ܘ�{T��ԐE����\ͣA�/&$�������U�]�_	��P�iڛ-*3W䉎?�.]���[ן����e^�$�+%?Q?țQ�q>��H���>79����,AW�D���}�H�2Y-��xr��k�Q�d�T?ګ+�����w�u<XZc���P���M4Q��W�f��&�� ���'DZA���؟�hڀ�m����"B@j�8��
P�N�p���^x�ͣ��}�
7����
��b���~��������i���R88�����O:��4Fz_0*�:z6�ǰy�!�� cy6��z�����>JVԇd�4~������m���w[��� l�Lm��G���z _�&b/��F/O���6l��5۹ ��;��%6���.�/^rוEl�V�m@; �(��R��c��ek΃�aK�J幃ۻ�Q}���Kw]��J����<L���-�>d\��L�EwS{��������2V��^��.���w��ue@�E�Ik�0R^�;fw��tf�i�ݱ�.�	�_#E0�R/x�i�'OQ^p喢�'.<��t:f3����t����%ȯ���^�uR���Zⴍg䆽\P,��oM+�n �����L��=�be�;T�^:ѹ�����-� W���9��D�1�p;oDi��0<�P���3!�����_�<5N
��CI��"�|v��'��nNX��&&�wL8���m��OHg}����#fW͑�i�a��nΏ�y��E	u� ���cx��d�_�\*�oE%Os��6�7���2(J
��S�W��y���M����2��_3���&�oX�~{�ԥ&�^*��h:q�X6��_&9e��sJ�p�g	N��u���]��f6�׶䓵�g��Gߚ�2�R��{�n�\�1��3��ny���EV����«7ǈ
�/ӈ�ߤ�M4t��-�E��|?(=����&w�C�!Ը��2}���^�Q�NZ��в�$�֘����-��� z�w��y�3�A��H��n>
z�wi �91�Y&���E��4�H��	��(�B�/�b�ޕ���,/Lh�H<_S!�DTm��*-��Q���0��7�v�����^�����+��6�ԅsc����0������ؒ��o�q�pe��Y��0�(�ܙ�Hz:kю(�D�@�4�����\�vGw��߈:��~���f5�.�霉>��q}��D����p[�f�=XZ~�͕�c�x��zޫ]�Eς��R��Yŵ�B��g�,;�=�t*G�P�K	#����Ҋso��)�z@v�\�O�S��ve�huRA���k֤�Ap�o�;�P��FG���`�#��Q���/�A�!ҵ��(�R��*zL9��w�t8�{V��\����d���c��H�|Fj�9��W���;F�[��H��A����Y�πt�{9�#kC7�guiZ�$��S��$�\m�74qɒ]��ē������#���BI���Z�(�o�C)����raq���/)7��rU2�a2��@����B�%���7�U��wf��0V��,�������) ���Et	A�2`B�h�D<(|��}�ߘ8D3��l�k���f؎�� �%���<KF-���*���5GB	mW�-E�;w+Mm�o���n�O���x8u��yyC����u�=�]n�
u_5Pf��)T�ؠ�������o�ֽ��A��K���~;�$�/��j��ǧ�M.��]u�D�K&ۤ'=�)���ү����cE�:î�gPK��!�W�N��rN&$��t��@�?�ےoPD!=�#��4X+vCr�0�1��?A�.Sܿ�;�pIP�/��u�\��X�
^f�b{��$'�Y�Cz�N���n0M��+�b�k���������3��l�=���tC`T���>�Xɮ�T�S�Ǥ�9;\9�Okz��\~l�������ENF���f%4�p.o�wK�D}V�v�V@u���>ї���NAd@]�,��e�L��b*kL*U�Է���|�}^�,z]ƅ[*>d��"7�ʥ�x��	��bb�6_
��T��}����CE�^�â���潫7F� ?oa��5ep��aH���$��z�3W��~��0�zr%�>�6�5���5�a����,IT!��ݝ�����@T���}޶�x\�ަ�A���<ي"ʌT����ҿ���@�ɺ*#f �d��ك�^��O�<vԚ��9f^��o������b���_�s���ӀS�laiA"�T~���cs�t�y�=��WB�ur�X�6�iL��B&��<�e�a�ݑ/-�;�m2y���R��Ō�O�����V~�)-cR�?�i��>���>͉?�=O��H���#7�x�h6�X�*L�2_>>�Un�05"]G�*����^1�?��A�bn6�=�$�7Ry����mo��w�\q>��B��q���q�N,��VP2X��6i�-@��\�qX9�ʣ����tC$���+�����b4�}�1�fj'�J��Ǖf�2���jf�ь�]_����i����L�$�6P��L���f� Q�}�'l��O���&3��ˁ?��}�l�!oĔ�IR�=BReK8KTv�(�ڟ�ʙ��hy�W��7iQ�/~2O����RF�\Zl�����P���˴�?�n � O�W&����p������d� �`�)N'�U�	�Sd���=BΫ�`��웂G�%�@!O.���"%J��Zde�ӘW�"vھ��xG��&�Qo����-��U`�ڿZ%�>����;Ҙ�)h�Fi�v�R[)ɩ}�|U�j���Ѽ%R��C��i#�А����\�u�3�/��b���>n�Zj�d�#�3�ʧ@����9s��<8@��(�ot��q��bv�=]'iU�I#����q����8�3�V�I���Qƴ6��fv�]�Hl�%�\T���T������b�Ju�	y;~{/��(b^����#&��z ���9O*[O� �8��~�p\s�u�DҖ���=jf�c�o�cwI�>����a���?4oA�Ų@��ޒ����S�g*t�ɥћ�!�� �d+���S_��Y��M(�-{�A���i;���Tl<���_�����2�+�)�*��'���vn�t ��n���j�-��nŕNH\�b�/���[�Xh�!�ڕf�����2�Ϸ7n��@��v��(Ku��)�����c�����*�Az�`��&w� h�kP��1�/h������L9��4F��iނ�.7��
ڟ��2?�X�7kf��m����;rn��5��ݲ_�~�I��ƭ]�m!,o\��y�aI��Y�li��Ul-���6
8e���st�&�����}H��ğ� A�O���F;��S]��BߙI�D�"�x�:�9KjI��8��XH�m�C�A��䔗۾ۓ%�+���*�:Q���&c�:�oI�mLࢦ%u��+&������h�:�x�M�9�J�f|-���� �T%5��稣xU'(�R �W��s]Nf�J>f8�BhV������n)�U{��p���΍D7�ԣ���^\8-;�P�q��s���Յ�h���1���N�C����dJi#W#����	;4=G������>��U��xmll��us�|��`14��� ����#��6��s�;aX��Wq�`>갮��8=[��O���5kha��/|Sʝ6A���y�%�h�] ��k)L�ň�cq����Ny>ֽ��J��$����J1�L�ڙ=�j����wl2႘L��OT���[��aٷ�^!m�z�	�4���0;X���~���E'k�1v:b,�g�:�@#�\��Z5X���s��� ���&F�G���x������?��or��wA�z��4�g�!�յ�{�n��4����m��ܛ�{���r>.�z��k��� ,�ᖢPBe�E9��-�}eǜ}�̐�=m�m_��Jnȏ|�{;�cȘ�Ց���@�zL�Ėe��̏3�L��a�@���겒u�'�f�J�H>�\��t? 6��ږ�����͏��� d�F�' �"�0+�_(T������ub����uJ��
�7Ȓ?	�9S*��������T=���c!dr͠��}��5̽lj3LڅUe̉}RH�}j��MV�j���b�}���.�����M)�cQv��d�xD���2	��y�X�F��0���7Q��N���L���J^�w�*G��0Z?*�����- vfn� ���������\�-z���3\�T]8���OH�$\�̃f��u��$A�Q�9�|��\��b�զ�@�#^���)�fS�"<[y�eGI� �Y�b���E5�9����{U^������	n��X���mͳX��tYa�!�6ꗆ��p���i�d�̩s�m��(�c|f�2rB.a�4JBi���.�1,�����͸���KS�5Jϐ�.�˺�$WU��:)Bb�cqg��0@�}������*�,A�G�1��������o#vsn��m�&�����!@G����eI=?5���آ`m��&��q�~)!77,3nf���ұOM���ĵ�aM|����'9���b��׷ot��X0��&�,�~��U���8K��7�\�_��#�Ǳ���%�xeW���x�s�/C�Ԇ�'�+���-QQF���.��1��D�7�00�����}>���u��竊�V���[��g�d��3n� &E ���%��d�M�B�GN{�.Z�I_LHZa �CG
x}فt������Xt�a,(O���py��k���z��?�.{�BKW��Ê�݁�f�?r�G��e'}�p��uw�*�帅^U|3�Qk9H�.m�˱~r���6�k!�Pen��̔�i�N�X�Bs�w�^U�d������t��r�^�e9�1O@�aGno���k���f��KS~.�!�q��jL��\|���-2@�B��0+{�#���~%� �X�l�|����c�=�:SttC��ZC �Fx�_e^&�''s�YHIXK��-م�t~���ɂ%��>}��� ����+��j[$�䵚�Ma(��rzk��c\R��Z���|2"�X]3�ܮi,�e8)[4C�ơ'�8J�SQMEZ� ��(�U^ M��q��
�Sl0��NIs�@�Hp�f�u�( ��t��)5�*�7+�r�h�O�ǌE:�Iͽ�e�"�������ϸH�y8�.l�^�)��o���~SQ���u����=uv�c~�[��z�v��u�5��HA�%R@���9�N���WHY��Q����~M�ZR���`�u%׆`��q�� ��de8�ZQ�ޛ�ϗ-}1[߫�nZ�l�uC
��
�7�'���w:�0�͆�U�iBG�-է����B�t�w5*goR�mv���'y�{ʹمHe�=��2(��<��x\"�K��+T�U"W��4\��KZVc.�|�/;Q�O��w�駬�_��"��˧"lJ���{U�j��^�|�~���T��=��Sem���tbQߟӂ簻\��R6��W�V�z��%��.���{SVI)]ed2�9e��+�F��;/X(��G�@LiK^����7�Ms��<@��X�(���jD�,+Q�yt��'v�d6B�̡��,^PU��xkQ���jk�h��)�vJ/f9=w/ �[=)��J��2 �{	2�%	}�����Y?n-+�S$�+l�Ֆ�ɦlfK_��H�bGe�.�|�ѹ����cq�i��0ad���5q�������ڦi��w�5}"C���c*�	��V>t�����K�Z�����:� �CM�Ѥ�������2>i�U4���V�Y�ce��z�!��n��#0$����DG�h��S����~�?��+�����/)�wߎ���!���Ȑuv�U|�i�W���	UY;Wl�d���9_"B$��ݑ��4ь0L�Q��$BɃko7���
���A}nJ,���hqw��X�<�?�����տL��Z�n��3S�\zɧ74u���q�v�W���3���*|QDrP2r��q;��SD=�}�hSDě�{֐Yg�$�
�"�ۑ�ň�F>^�i�+,�����\��������7�~ݚs@Ǌ==�=֍��]$	'�]��Y ���M!���H�����H/���A>S�)��Y�r�������H��0��=r�æp����HT�D����}�	#V!6��\��u>�x��)�j���#y�T3�ŝ�_����%O�"�ڵ�y�ƚv�	u����45�\��i���X>��HWf�ր���Al�=DS51�
\�򈖂��eC���v�M�?�e9T����M�Ѯ*��_[�uRN5BԹJ*�e@S�5zoX�g�<��6TkHM�YV�;� YÇ�x�u� �`]*�����

`���*RР�� ��"T@�'K_=�o������������¸`��ҰM����V�S�;��a̲�7X �V��T'��`U7�Ht}�F7��(�	�8��(a��dK4�K2���#P~�y�Fi�Q��w��E�����R�&��p����ž![.�=����5������R�����F!U����(��N�kP��KnVGxAB��>k���@��A2~g��Q��)[c�p�PR��v2Y������,����lJ�   e�-F/���}��T}�1�GҲ�|]���U��u��0�l6aݿ���C�ݭ���7��#�R��[����M�q�.��D�m7�R���&_I9>k��iJ�����ܲ4#;�ƘC{�q�j�p�(C��V�_�������\�0 n�c��u�f�\h;Q�f�K�˘�	(��0S�ͬ��ؖ�v��q�=���|��!5�4t�Ϯp�8��J�1�:�FNNIǖ.&:ϯ����{�/�7�Ӿ�J�xt�f�?:����~Σ�w�X�WbY�9y�c�7PCF����{2�%���s:3X|�юxDϿ�gE�t�ya�Q�-[U�U�OYK�scM�&����n����"�rXU����/���#�ƿo�+�Ÿ��s|w��������U�5�̿�r�텯�e8E�tӴѴW޺�SM��sz2�y�`��!$� �
Y}_�.��]�E�k��v�8q��@)T]9�����2����|��y5,ҳ���L���VZ]��{���mui�A���NG���D�򇦮���K>�@Y$e�l�iD��6�w*LU�yi8p�FC���ު����J�R��g��uO�]Q�#s���c�i��&�p����7!�t�ӝ����_�(Z_��pI���MΥ�-���إB퇮�eI�`��ÿ.�P&ܳ[%��L$J�M��q��.+Fv)�)��z�'���<�e�_/Þk���i��0����;G���05`B �|\����{8s�~5�T��d�{��g�=�a��p�����KÕ��
 �#?[R{tmz�'�uL��k(�<��?ldU_sT+*]`�g��f�q����9%>�OJ�C\6Uo�".OY���R�Yj������&s��>e&��x�@a�3��͋V���V�.�����4B�#i!��9ٴ�����G(��ØC<g�jk�7���#&(S��Q��J�9Ǒ��u	o���$[Y�PDފJ�A���6dW������:��O�����TJ��UO��-%���k��%%Li�T�ݓ�{�:3��w;�9o�B��݊��A 0)S��ş��϶�q�yi�H��\Z��. %G�g��c'�f� �w�؉!��Po�t/�7$�e[�d�|%�����!rv�$��=���h�"�� �M�)�-!&X��>3~͈���g��ʘ���x�K!�~�gV�[%ْ��D&�QA����M��N���q��v�0^�;�:���*�l�
��������o�2i�vI�p��޴�DEG���y:01�U]2*:p\��I4��@c��/�����A�1F��.H�3�39=9T��T����xzn���aZy������fA6��|6�����m���9B��+ە�3��8݈�F�I�\�e���8!a�O��Cf���P�C�+r������O�[/�����K�ע��Y&�>r%�Ԅ��Q�N�Z�k�0ō��\�o��YϷ�|�I,[���U�����(�<v�f\ֺO���d7���V܀s]N���9"|���>0��@���J۰��TX�Rg�1&l���fk�o����ו����r"�������GK�N��kd�B�8�305rg��-6a���jI����f��%L��wS�iÞ�_F)%y�J/]<��lx���3���y��5�ۚ��z�!a)��x�q�/��",��x%�NN|��D���9,��A̐̕�6����KTRD�ԬB�����R)Om@}:�0@��(��0k�6)��6xY�.�����	C��;BŌ�C]��x���k"2��Fl����j���w��k��G�i���_��]m�U.U2���Z����_	gEa{_��u�����S*�@�9�������	K��敞��zh�8�[a�e:������"o�,6����d��o�5��Ld�Q4�G�� �J�h�Ԇ�Kq�0�3���o���&�Ñ�
3���y����+�G�p�m���|�LkB���s�O��U��0����*��D����J�{�"�u�Y�
����gv�/���\YR�G�f�)��(��c��/��t0���ìC�KˈF\�)UQ�&�\�����rPQ�3�z�8XZ�\�h�Mt:�폝��p�*�n)��F�\5iÀ�����YB�0����j��njW�����݊�9?n���פKA$I��zQ��ؐ4$�stJW�贩��2[��~m���~M�=�lb�@��U��_H�-��,%͛]�e&^��C��P����;\��R�2�e#�<%���5�.��2t��q9�""E+�@���ؿ�w�n~��E��2�����8��X0L�������z/u�#��a$z���
�����\�օԆ�q�?��{)�U׿t�>~i����t�`CJ�*��zc�3K�6�мz��ÁM�@�Y�TF5d�Dn���N0Q���������/Ǚ�RWO�A<8�	<S���K��`6r��b.�?���󪼹�I_�Կ��}XpHQ�Bi9쏗*e>U4i��>ڶ��C��q�D��1����?�,�c����Ipc�a�������Ɠ�j%ZP%�+vU����ZB?N���d�I�=
U	�)A�Ř�é�\�%��;����#h�XR:O�nfd���ꉑ'ᜄ�h��(�1<���)M\וE������:\YN��p!f]-��t��4�Ѽ�I~�!�/�3�*Q:���R/�^���]2h�X�}�@}_"�����<33�Ж/Rx�Er	0O̷�9�� %�c��<sޞ֎n�d�F���wwϳ��Z{�tC.�J���P<�� ���B��m�-�0�U]��R�o'��<�r6����ʱ��t�P�����j�
? �7 -��{��C��eٯth��t����Ep�}r�V����nU-¨���:�*��u�z�}��^u7��s�UB�-�-lQ��̆��3�M�[d�����}�ba�`Y��d�>���mQD僯��йP˵2��=>�L�2������5����$q/�޲i&� �$D.x?�:H�M��x�q"��y�@��H^
ղ�r�y��!�6>@sz�k�oTz��ݭ.��(hE�+7ѫ`?C�OH��o��K�|4Gۚ@�'�m�jm���m/��%�CwD?Læ��0(���v��b�8S��4�Y�Y)>��@���ˀQ�>w�KN×�1�I7������]�M;�Q��BR2au�̿�<U�?F)w)u�/H�gO�)5	�t��af�T)�뱔�nk?�"7z1#���S]_�f��z=�����䷐��6ܛ��2W(� ��������sZ0�iS)*��4���`B0e���O0�S�Oy�֦�6���T��G�1x�E����'�/:�MG�����J�]����y5�)'�yՔ��F�?��".�	����h} �q�=\�Λ�@��G;�~vt}�c��L�<v���� 4�E��5��>��|pƂM��q��v}A�Q��1���,(6HY�h�Ø�1�|k��`�Qf�G��3ey&�u� ¾��j�����[��A�c�k�ό�ybuTy/r�T����$�l!��*��k�8� ��b#}����;z}�~�/���PLϒ0-��+|����wYtɨ�w��s;��{�ੴ�>O�>�͗)O.��i��%�D&nJZ�H�z5:=|$�eX!e��o����[�Qu��W8�4��x�XY$�z1����}t�Ӧe� scP��-,7kq*�Ϲ�����|�����m\mdy+aP���D���B`����8Ąn�R&�ѻ ÿ)J��3[�[,Nb�{�P�����i�o������R��ǁ?��3鷠�bg֖�c��k��y�+�=�|������S�Ƿb��������v�*RD���}�_\��C~�9�^���jll��>��2�w"����Hk�2�@��-��0���sK@��?	���0:�L����@��5�Tp̃:7��}���ŧ/�Lx9&������/�Ót� ��*���>��"�p�Y��+mʛ~����5��O�+��R�[�xj32{�Z7�L�Gr&�)t��tioG�?�Ǎ�?-��?��[�˓���'?hQ=�N�O��8��-r#&�ݳ���Z��DR�ᓆY��t@g��@�o̊9���xW��<�?�1��m��{c�����ᛀ.)܇p�ˋ/�w\�m(_9��HV���H��b��Py��Wn1����xT��+>�}NL����>\|�G<���?������|�嗩��OE�㶯�A�0��梑�/���38QP��Q�'�1�K�.6��I�6Ns'n���hqjƛ	%��G;�O%1B���e'C���Ho�P`j��j~����ӽ��Q��
2iL��t��
(^��K�gV9�R:��Ǯ93e���m�E�e���z]B��c�c/�T�|�5�����s��@-g@bz�E󯼢���(@A"����S��*�k��ٺ�l�ҼJ�##Zm�~����h��~Vbk=>&�O��3`�:F��<Je�۲����G`������`NZ3{�����uSK;	x��L�
�S������v%_�&�����`s�BmuO�1J�[�k��z}�o׾+!�0�E6(�R���t-q�?���qH9�5r��1�z�w�5��X�uw�������-h@0 ǳ��*z#Qؙ/����s���� �weBf�J�n<�`��z^ȸ���y�J�{u��ہ��>�gp�b@M���x�	oH�(��MF���D��`���T���p��ᩉw��������̰��A	�Z������?=�/����V�@	H�pI��Νzk� Ū�B��(������H!Źi����8�aB�0@�e_�bS�>l���o��j���b˯\O�I�U�;�0Q_����qq&���4��>Kz�V�v�&�#hlP�����ޮ�
��a&
�y���%U�h�X�Z��7��&��A^]���m��Lމ�I��iX�0\I<�r��$B�z!_yvȐn����_���X���95�m~��6::sc�V�>�����%-?��Nn�0kRl�a,�zU�BH��_�1��_�����e���]� ��;��<��Z�U��=?$�I�1�t� �����1W|3��Al����9�@ؖ=�[6�[�o�ު�U�g�v���!���_�)�;��<q_'���g�<k�����Y0;����Qא�9�-ɮ�=���.�<l�y� 'Q�����&��@�ރzEa5*�;�޶��JO�'���7Q�_D��`o�d���-�� ��I�q���)E�[V=ޠ���/C�09�5:h��:����hlZxF�hn�N�cс��	��gP�����+�	����#�H���X�f�vr,<A�" ��ou�ak���
[IIe,y��/�7J��8B.�����b�*�Oe� ��Z��a�� ��� [s�U���*I�[��B�Fw�O �/�d >���y��-���K�.E0 oP1��,-��/oï�bv���N�`�f�`�Xq����s#�)9��^��&��[P�Ζ�4���L�����������xo��i�_��,�4�8��3��kJ4qt��>���$��������	*0�aݥ��e�WB�ҥO�	,�I �Kж��)`�s��{8u 7��6''���'�6E݇Lg*���D��� �]��Z94�ql�:.42$"���W�}G��$x����_�
z��f��af��#Κ�D�"�l�m���*�7�;u4x�kY3ZuPQ',VT�j����9's�jq�n�P]��w���kʙ������]8y�S�eDjp]�Ac�-�����V��ayg�V���/{�����l���Ur��[x]��5��!,��rsMrW/�O'�3��C�!�q~X��r����!�۹���ʐE�=E�����n����
��"��\}P�g~�t]��؄f���ۥK��%&bʓg�z)��,}n�>&.	����DG Q�=yٽ�Ō�D��1��!��#�*�������2����c����CrO�����6ݛ��aڭ�b�Ӕ���b1\pr��f-0RԻ��"�)�*�v�id< �I�R4P� ��S������B_A��X؃}�%�yO����.�ǀ�L�<e�/r\�Ǜ���M�U�@AF�Y�
�Q+^
�8�m�pL&RF����M��Kjb��6N��z������0��5B9[s���"3�I��-����ph�/���O�Ԯ�c��xp4������ꃙ��E���aJ;���y�������{��"�����p���wX#'�ǳ���(u�ҝ�F���Rq�V�.�0Q5�����	sg�:!�M�� 3��A��\�3�*~�KaZR �RUm9� h}m-�!�{���DoOk�c[(�����yp���#�-�Rq��@G㱪6 W�`P+�TVO��|�'f������?���#A�:;�i���?3��?aE!ζ�U�I�a�vRLþ���G������E�@Pe���9h��U��t�����m��L���i��Ʈ�{��,��D)�8�$,��&��faa՚q�;Y��Y%�d�zR9�Hۮ�D!�+��:�8ȥ\A��ҏe�3
1k�O!|��a�>�?�*ij]����Y�~R��aU������}��Y��X?u%������aX�5&x���ь����Y� 2^Ƀ�h� c����<m��`�nL��&���9Oi���bk\T��8Nh�-uJG��ӗ�|�m��:�d?
a]K-���>�&�K�c�-�{ӻ�����
A��K ��+�\H��/:%��g���9K���J�E7���s��V�k���n����&���
��;��5Ur�09 j	�r��j6V�q{��#������Ś���� ���
�^��Y'��C��8���ȃ�Y���������3xZ@���;]S*J�#*T�����u��'R�3^}��y,����t�ݟi����-�9X=�( �຃3��-�� ��t���*�=�����Z�FZU�9y�`1�w���~��Uf5�:y�F��M����M�^p��������/JCĠ3|�\�|WU[$n5�g�I���W���F�j��$SA]0�%�a�2*)�1FYSԤ�cF��[��D8.m��"�E���j����j��-���|��?*{�M��@�o�d9>�w	hWw��{�ѿ�?�V�m&�� ��W��:iP���т����(��Q˳��H�ϑ�N�B�1{tvWdU�{��hnX,t��Q� XA�k�/O�8Z�5o����p�n�J���TF�Ƙ��[ߘ��L1'�D��,D-�۵y�p�Rjx�qF����f��z�If)4Å�n3"}�co�aE}��4�9:W��F�DK�	ky^�KU�R�Ǹ9o�&%v��f�Xc�Ю,/�Ai%eX$����~ztq���cw6�o*8�I��!�����7�k���j��$27�fM�����e�7��S^jX�YT1ȁr����Mf�+:x��n�C�����&&}pMjA�u/|,,sD��;.oykL�Y(K�`�zW�{@�S��^ܠO8÷)�:F�O�T^1��+�켢}��W���.�zK4Hl�V��G��{h7���^ܿѝ��@�+�\��,؏���K�p�v,�o���8�ٖ��I�A!4MT��`�	>����{�[s`!.�!�����#wvD�G�Kw�CW�6i��d��T��XjL&iXM��_�z�Y*��t?���Ϸb���-�y7/�M�n�|a4J��OPzj��i���/�}]�߉�F���m��Ԗ~��lY�i)��*��o�$�dJ��3���:�0g�㴪�β��_����ڏ<�hjo��Z�h�N�А�F��j� W�'����{�߇Ӱ��⸳J��~m�U��8���ϼ<:ѮRޥߒn�ݘ��u��q���9�́��$3��Ҧ�;\̠���$�k8�� ��Y@)��#<�Gx��/�tr{�#_LS� !��o{P��|�!�m��K�=t{}���\n�E��;��c�"vA=F\�rV�W\.����ݪ��=ڤ�4��Kh.���0�CP^�2���P*��ܙ�krj��'G
�'���\w@0��F�3�L�՜�v�'�*K��r�Ntm�"c�<s��Ah�TdcHŕ_V6�T�K���8#�kzȐ�ZP��+5G���q",����@/��0�[��Rr�|]I��TC]:�^b]��-�9�J`�6ʯ��3q�����ikH�e��j P���P��պ�*J�=@�Fl�"���t"T�[��$l�B����Bǰ3����I{U�¥R燚�����O!P�ڤ�ȗX
��tq+�� ��뻧~�藥��1^����^-�L*����w��c��>�з�^#օ��U���1o����õCޗY�ذ?��滆l�K���h�9����B�
tuZ Y����Zј(��(�J�7��uc50��{��^��=�"p�G��'����o�w ��{o����2�����>�"�( �3��!5a,S(/�@w��F�D΢��W�_�I���N��<���G�v:�ȴN*
�m;�P��������6���k�Z�(X�����y]h�`_�p��صA�b��I�>�:B�{�3frse�>��n?�9B�ƅ��br~N(=���� 	W�"tҵ�L����7]ƙےͪZZD`J�"��s�}�n�`%�
�RZ�̯���:豴F��W{�BD�/�:���Q'vüT�oH���K�����x�O�|Mohc6�����jsU:2_Zن�|���uQ4K�.B��#s(���a��u$��`&���6f��&O��}[y\e��x�h�S*�'���3�y���.�s�$�ϢP����l�#ӯ ^�$�)�8�p�h�4΂fH_�"���/c*t���W" p����߁b���J�(IƊu���*OE�x��NqX�N"2v��^���Z��t�.?n����"dsd[ãW�C�#�OȪ����U�-v�U�=�۠��A̱ۅ5H� 4a���E��<C[�Qȏ�-��-�t���.�p��#y�-nw�;O�wt�vn7��ԩ;�BP	MB�c�l��Z�}ñ�52�2PN��74=7�1Ds��>��oeJ�/���fB��~�����^�{#��?����}������c[z@��ʄ{х���,��u�n��dT�l2���)��n~�:���I?�}G,4��}([���7]$mJ�Ux��2/�\h#�TA{T�{���g �nI@��ch� N,MO������]>i��0�8�����*u	^}�~�+^j�m��(��%�����ԓ��J[��O�9K�-L�^�7ߟ�a��'��49;����=��\3G����yd���]��C��k��$�SHa��_z��ۑ.n�JS�z�-lD%u��������K� ��f��r���W̛�>?��#��i�>����&I�__`Y�}%tk�/T�OU4�8�H�1���fQ�d�k"F*�31C�~�,4T�=���S�,�r���L��� ���B�a�x/���6Z�	�%�3���|)' ���z�����?|N�؇�r�3>�,�1t�/�B��r�BEA+>_t-�����O��i�H�NYc�/�{�k���y7"A��CͱܑQY��(���)J-;ET�����&iN"G�`E}�x�[���sx.��I>S3�"$��YP�,��239�J�G^;�#�m���l���L�ag�ƪ�J�J4��9����a��ecYWќa��wߦq�	>g�C�&�q���?���U�l��F���N�a��}�<we��ER�������d��΋!������#��{}�o$19�<?��8���"���\�n	Qy:y���|@q�c�� 1{�����"�N��+2�!n����C�8��\-,^!l9���~��V�w��(�#�3ң���"�Ӌ�z-���wXwPsm��15����dJX���(}Y}��kW}�͆�����s�ݽ2�2��"�x#��b��� ��������<ޟ���������ۇ���4hw�MC�Ga������f��?�w��`&�x;��O���lMY"��l���u�E7�u�`-;�,/��{�n���zI5Vx�`��w
�e�q~6�g^��X}�qԭ�G�����ț����G�-�Ɉb�@~+ro,���[��E�X�_��QxoyL�tlp�f]�@�L!�>��C�
_�3�1��}���s�e/�#^�Ҿ��!/�mR]�b��w�cj�W@2�#(&�qF<�0X��l���
��G�u�m�x�z:�`(��7E���u�Oj�C* FG'tdrG0�>:�y��U���H���3���&E�B@��*Q3z�a���)ޯ�.Cp�25�[=�7�l��?�@"�g$�˟wM��P�gU�)CD���~�>�X��*:�=C��t]	�op�D9N,j��B��ΜX	*(�F{�?5�0�Jh���L��meѠ~�U�O�/1������?���xOje� ����նU�[=�q�5��"��mr�`�h��m���a^���5�T��\�R�>d'�,�~��Vm��$��Oe�l4��D�� Y� �^v��2��@fn�G��g�f��N�#Y�&�Ź׊/��Es�WqSSXN��Q8}��������$���2�ς#Na����>�7�7���0 g��"]ݳ��G�W�x��7�Gpe��]��ټP�M�C����F���/w��3�@���S�'�Q�����/��!�����Hϖ�k�$�uZN�轳M��� :�ùI�g�p��z�A�d���ID?�~ԕ@{�E		�`�������B%�&[��g�N ��e]��C��I��o�L�x���|�x|��$� ���J����x�1�@�ixs6�8[����y�m�^�AQ�k'�������}rHR�t�����97?�Wb��H�Fn�V]'�0eF.���Ȭρ�a�ɜk�Ku��S�gF����Fɼb���dE��0ڤݪu���%y���g"���D��qk*Gt�Ε��=�e���굑�#���t��ʈ �������F�U�C��r��,�t{���<v�ZA	�+Y=$T�R*�Ga��s�Y���Kc�.Ԙռ��.[��*�m�����μ��
����%��W>��>>�����!�t\�g����39zt b�W�UK�l�(䭟�L'*>� ��18�hǋ����C��0�M�䡲Aa*�>��3�K�d�+������7���?E�ӵ!������G�z�L�y�9�Q�\CԣK2vC�z����}L�-Z���"�����>!��QL�]��(��-O�,n��}�Y��)���� Sk�4�����#��zp���.SFT3ܖk�>n^K����a������M���=�5�F�ʹ�>���|����ԩ�^a?�q��s���+��a=�)�x��T��{#���rvt��{��@=��BG��a�Aʆ�Ƙ7p�M��[�����ZKg�T�HC��d������!�
*Yi8�:cG�cux��y!ޝ�g)*��(�Y��^�CR}(���E�7}�o��:K�P�Я��_bJ�iО|��C�[Z%q/���
[8�pT�@/e؆%���YΐZˮ��M/$?��0PʙW;�-�Ƞ{��L��29�F�_y�yP��#Q��=b��_�G�Z���_�a�K�os�7SQw#����U���a1���T#(�����@�ܥ<����8�/�ւF<G���Ʌ#�9�����D�����\-����ű ��(K��CB��#�,�O7��yD�ě=���l���CE��8\j�l�;|h<�b�f���1�s���Ǡ�6����%y+������`���)��5u�Dߪז��S��4��oK�,#�`�ub�T��
���iƕ�8	�j�?�f�~��`�6�=Ѝ�����c��U�a���\�&�x�"`���y�[w����@�Z��Z�<=1-�&��Uq��=����CЊ�M�o%��t��K�[����s���f��Ԋ?Jo�%8C�TQ�)���J�/5V����uZn6V��l��0�h��K�XN9/Њ�mOUCȬWf�p�fe���Ǩ����O���cH��<Ӈj�RNqP&C�H�?����v��G�I	\M����\�O��~�W��w,˂�8V{�7�7oc
���m/zD���|r2L,��O�6����^�ͷ�FʹU��27�%ب*�* �!���;���\R�ܴ-}�� ��x3���ޕ�'M�xP񂃼�����h�1��YuN}e/bM�&�o_�s�`*!����$����3���;�΂�
�w|	3�J�q}�b1��
��1]GL7R"!�����ՐJX��b��	��p�M˥��4�(�uw����LO怍�t�>�Ft�̿$<(H�/���N㻅��&��9mO^b�z+PL���"�x���G�W�~��l��Fߴ�����<��~�>��c��'���c�šU��O�sP>���hO]�GC�ḔFU�D}?�u(L�_�'�"O��2s�`�V=�7������f����C]�i�t䷾Sܶ��Ƨ�g�����?���n����O�Z� ҥ�1<h� ��杤��	���(� �>� �����%�MU�����q�@{�d������ھ5��i)�)�xϧ�EC��y�)�2�:�R�����)�f�[��=�.�Y�
�WDk�9��#��#hzZ�U>�]r���T�s������|u<% w/D���m,`(.��7q� �੓�+��<ӡ٧�����0�Y�
�,m��K�<&�sE�� H��b���. h�k���0���'�jQ_*i7m�`�o���7	
A��=]�����GX_�k���=#{35�%AS�����B��HN!n��4�G0
�A�\�Kز�rb�hc�͘>�c�UWrgJZ�Z>���m;#E����P�"�:��1���*��.�f?��k�yjPS �(+|:�s��$�$��?�B�.�C�����뱠�h.=�5��JWZ��D�
�ͺ΂���s�h���D�F��e+����D��j�<PN�bZ>�-F���q�Nuz��{�0�!9ii���ΨM:��.���Uy0=�K]N�6j�r��	�@!�-�G�L�J}���,UE�[̻�_E��<0��0�۶���h���V��\��ͼ/P�/X�ǒadL��u���������Y���3S��Ȩr��{^�&{�ӯo����NI�n�!�ǲZ�~E 	�d��d�qǣ2RT�ӫ��!��<�p\5��Z~º���&@�d�S�:f&�w|�����z�[�4�J��)=� K��)��6͠���E@��Ǻ�E�rU�a�@vvsM�_V-��kA(!+�E�L�՞ K[�{���\�B��	�:� ٓ�7X[#��ȧ
0����-Z&�=�
�h�N�?\�q����duV��-�]�k�j*wW^C�N�*?�	��ES�t�Pv����(r`.(6�v�dh�3 ����o��'5ש)�2�F�}k�(vN��x�*�]Y������;��B'��CF�<`�ee3�6qF�7�J(���Ͷ��xs��][>"�A�Mi�NZ������x�W�Of��k8d��W�p4��訚��]t�m��,X+�_�2���&G��W$�l�xdf�BU����Q�Oܬ�*��`?�%���}Ӭ'7�ŏ=P'�IT�A�tP�#�J1"������k_ͽ���S����CD�����
�j\~M�F���/�m�!�M��=%��&��yM�^�#�o���;ݱ�;�ė�0w��E�$�,e���d����J�d��c������:��i���]�N�8?�{�j�^2{���V�I���`���u@A���.�@R��\h���K�!&_�k݆�	b-��瑿
W[�`��-�:��AQ(#�*�E�@&�}W�rD��D9+�Y;* �	`����Y�y-ƅ�oh�JK��ɞ�tm'�{�4
���(���灱�q�c��{_�Q�sn���wz�`KH�aR;�f9&�*��R�)Q�aaX�>] 9��>����6h ��x_i�E��.�*b�߇�kcͷE�fʔ=�28�G�Aa؉���ğ�5�xa6�9����cF��G�u�Y�R6^�5��W�;�ݍ�BD��4�����_E������MV���������cq�����C�%q�o��(��%��N��qF^��H;Ԧ��<�M��f*�Q�rf�� ���AJ�G�x�S%U#���d,@��D�#�4�z�p�\�p���:=��Mɰ6l���r�;��#=����`#H�j|�&�#u������{�ES�φ�7WDwG�� ��v5r�^ߎ������2%J�S�D�#P<_�	���u��iҩlO�Y��|��.U���'\V/&C�G��Lw�Ƒ"p��4���c 
`z|�' �9�ԣs������]�ƆhĴ�C�T�Ҧ� H���<� >��OgL���b�#X�X�l?����jj��sͮ����ڑ]o�;�dk+t�g���#H�ZRV&p�C$�#�A�S���:C�'�EC�z�VjЮ�ϲ�St���D�`?��`�CrR�z8�=s��������nf9K��&�+m�E���ؚ]VР�l���#���>�ԇ�;��-J�)��Ɗ�V��[��?dj̣���@>;�،�h1�(]=-�o����ΩG�d��`ɇ�@ɸ���C�:]�>��*Z�����te�F"'4���;�n`*NS�!�߃�E�s��p {����q��x����;���߾�)6�T�Z,���tG"4ߗ�\�N�бpC���xN��,�v�0F�:��ܸ.�kA�)r�0��ҼCZ�'�[��B���g����qo�ת��B�Z�N3뉞�og���ڭ>F�T���s����dp[��Ǣ��ȃ[<�;圊��Oj�I��=^t�]�������qFc�" ?��j�$��pL
��cgӥf��C�C+|"�F�$S�_&����w��R�NN���ܔ�O�MW(�^,�dO�uc/� )����G͵�ui�mx�>;��j�H4�Ƿ�d��H�M���wLY3]��u=N��x
CYя�r��3[��&S���[�����=�]e�'�$�~nm��~4��h�b�*���b�Y�mk���<	~��S�����9�-�s˗�[���������8i֩�ß{v"�&���ڶ�$]SWt��%u����	�%g�x��%21�pdʔꗋ.ӯ�w<o�a����`Ƥ�{Vܔ�d��Ke��$��)�4��ܤ�('[Ï�4�ژv����{U�ŠN"".b��0�3R�*�C1�p̬��%]l��`:�R}�GP��ŹUhzpL��G,4�Y��]In_kG�!��O��ί� HT��0�H���PU�欛vvYঝ�p#[��� WB�V���P�F��w1��(����8:���"�y�BluҗZs�v!�@@@a�s�Z�E�x�~�uL4Ә�F�(������? ��@�9[����Z�f@����@�-~�M���e
�����Es�LX�ڹ0;>^�򪬤�j�fD�,x	Z��K��?����o�L#��'�p��X����f�g5���ȗ�٭f��� 7�)fO���l�U�x����)��f�`z�W����XYޜ�t��z�\��T>�6Qd�W�˟��T�v��_pI\��G�&���O��Ui�&E"��t�6�.>�����i��zU��	�~�
��X%k�V��!&a��m�q)�a�0�@¢�� �ѓ�'��H��(�k�������vd���Z����H�`~d���F9���m���S1�>��oVd��iq�c@�@_��j"s��r��ǔC��%r��h39��{��pj·U8?��ެ|+�@{��l~X�V:P}���i:��l���Kə�Z�u'�	i��~����!M��?��\�A���2�ߠ���&�}�������r�Kv=��u�H�<�3�>�У	�ݪ��YՊ��� ����-�e$`���T�ga�Ӹ�7���Kg�`���zh���Ͼ<�(���#�0�jڏ��nnmw� \��3��a�y<K��O�ѓwA�.c=�]w,�ޡz���ep�=�������uV}�H[��f�b.�[ *~l��<v|���R�*�jB+�����T��N�S<3paܘ3��6Z�TX��&�O
���3:�
��R�{l���%l�� ć���%k�E�ٱ{Z:�����<`3�
�/��y�}���{8��~��߲���E[n�>~"�Ǜ��S�O�&n��1��M[��������*�<��rCs,��T�1�Mh�E�*[4�0���e�n�o��hg�]jR�z�����O���*o"*���� �-v�,"�� �
�lq�#E�,�Az���BU�*��-30Dȯ;�U�^̙�!JzǍ�X�Ч��7�����8�G�:�z�C�ڎ]��q��x���c���/&o
��TQ��]�H���"��b2�se(1��`���Y�=~���p�D$�0�3�P׈�8�[�y�;p��l�fpQ�ѾI��Z<d�~?��9�ͯ�U�C?P��i�U���p	��w�j)�\�؊�/��m}c���:Q�Ѩ���MD�q���i��
��1a
�H��M��k�:����_��]�X�EA���w�W�R�*�/�	_�A���3�P�w� ?���RS�[���Oo�qB��~|����Xiy*��G�Z-�P9N���	�
E�Is'_�j�Zb���A�6X)j��# ��Y'@�bJ���\z��f��v�5x��L[�Z'�5�W�I���U��V\��J�+TU�v����X���0G�k.)�M(oλ����]X�Tx�I�)S ��p+#�.:ݐ�9�j7�
�M��@�JI�q�w����*�q�b2�"4��z�}��A�e�w^���˅C��l�v؈
�6�[&n�e�����H2~E#x�Q�9�<��
�Ե�-*�@�����q�ӝ���@�:�I��Ҷgx�.�ѭK,g ��Z=���m�]�u�\K�=ېb�]@+"������I��5WM�{�r��;�F���p39a���>J����e�s6���.m6?o�䫣^���Yd]�����L�l�;CXV �V<2�rQ)�}������ĢbI��\-��1�)ٵ�	,EY'L��ZTu�q���FP������-�����ۦ��Q�U�ɉv ����_p�P��Y2A�ğQ?e��峉jCb��8W��,��xDzv��T�YEĥ/��D8�o�;���	�2�H��`ܸ{�W��4`̇Յ��q,���g�#�,��o��Y�?�};����;ڔỴ���.5�I&q9�T/�B���y?4U���{�2I��8�N'�r!�������8$z U�=O��%4�#��\5dYQTW�t)
��Ӽr���.��Fr_r}Fw��@���l�[E˵"xH�E@�39�[b#��b�q�c/]�D��[n<Y�t�@����$sl9%�D���:u;Qr�Q�YP���}�ًДz�
��l���?��6��=~��oŭ�v�@	���D'�A.s�Zj��H{O������@4���G80�Yw����u,Nt����U�DZG�Nsg�
 �-�{W��<���,(!� X$����X�ܙ���c���'�~2%Bo��y�߾�E��!ST�߲-s���%�>\��æDo4�I���6j���$�\�I̕l�$M��v�5��BvF��Tb+yT�T���}���g	�gnJ\������3�]����#��4�!_g��T�M��
���Ŝ��`�ԪU_D^x��Q,j��N������.�_��9��z �-�t3�~�^�&�	e>l�ߪE��l'OV���^׶�}�'�=ϰ��)H����LEvOWh��o�w�,����������e��/�#��1{n��'�L3�֣]�dR6m�yQ	�� �N{Ν��� ���;׆}\�r�L�7<=�788���Z&ۖ��lj�j3�f�c���s�P�&M,	 �p�V�>Vhe�i�Az����CH6�*w��o���V�@Z�K��ЧX�o~ѱ��pF����w���"��[<݀/��<��m6?M���E���9�����^�m�'��%�����p��]m�*Q��֗�P�'�>3-��դ}�'e�aZ_�ĥ��
� ɞ!�w����B�r���ۅ���?��K
��Z�w�-�AS��凥M吶�0�.V����W�|r�+ �K�3�e.���3�!𥨩Fm6-��lu6���|q�����:�#�m)���bWR�l�\<^�����F����c��du��G��쇚Y`�a�?ǥ]/�s�0�Vb-�~7�ؑM=��{{��]7S�|@�9�bl��j�nl��F't�Z��%{��͝HF��H�9�a��Y�����j�ƅ7
���Ra�O����rV�NM�j߂qՉ��:8cP�׃L;0�KД���twf[� t�)����l�q���?�"V*��ga��Q�)h�4j�P��Y,�e�9�Z�uz'#�H�֯.������|�\7��l�
���`s΀���Z�o�w� �\&��/-���2M�l�KUȭ�Tu^����՟��Az�	�ی]t����L0wD�J�ʳS��%��h��~I��}��R�(�R^4{w[��݂�
�D�y����/ҡ�C�Eq�x;�Lf�ղ������MӸ#a,	*��A;]�i$�![�xQ���dq���*(�Z�Q^)?},�n]x�&rg���v��}�����������2+߁��Q#�gL�ю�m���m2h[��2x�-��o�r璢�Ԍ�Q�3�p�A�+�hȭ(Y���n���:����O���(���Tӄc5#�R��}�V�4��Z
��CU�z"Xɬ|�KG���B7����U#&��3��:nĩ���ꗚ�=O�\���Eݼ��F�����l!
���[7-��n��_�l�/�/����"G���=xϠ(�
�ta�����`�G	K�>�=5,��L����i�e�}O�vܹ���h�-o��XW����t=����e$5 xz�|�s�8N �����)Y�ưZA{�q���Z~G�$''|�?}�Km��2�Z9c�R�ն��'29-
����0c�����/r8Y���7�E6(�,F�]�M�f�rJ��R&t�Z��U�t����2����}��	����s�`�/��q�PX��$v�%#gr�2N��L_8w�N�e*`Z�����H儁T`ΰG�'�cW�sf�������&�P.��LK��c��N{��ꝧPz"�7�b����v�@�[���t|N^��	ꁝ�ecb(樝���I��ڛ����g�!���z�d6���}���+B@(N����hp"`k�#�K/F�בb�`�4c�5?�0�%�$B��zA����D�@K�[�xbD��2h%�x���	���r��������W.����5� P�V�{�׭����	5�*Rj�Ę0�I�Pʸ�9���K�,��"��rikx�e�
ר�W��NS|1^9j*L��Xw�rZJ���ʄ�M�S����R
�Yď#3���\1���iH2oc��oò�0��2R�����r�z�{+���$z0Rb)QwA�R��tw��:Ca�����nk1��/z}�ʬU-����"vi21&�'ɻG!�fk�N���0�-܋���ICP��;ɖ�/ɓ���iUn���Y��ﻢ����B�("�^�R2n	,�Q9(���(T�^}l*O+�7o�9�͡�/x�q|�?�㝟0�>��ݵ�R:�e l���7�O �^��=�(�}���]�WҹSk$W����_&�f:��W��e5e�m�ﻏl%H��j�8A7@}y���1Q���:�ِe�R���8�ިQΐ�{͜��Jdv)*����c�+.�$D�,�#,���]�@�lJP��f�"'�7k���+����9ۊ��J�j(~�ݡ�Y7@�φY�ۊD���䶽�DML�鞓���j�� w�Va�Jkm$E�v���N�%�.�&��'}�+����⋕Ћ�p*�%7��w��4�?U�O7�W�O�Qi�syt&y!A2��Kdo�T� ��!��-+%=b�'��/�n�sd ��}����4o�2�['�KRd`�7c�KO*��8�ai��0v���� �� ����ΣR����3��A0�ss�h����a���?��\{EI ��������s����[��$.�,���c�yT��w�r����)O���}�zܡ���G��	ۭ=e�O5���7 �u�L��<b�Q� �,[ߡ��]k�T,̒��-�zg=��g�+��9����GQ����x/0����D��-��;7a8��E��>�`��}�t�����[U\z��cO �ug����ug2{��M[}��Tc�p�����Q
��юx{����S�N�+�L���g�4-�-�7���ӎۆg����A������g'qfg�Z�@���c׭�w���l�Y����00��ZV� �BҴ6�G��s��}����}`�4:
��A�Q��y�#��d��W<����q&����v�j���w�7���>�f��G; R[;���-)����+*~F�������)��]��q5���l���H8w$��r���3�$�D��?Ο�q����3K�����w�t�A�f|+h 2H,���1�ۧXʣ�nK1>~����>�gQc8#/����7�Hv�Nh8X�0�4���t�u<"koS^� �u��q#!��\\�3�/�g�����?�3E����!�����꧎�����x���Y�>Ǭi=���dMC=�r�\m��v�hjK/ԴM}�Y���]-� �8nX�I2�䙟D�l>��v?m���)��H���N��yF2�S�W~va�}�0KF�%\�}��O��頴��ɲ`˲�>J��Ɂ�~j��*�M
-x�CIՌ�������A֟�A�z��uT�mh� ЖΖ@6zQԀ�̥EJ�����Ҝ=P��Bv�t�PP}�_����i�k"f�~��ɵ+�0���?�7e��}�e才�UD���.X��o���J���ӎ�Sf�B2��Z.
T}VY��&���QY0ӫ��!�T#�C
��\n��̘~ӱDD�x�~��NQj����l�4Ԍ��V�1���L��p�G��Wޠ{�1�&?�T�^<G>�/e'���:Ʌ�c��BJ7]pKHq�Au���*F�rb�
�	'M��fÎs����[�)a�����BxV3Hl�O-\M(�W��樫}��\%)ya�'���R��[>���Ƚ��l��Rڵ���BmB���]�+%D��Ъ�U��+��9�����N��u�XzK~�MD�@�x!�%B{jqZ@���~��O
4����N�d?�Ϳ��H��{��h����Z;wQd�����=���Lf�"�
Ü(�+Z�1�*2x����I΋y��kxy�_��� \��?�ib�Uo��i@9�S����C�5�$m��Bܥ�GkVSÐB�d�[m_[�WϚ�S��ROϠ�nB�O!�ߦ�'�֘#%����C	����eE]3��V�&�=Qf�4=OS������F�,R �?�v�x����2�t�����ɌY���~נ+KT����}��nZj�@����}N(8w]�	1��Gm�eVʯ�K��`�R�p�i��QM,��A�(C�sX��i.33O���<��3�\e�d���f#/*��Ђ�n�3ZR [ב ��l�e����q��uK��׉�Y0�l%Ų*09ANh��r�f�0���qԋn������
�KU �,��	ȰYU��\~��ӡ�|��j}���hb�@������^Rn
����f����u02��K ��	����tK�܃�J~T��Vi��^T찣?}3�b�A�1���dLٗ�Zԉg�T��MB��W�7G]�^���d@[s��l+`�R�_�.�9�㩸�����&j1���D[��8�햒xKnp��'rl���cF+#ݠV3��ׂ�{�8���"{.��T����JΨ .+=���Q6��B&ۆf@|Td�WȽQ�r4�K�4�j_�j�7��#��Ѥ�g�<'h7v�-��.���	�CP��l��(y.����J�挵$���{J���L�a�2��Is�Gw>�s�n�Lѥ��L��H�Λ|K{�x4�J���+����c��kEl��~��s�6	'���U�dM&��=�5Қ棉�!�܇.<'[ttO+(*e��E��7�����M�G	�
g����K�v���S�����a%���q��*�"���� �[�|J"�ऴb$�'xa��z��:�m�S��1�B�hm�Z��7�=�aF��M�f*�O?��D*�b� ��_w)}(��%yzVy���z�%�(�(A��b�k��o�B�͆�C�.��)���:���;Ӫ@�.�ɀ��w�'g_���z��&[�6=(QC��(�wX^,��H
ځ�l�4��E���*%8W*��ߠP�$��A3��H]�>·����#h�X�k������ȧt������P,+�8�4���`����!ѡ�v9A���av�L"�$G߫ʺ�v�q#��;l�i�ob8^#ŵ��wvt|�d��+Eˈ�����عj��n��bH����_s��,��OD���N�pm�� ��K:�9\��Q��Ю�B5ߦr������.��~���-�g�
~���h��@!]R���S��	��$ �㐗�D6�́����[Y�F�(����x���e?Ҩ�se��0�Үh6��%�~�"a�:� �";rS{��)gh��S��U����$��n��ܴ�9���\MK>��zƸ�|M��Wi�9��@hc=�ۂ/�4&�%�/M�ثe�f4�p.��,�<��x�|���p�}���*�+}�r;���Y��u�aZS��T,
N�)���/�L��:0��҅-+0�
ن.�e"���C1A�"�y��c�B4�~c�
��m���b�9���2'�q��?�T�튳[����p^��Pe:x��d�G�Eiy~V��w�U���O/*���"4�4��{Li�T�!��hj�Y���~�	/�h�`J��}r��*�*K�_��^o@��n2��t��M�����L&51�%kH��f��>����X;T�Nq}@7ݢy��9�'-���	O ��m��XF�G��`Կw.>ZN�]')�*HE��&��|U��D>�'&i��0���x�������hDDd��x�Z������'��U3�����pd���Vⷦbw��)��G1��J��p����3#�H�\��eu�{s���s4O���
�h̕Դ�Z�I�/�z�D�6מּ6ƛZ�0��
hD����u@A�lJ5H��t򚢬vzò"KM�`���K%C�'�e��s{��������"C�J�K�q+~� ��Ņ��.O�u�|�Ґ�E��4,���Jܸ����v�8{�Ea�U$�j�>+��NfD)T=��X���)@����;���΍��f���T˶�]��T~�� n؛w5܏q�$e���8�����t��I�
��Hx �Nx;�7c��I�?�۶���+�k�ݡ~�D���k_�~�I}��U�y<��M����m�.��>�լ.���L��\ݚo�pn�������Ѭ���o�8؟W��).җH)��K�p~��a���xZf/:ot�JN���P<��X�]�M(�Ȍ��]y&/t��*�]��z�g��G�7Î!�<h�I��?��V~���.]��Q��};��� ^(���n��@��;h�?��?5V�E�=�B����O�t�O9��3O�/�� �-R���,��d�4��82�ʕkY�:��B#�n䣔�J�����J9�č�$e䓠��dЖx��H~�Ң�<��.���p�?2P�hh��T�[42��r��+�TS,������=��fkۘG���l�C��dc#�X���lX��Hy[��ߞ�+��#���d "�@?n�l�x����8���Ⱥ�~J�ܩG\�{uP��MZՌ2�g��0\����Pd@�7C�q�ܳ���Ũ��=@��ks��fYI�<>�u�4�4�_�Q����xHzf�a��C�����tL��K)�ۨnJ�@�f�9���C�i�]�!/r��U~Ϳ�[��p+� �^
�ˮ�dU�T�(�g��U�u`H��Yv�������ғ��qfa�[~!�	j����\�p�j�H����ɝ5�Ǘ�Wj)�>O6�C��i�$uT�[SW��'r�����lw����b��z/"�ԥ�H�-��T�?�l5V��ê�Qh����R���y�ӯ[��cy�/e����[N|F�����BQ�n��~�,�%��ݻ%z�n��
L�DF�̂��(�n�r��)Bn�I�a�_�3^��g\��q\���ې��%"KK�~ ,���K;RE b-��e��i^�{�h�G����f\�Ob%n�e��71���1��e�4=�P\v��t�(m�E1,��h��]3���	�,'+Rm^�!_��޾
�+�f��/�_2��e����v��Uo�**�gY�#u-�W��S������^.�����l��R�f��*�W�c��[p�ԑP�RQ�-P�Yh���@zР�����yc:�^`(�':y��R��Yp,�^���Q#PnT�~n֙Sw�_�%��lr��~�ޖR[�\l�w����_��R��RՉT}�@�������k:�{!]�	UU�7ꟁV�7�����G,M�e!<ոի�\E�����t5j�(c@X��4C(D�0��	��Hh���f��p��5^�&C6*��	O�<��/�!p�_��\�%@F���w��R�{*�{��B&�A�R/«r��((�at�xV`Ub-p�[b�1ׯ�Q�6��ې!F��W=)�$^x�Xߜ�E1[����ԍ���l�!�ia�v3�?�_���s!{J�Mǅ���yhX�e�]�6�V����Q{��u��ή�]�9�%8�[u���6�_��w��6l�g
���\X��A%Gi�i��C���:�]c�����hh�3��\"6�|1m-5�0gj5ae�W��L�Xd:/���~Pc����! ��O���'g��-��Uk�ݶ��z�m�#��3.^��[�J�%7tRq�c��<� �5!���^Tz)'SH����5]`;�<e�Rl6T��V�J�����s��Zǩ�?BW�o4A/��
�_6qz�MV�L%I����=Z} ۅ,}�Հ�_7���Xֹ>����6P�Jȫ�M'�$�OϭP���
Õ@��i7��k��`��s��Ш�J7��V<�T ɶd{���}�ds��.�t�ק	-t�W<��1�H����ۭ�YfL��ٝ���v�I���}�(��X���t��Q�13�o<w���͊p���t�/�B�f:rL}�E�:��:Q�*���Xʃe�u��A�-��]C�x���M	B����ֳ�	�-����K@�BE�Q$o����ٗ("V�l�:�����������%���q�9� x]�chÆ_��D��`]�r'��d���7���h
}^h�H��w�;��nG��[���j��=O[�|n�E-�P�5�P�d��k��[Zz=�`�j���G�^�(�l(1�v͉-���dKew�u ���
'��D ���W��eߒ�-���)�����d���-���\����[�I�pR��c�)�ݲ�<�c�{@��S2����'j�O��&^Ź�X�����"���	p��nf@����$ǒҖ���;K���zy.��{���_k�����B����H��k=Щ��%�h�k����;@�5�gP�K�� R6�j���흲��U�%_������@�~��%k��7��ݑXX���n�������1me~�XsjN��V�����!��0�{7E�� �!Jj�E�(�C�,Y���X7xf�^k'{�>���`Y���oLL����Rk�S�(~A�L��|!k���Ҏ�/���Q�
������Gx{���h����A��@�Ċӫ�]�u�����\,k�Ju��µ���>��� ����w�D�"ƴZ�[��É{�(��t���#�ܑLZr��&ֽ��.e�+�[.��Y�d�?i�`'ccj�y�xU_P�V�b�܀�er�*{}�_"�9�[V�� �9�**�z��>6��DBX�塾��}�&mS-l��ݪ��}9Al������(�Q��N��6��*!q�=)�_(-](Ֆ�Ot枤���=g��]��~��R>�
�R��j�B��䷱�[�6�=���	 ���9���ɓ`��9�} ��6��@�Fy*�98����di�8P���T(�WJb�A�b�$��b��\��C�
!9��q) Sp���>�"�	1%�7�<`9������a<�1����� 4^� ���ķ����<�-��'��#zP�յ8։��~_�^[��,W:�S(�!��Ԅh�k��?��
$_]A�3tb��3��5��ɦ����n+-�7(��<�9	v��&ی�Dz!h4��	K8�y���g@�������F2���?h�+Nf�i��g��m���_^�-��]��_#[�����E7��א�vS��i
��SB�zX9nm�G^��D�n7����fo�JݴxK�:oߗ�.���:�W�2�'�eŃX$�1� E����*;���'͢�Gl�/�+���ZE�����k"��(ym3Q��r�Fm�%�� @2�7IW&�޲.����"����% �$���@N��r��85��.l7����0i�0&n��|V��z�]tu%֋/|֧�nDTC?76�8y��\*^��-M�=Q^�6��
.zV��%K��('��ow��M�+��-�*+K��-ڱHA����Qr���������#Z��6Pp���?^�yMmΧ�E:a
�@�=3~��A��7s�$���g����0��̙�D��'zS�������7�Y��%���O���-���[�H��@ �=";4�0XN�/Q���c`��.kL/���iO��c�Od$
�v���؉��A����kHa`6��(pl?hH2���r����;��(*�����T{�-��bi���S�?��v%����?%ٓ���"'ڮ���U��P	kP��Bz
�UJ��c�C�yad`%�����wί�6谥c�����b�$�o՛[�S���`�t�0�+	X��^LA|:�s�.�^���|��}:f`�D�A��L���䩿aw��Q��xY: x�t�8%���R�/�{{?���8p/;���OQܿ�iXD��Yy�7����T
�o�d����޷�Hv��NX�?���}��ʘw����ݮ8a�%��2�c�+OI�ͱ�V�8��ʓ�+��;6�$������b>:I�m���wX���g궪�%�P�i�qe�Ik��W�BwN2RiV�}������E�
U|1�3r��sz8p�׎))nxĳ�)���
��Uט/T��Be�H*�Ed��� /���>�.���ߝ���}H�lv ��:Ƨ�0����T�Q�k�ݑ ?����nb��'���J������f�Z���nAY�;�,~�1W]o+��>�wڋd����.�Ix)��r�;�C��5q��T$��~C2-�U�jv<����pj���A���7����c�)3�YU�w�mj ЇB���S{k���Q(�57�JW��]%WF(��/�Ij)_�y��"�"Z��� d�V4�0xE�q�ײ�b">y�8���a�I����|�ee�ʯ��w<R�82���!���g�''� �m����0��Ee�M���L�=���*L�~rqd�L�!�E��u����4��o�7���	��4�YHJ]b۔;_l 9ZEA�*���j&�B]��vz���C~�����3'qB�Z���|lhOc�5:$ض��i�H���F�ϣ'���9���e�=�x���i���>�2�%ףhC.��)���?��j�9p�,e������� ֥V��C@��Yf����k.��;@���:y��{l���f��C{cXE���x<�SjS����e;�AhR�L������2����|tC��pW/S_�T��N�8T�r2�+�'���=J(�-�X8�e�{�)������K|�"|˝)+l�槏�=��-gW�&͡�(�I^�B]&������io���Zv��B`���20ߘf !#�$�3ݷ4f�ޅgk��t�j����2��Ѭ��?ғ��ԬGdcҟ�${r�(�U󬸸j�r �P���
e_	�{��!�\�Y�V�
��)�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�}�\�$}�����,`Y�U�m$�f̾rc[eR\���?CɆt]a�B���R���������ʥ�+�[���R��0'>�ϋA�����/���;㭤3�r���$!�v	�IL2�����w�џ�p[9�v���t�MQ�Tz���6��M��R&U�֘�ntG;����X�V9���|���:�p��S
�|�beB�n�ؖ[A���#�TLa�T�;�7j>X��<6S�ɒ�ȩ�_��>�_,ڻ	��H'�Nh#��̐'�:� :�2�q�+u�I.�YV��F�pǗ�1(2� ��I#�m'��x�`s�O	�i]�i�Lpm��i���CFAH���Gd!�Z�֙�eHήC1[�db�EJs�_鎇W�VM6����6K}a�U�*���S�v Me�����DZ��`�^�����1� ����W^%�=�s:�CY�}`���+a���'B7���^��P9��<���+-�o�'u��������>��5S5�h��Ò�]Y����6���.�M�V=Ckg'R�U�!ҟ�*3�0��s >��GZ�0������6W�'���/K?���YN������=������K���n}i���QE��Qs:ݜb#�C�zC�HzsB�-K�M���H�����L	�A�(��m<G�t~æ�����.I��ʲ������ЪU��0�����o���<�X�JT�F����*)�������PbB~;�6�����R� *k�|ܻ!����쥿���vD���AG��|���ܑ�D��[�x���Ƶ��\�_���$����>��i|OWȞ�Y>7e���#�<�ج9~����$�Dy�ui���3k�3�C
?>G�9���O�����W`�@��D���_�YĚ����g�Ho�[g�i[�1��<>s�	��T�K14��zs���q�xnbd��[�����u�@���L;�؄������L�S��a��;̞���2��I��CK�}��:*��MB� �5'�c�n���su��P�=�eO�3�Z���O	�т\����Z��賨"f����af&��;�AJʆ�Y�"�q�S֎�3h�եZ��x1m��
�^��順�K�J�z�G��f��E�Lٜ];�
'g�|w���&�-/`,��AV��bh�8ϛH��:���ۻ��w݀��S
��/�z�����\��򠡜����(���YD�����Č��6��3��f��j4�%Ԓ�=������[��jR�:^Hm�P�%h�C�8�)��!;t.�G�^n���fG�������f��F�AJ�Pf?ns̛��UtX�iFi�T~�����
��h����륕M��F����(UX��� �t���½G��c/ 	��M���VWkƭ��ȹ�6\%��>�A1��_k�Ì�E��C���y��/�&�7��-�s��ܪ�������?6��t2J%,'$��pԗ��]x:��6�+yJ���F�����X�k��׶�- �t��`Y�otFwD+�{��o�*��~��ä��Ě��k$;��ld�V7�7�J!�?���s��J�/3��a���C'�v�]��,J.Z�R�nO��4��� Z4���N`)@��W�йj�ƫal��nȈ��L�ݡ��J�{~WEW;R�V�Cn���>{��b9��2�Ō�5[o�ҳ�?4���t�(��r��w]s ��'���MU�DZ	1Y���1`#i������"���/>�(�f����2��֏���Тe��=:8�U�nd�t�'x7��	WWܻ�� �Z�OF�g���>��w��1���˨u�6����:�nf�tP_�`0p}:��u�?c���E1��2��/-��3�!f,/9��Q#J%7��@�
���nYX#	��7ϗ�����K�m�0 �ޭ���P�Ie�[c����x�3o��澹�+Խ0�b܁꓏����=w�k�U�q��d伿W��z���"Jkaq1�>N�#G���ܟ���,%�P^O�P[0 ���ԕ��m--�TF�W3��ԑO��/�6~�� ��d5�Έhe|�G�����Ȥ~B(��N���FK�6��h�U�^Ҁ\;?L��b4#0�+Y����g Hm4�̳��.�숗�1�T~\�7:[Ú�8`f�r1�?�4Y��'�	�b\m,�*%�t<��r͎���	�7���b"���P!�%�b��y%^���	x�m�����|���̪6��H$�)7ֳEHRL��K�g4�*B���A;�����In
�Q�G���/ė:�a���
H�jV�M�/��%��܈�4�������T�A��ZHF{tu�ٿGSW�á3R�F"�V�1�����MQ�,�G3Q��c/��6g��3��N���6Ԑdy�.�w� �������Ļ���Dz�Ȩ��ە ]ts�����ŗ�i[uo9���Ӑl�Z�5�>e��n{�������o'��j���DCa�J#��I�X�>�'��k۴�S�W�Eb�**��Ѣ<�Q�s��0�(hGv_⏛5�a��O��U]᧗w_��V!�q�F����=�^̯�l�;�9K�}>cSȧ5oR�#����ߧY�[%i?��[�hh�wUb�g�f�=Iũ{q�����Z�`Oo2�0Z�sN�V��Bz!��T��c�e�B��E��R�gOm�F�YJ9q-W��Ԅjs��5P|���tiFb�/3'kpR=��9��杷K5��'_��^���W�GR��B��}�{-X%���$�L`D3Q~�����������ݳ�a@�է�ӱa��� ���[�x��=�{7��豌_��BOx�
���]�0r��Q�x�J1�}3^A9�~BG�5�Ν2[�>�zݒ�
E��"0Ȇ*��ۊ�tB$�`a��ɷ4e�R-NSRv$���m,{-V�֪�L0~�ޥD�a���`�ȃd�h�����d�����L�׷7b��p�=�rZ}Co�+K�x
jL#���rIk#"���t�[xk
��.bsD�\�U��LP��Yx���Bs4A� ��L�C��J���ÖNG��?z�����~-ZW�G/s�$��m��+��O�s�2ym����	
�A���Mh~��Z�H�Nh�oy��m�AP4�t9�e�8�}a�����~�����盫�P����"�)]'7a����}{,)n����q3�ۅ���[�����|C����7�A��"D1/�]*�1<�j�+09��P�;�Y|v��ԕ�پFN4�'��#����� ��d�g�z2D�.B���O�zV%^���g.z��A����6��H
���ڿ�5��R�6������+�`+]�,&rЅ?Z�o1r�<��ۻ�I"_<7m�C^P琤�l�K5}�(��o�j�yY}?iE�d�s��9h< �d@��RBh:]e"�TB3�v #|����/K�$c��գ��Za;�ܻ$g�w�<��0Y�<���Y����>��hZ��}�n����}�;����*r�Htٖ�
Ɓ�;r8�r��1�+&���_~��^[�6��S��8f�1K>
��i���c��#����"h!2�!��v呲Х���'�erNR�?I;�s�}����x:Vrfnbb�ԥ2<6#�~9�9e��[�
'nuNc >�lN+T��$g������{�4HG	�1X�A'�c�D!��gE$Q�
@o_s���o��%N��aams+`ɱ�rH��Y9�"��8<�i�
� \�\<C��4Z��7_�cs^.�_a��=���#C�#)��@\�ƲY�&��3��9�#�#;8���'}�9e�D?����HCTP��`Q��>R�=��M��n�C$���u���COSu�Uw��B��9�m�d	 vx��w`���,5	�Azf��幇�;�xc���!���Kd�<+cn�6�Yh6rW�	K:���M>��P�iKs)a��1���>��oǂy��(1Ӥ[�"�fo�M��ו��>
Ľe��K�T�N4��t1�hSk!M�&�O��ê�T5F��8�-����$���hm����`���Qh�"yr淺غ�ڕb�Η�=�2���z���AN���s(�_��`�^�����nX�9�[�I��$�Nl�ż� m.E�;�@����g�����ob-1�O�>�hВl8)Q�DJ�ʒRa~�+s��;cB.��6���c�����h���Iu#��JzLWTJ��^�&�,���N���dC�	;��=6�H�hP!="�x�m,���`j�ɳ�!�o7L�F�9�/�÷�CW�K��s�νpi�8�~00M^���߆ڭx읳 �/�48�S�a���,uM(��5��XI���?2>��^+0�J����A����oU����=nYב.���Ft���V��#R]�1�����hЪSV*t����4��)5���O��3)��/vӔZ�&ٓϠ�h	����T��x�81#	Q�K�E���c8������fAsA�plxik,�+Myf1���<�5Re��Ǝ��:�9���ф��O�i�fb���vן�ָMSU#��:������i3F�}a���PLᨨj֮!z26�q���G���Z8j�JR���N޴~�s6P�C�'�<��t�Q�m��n�鸧bGiq���mAp�&#��rz�iy�\�2�PgG�2���j�.	�1ϦbX�ٔ/��i-�L�k�B@�0����K�?������a琵�7kޫ�c,�� ֬�JTL�O>�0l�Mb	�F'(_�t���$ሏx�i�=Me��@@�b5��n��Z+��B(������}_�΅5�P8X�;K(b�
�����-.Qu]��0�t�g�A�v^
�@�?�A����U������8�"_K�b��n
>��u���W�P*R���*KqM1�Q��#y,�"A��Ѯ�}�����圢�9�!e�y�=��c�#�ލb6x� �%o�������Ѩ67�<��N'9����I|L������І��-䏾5�6I�	xN��@�z�p��PD_du�.W(LMM�� �����a�\ˣ�jw��9V&��Xa� �ӴՒ�,�+���'��|ޗk��4�T[����� 	�wڛɌ���5i��Jx+bG��d/�����Dzl�Ճ[��	[�����gz�e�PЊQ������Vp��Ϻ���ʊ�J�h'\Zt=�8X\�#-g�����{�=��9��Ѝ^�����:l|F����^�)2�*~���r7�iGY(��v0�d&���h֝L HWp����X��~]%�B������g_�
�?�D��^A���p�NO�u�)�'��;�)��qC�|m�� R���w�A�!=1���}4"����r�o���S�V��]�t��5ؘ�ag���n�v����#`$��ٻf<�9*��"�ߟ���hG��9tC �vѾ�&W� �2�n��jñʤD��e����QY�x������4������}+�s�k@֧�%֯�i+t\�����FK��y��� $:��P�*i�����!0.�C�)�'���J�^\�,?Rg�&ǹ�D&�4O��I[��|em��-ئ�;�2�K��4AC��ǅ�����'[rc��)(i�`����k�6�;dɪ�J��T��� <��  ֡��CA��a2���]�l�*�^x�O�Lb�3���H�Qk��e��b��N��D�D;7Q�����dwKMe��B�z���0�U��]��Vo�tw#�}�f�?E��7�,�<V:�]!�r���Q�c���qF�s�,�b�?��Q̻ҩP�]��o�z(A�ՔC�xx�.ܝF+�*&N��B�
\o@Z\�]��B�D-�U]��ά�rŝi6��v���$<�O"�׾	$��xyS��0@i=��\�mJd	]� �>� �����;�y�ɰ���~��3�Q������ǻ
�D>E]�y�<���6cL5_��29]��*5Ryc��F��`���ɨ���]��θWe�an��dw���Y���ON�H�B��N������lI`�"��4�g+���Ȣw�{ ��5&;��_�x��a��w�	\SϹɄj:]�Ke���r溢� �@ ��ś��T�@��˟a��7	���}�S�4��[p$dGP�'(8}��&���g��������H̺�7���Ė_tl�Ϭlyv�Wb�e������{E�Zۚ4�P{Sx��e��2qsH�dF�g�4cs3Yn���I�`y�w�5�V�w���s���)���K���F"�!-����x��t80�Rt\�Pw�V��L������K��	HtB�v��.�"�v�r�U��������.ZCW��^~hJ�A "@3�RC_�K�lj%l�ZbR`��&A^-�X�$�!�u���+�R Z���0^y�����/x̒`���e̥Sm�kH��^�$��a�����A�'8e0z�H�u�&R� ��
�_m�^V�<�.�9���D�Ԏc��b�7&�%s<��/F�uV(�+� Hn%�D��5��QV,�������&�6�U�,s��_irHn6N�y$V�-�癓��L�j{<a���g�@j��'���:��t�n8���v�(��D ۷�k�Ը��Z`VL�c�L--��ޕ�v;ݽ>2�I�Z��*��oG�]�dk�����^��.DlV�)^��N�NȚ��v�M�]~S�Z�"Y�K�+���� d��0|��Д��"�Bc��24�2$�ap��\����H4w� ��	�ɖ�&�s1���p�W��-lh���U�au��,�QE۪�i�*��MêQ�����Y�Y!׉c�Y_�)�:7K�dEVvc�q�8��tX���@�$l�������tf��E�_���y��4�!�K���>5vZ��4Y�5����?֟&�c-.f��L��ާ��,e	(X�}����,�f@�d���4߻�M��`�7�x�y���O������*b�4F�mǰ敌�]��S�D�R�V������ɐ����}V�jB��^�ظ��L>����NJ�6.�f;,�=:������*�U[��5(~2�c6������#]R��qM3����o�9��ܐ�T�f���TjV7�̇N�R�3�9
<a ����q2�#W�j�Ӏ����$�����͠�����@���z�_Z��	���цp+ϭ�m�,�v!�Uћp����.������������S���.�8w6�:k���4�@v�ĦJ˃����2q��"�u��0��XV�w��9��w��=BQ$���E}�,M�ƻm��ǌ(�*F1����8lI�.�C/F�J�3Zqn��G-j�f�;�w[pGl��4Xa[�5�5�����,s�B��z�V�Z���O��Тd�z�@>��
 ��O���6�O`V�1(�*�'B�,j{��U�cP�եM�}�ѣp�����0��t׸��@��`�����7�>� UrX�uk�%�i�t��Η��f�QWxq�됧�A�}����u��㥿U��?��S����N�5q`�vRhI�n�B�����tQ�%�C~�aR���WI՞��֢�	�#�l�(~�VI�ϖ�G��^ַL�#?ߦj٘*(Ȋ��Y��:��~���'f�<��ؼ�fOY�dDo�w���I�!�:�ɛ�`� �W�U(��+���3�׈�2�_���_$�����	2{Q��|wi��I�Ju�'�o�P��{�����]�~���HL�p^����z�K�f5� D[$S�{@���7_F�E�!�	���7d[���aCua���}~3�F�e��F� �@�����7�ZHU��.�>$���[����c��gW���6/}�%2I��:���6�{���c4!h��Oj��	��	Y���3��>�Os��g��I���up!��@��M��,��J��R��%���D�T���j����������3�r�[�����	����q�x�a�;>�u>~،�k*�n~�M����4�<�m;����I��ϼ��g?r��(���R�?�>�^�D��:�R�T��"�����s$��HjD�����Km�qt�s�i�F���d�@}�zS�B�͏ܼ��Ex�3�U����]��#>�9n6�yssd�M F�;�ޞ)�Ʌ}�πƞ(�Z��<��7g�)��n|�Lst����� dd�+A]T��2�L��4)peT�pD6�qT�æ����?e�d�Q���\�.9�tqNtV�)E@̉P�RA�U����i�cx�@��3�<�.5*,]�l�ΓtV+ݦ�b���I��Мѿ��㞨m�K`tK�-,�,��0���?�"�,���Q��`i
�De�V���i��\��4^Q9��nHCtP��N�%b�*JU}�=v&̓pֺ>g�ט�-�ZU�3V���?�]��h�^Ҵ�e8���yK�(��!m��B�8Z&�~x�̻��ڡݿ��&��.BB/�t��#�)|�)�?��忤9��)��_��V&�^�n�B�Y�ޢwK�+��b��{J�O_bŶ�|%��x"�E�-{X{�2�iȂ@Č@[���q^�eĸ�1�Y�C�~*��M�Q)�Q\qI��4�����s2E��� �Uo_�gD�i�^k�k+�6S�:�@�3��HL�� ��xA�X��m��3���!j�GPh?8�J��h�s�gH��&lD������� �l��I��d=����nWp;���Hh\to?�uK�ͳmwm	��=��c����;c�/�V<!Q'Nlɚ�~�E%��Fn��VBc�T,VkA2a��2��B�����F�����  �{�]��sJ�������+&r� t��X�͢w��yїa;Zy�R�U�n�	����6k����g��og�]�������C~�vR��ttךB����q�̊��]�;sk%t�����n��p;���j�h/�l;� ��М��ti����C��6�7!�Q�s��k��+�Dc{�?9vk�~С�e�=\�)��Rr�l�.k��z�)P����v�$P���	�V?�#��j�	;�iA@�n�fGp�1���������WMQ���Q�G�IfV[[2���`r�������.8[��c����4���;稪Z��AP�V9�Gb�+�72���7�tB�S[s�x����FXxXȐb�q�\�������3A��Wna��-��2*�b����P��d�I("T����>�P�u���(K�:B��p�+4q5�%��0�G�&úd�ѧ[��(Kf�3ڐ����剂r ����Kc@�'�WK�q��h!�s˅�)F���P��gE{�5y����}�@�w��E�ʟ��cQrҬ�f[D{��+]��i/B)�S����"��KP��&�7��^�`���Z���.O��c�l�)V��_]v��f�I&�i���fn� 9�N����A�7/#�R�%-R�5 ��Y���[��3�=���}�x-#݀��.p���>�������kwHBZcP��GB}R$uI���������/��VV[p��#�f�8j6� #��$N���.� �\�x��\�
�j2��B}���$$�4_!�5���f��J�����IV�w�(���/	�����0q?���F��p�g��mm���X,�|�75�:��˒E%�`�¢���X������X�%���C���_s��~g���>UK̀H^S��P�[2g�t���&�)��}����pﾜ�S�43�!c�)�}��l��ؠ��B�i/��"�U��Nw��5���oR7�-_�$���Das<L�P�p �'�7�ݒ �Nu�Y�Y]�݀q8f�ƭ0ؖ�r��_�_"��"J�E�L6�TJ ڊ\�F&�d�:���av��b䵧U!�]0*ZzB,���� !�^��兄b-��XW�lN��K>�-�Ȳ�P\��>p>������`�H��&�d�*g�yѿ�;7�gR��v�p���JpW$fY7z���C�)�#N�L�['g�-���a�-g�<����] ���ͳݸ���.� ��?8�b�I ���"�B�~�h�b#��i$�v	�W�[4�{����	�O�,"�Zڒ�g�@���Q��q��+��3���*��v�g% �Z��g�4A��4����
�rYi����S -��h�a�#SM�y�6���c��%{ 7@��!:�A�;��PT^5�ߩ4ŃZ]�~�i#��=�?$3epn~�(iP���V��}�~f�\���·tW���T�՛<�T�����:��W���$ʔ�M�r~��y�z�������g�+*	��3��~Mpw���n�� �nZ(e0t+=��}{�m��R�	�Q8� ������?S6s~ʴ���'
l�4�cp��B��5E4�����$�}J��Z!1X#�Ѹ��Y�@���ܶk�-TD��K#�48�GAp�^� ñf<03�C����/ޙ2�6�^�7LuV2��p�&i]�j+W�2\8��N���@���ģ���6G����/����B�����!][��XA�wV��Ҟ�������`��-��t"��|c�x�<ȩ�_;�j��j�']�����)�?*Bn���H�靿���r,�:w�)�7@��Ȩ��w���I>�łE�EfZmLfn8$��aa�.��wFYƞf�*d�Gu����Kj���O�'�8�xR�㷆�Q�|} ����ջ�|J�6cE�K�P�`�Tk���g���E0���Z/c��m�}g��koŀ��M�����@���X.h�b����
���+Jc�u�n:g����u��`������5��P1��a7coA�F3"�� :FG��o�gw�`��N�O@pi8�6�!��8q֟��I��^'RK����$����ߴ�����֜�=AN-�֏j��jSgL���j.�dRK��:W��z��aǨTg�Y���9v�Y@��"��^Ou@��A�y��nT׵;����o:à��Y@ 0�d謣�89-L�Խ�4P��n�m���07tV<#��)b�GTI�*�ϔ!TM�tj/#���T�6��~�J �dI�Y�<5˫��x���q*SQ��)�;�j��ќ�f\׺g���]x\}�la��]L
#j�yQ���cN��n��˥۟L$b�Fk"m��"��ƪI0�~` �s���Q��/;?q���`�[���o;Y[,�#:x�&V�2ο��뚨,!���w%v�;ᜬ�T Y�0��5>�N�\�C�lp��w@Ѕ_W*6�ɩ�����tI�S���\h�lF�u�.�����ovh|^��F��B�wБB��N�8d��&G)��I�f��K���V����^i�.��@��=�i�N&ZM���~w�*�؎_��r}k�;,F�OF4pY�G��˖j��t�.
%��f�ˉ��&�bwv[�� `�#�!Ă4�{Q	���X��=����m[]sYO���I�ւ�`��'���W�o0��)���v�b���3��J
,U����g��`�u&�E3�h�ȉ�r��a]r� �t���k��b�r����n?x�M�k8(�����4��A|/G�Js��?��-`Nĩ��']�0����K��y���1�"��=]���Y�!Ewm�E�S66�~�?탖�����of����!L�>���-2e�<������م<�� �rn����}b;��zf�gh5�@�^ʱV��'���V7)�_/{�����e;�����C�)Z�ؼ�(�5��lڱ��i
��n"/d�]�h��-�P�P&�i38b�)M�xZ��556M�|���L�x��.�~��3^�����F�^%cB�Vi�4�.A/�W�������	�an���I�%9=���%'�%�F�o�K%S�}B��(U����RIE�}A�(k2�Cq���TL���`JS��>D@¾L^�.ֻ?�NQ��B�qo��Ir�t.��_�˔�b}�ޱN�A�#t��47\�bg_�Y�'a@���C�₵X������j��D�]��WWl;�����ܛ:��X��S��T�y�!��x��z� ,(��1�R�$=Ti�%�>�Y�%L��px���K��c6M*u�xR���L֬��R��(0����
+J��Um�����.3k�*�2<m��<KK��ͥ�8(���\��o8
�%O~�8p'k>U{[���CU�c�Z��V������(����h��ـJl�yV'��L�z�צ�=�W��|�b�l��.@��`��G�͗/|�_Go	m���=/�{i���"qVR�f
UCp����
��`�̊�����g��|IXFؓ<z���=��dc�zٰ�`����h���m�)�,S[�8 w���d���r2>�j-�=9Q:��.C6Gy�"MNx��������`��Ͻ�Yg7Ė��/���e3�LW�±=��k�ܨ�H>��) ,K+�݁�Ԥ�a��,���p���|��F���sˮG��CnF��Z�^�a�����O���$�Lm[�I���|��Œ]Pi���ZI�����[���uVO����i���n�j�@V�ֹx���\}/5��`�@2e �\*F9��CWh����t�f�hh����S�z�ıP�pOn��O3����7���'�bT�4Èc�,��݊+�$2����� ��a�Z� �hҬȝk+"�o�*t�� ��b�M��YC���5��#�H�,GMn�C��jB#�F(�"���W��͎�^amq9���S�Uª4�s�o:�����Л�u3�7�)�u��&�v!��~�-p�vF}s#meݢN�mo�	;�GZ���G�p���m1����]	�	�ǹ��,e7���߆
&����ꉱ�G`��8��y�L��eԪ�"��،��'Yj������eb���NPL>��|���3,�4K2Kj��[�`�4���T�:^q���m�`#Sf�i�Q�o�%샴���hۀ,���i.�fM^�@E;e᭙�X����Ʊ7�R��
c����Dqsp�l����@]
�uI�Κ�B�������Dvn�v�>��C�V���|D�P�BlTy 7/?�C�����/�ԍj~��[��tʝEe�0�,�uA`���f����4%/^��̻.^c׾(�Ǡ:������4I�8����;�?��,rGϚ���\S\�o��q:�ªCEį��
u%a��N�y'$��Im�
����e�\���F���LӁ>)�h2
�$T�����i:�vJ��P���Юo����A�bլL 	ڬ
��"pt�U��Ym�>Q�J��ʒ���W#E=�69:���`�%���2qEK�0Hq �₳8�}*6S@�7��P>��|x�-�C��[���Q�U 1�v*�]�,�8�Ӛd8%����Ii��k��[c�ԶU�qК:b[��h()���~�1��J��	)�����*��yI_d���rD�Qe��ϊw�^�n����B���۾����(����" T�İp'^14��_�1������{{���N�+��1])S-��R�R���t]�t��^��S�,K=���Ծ5[g��9�'q5���mB�Q.{~�g�nh�&ϲi�����0E�MK��a7E[!G�P���a���N�t��clG�"9�q˞0-Ѻ�rwn�[�[z�׀DC�'����;]��F��"σ�}Mz� �RGH�����m4��(�P����R\eG�D�������T*n�|��(�
��S%�����R�{n���t�܍��j����Oa��H�3W���Q��PDGj�DH#������_&��&�ǟD�B߄(@��� ��=�y�s��v<��G�(bHS�w�53G����/��_O�Ի��+��
4���Ύ!XT��NJ_Y�^�H�@�G���J¶��`K���r&�_3=��{��VL��A>]�ӫ�����v��>��DL
�i6ZkK�T�I��&���C����A݅��)�#���q�\�]�{���h��d^Ŵ��#�l:��Ǣ���T��{���.Yq���A�*>�ڌ����V{�c�zhGĚREc�qEȋ��9��t[�޼�q``>�1P��_ ��؝Sx�mߦ$? K2;ª�1��y4 TBܦ�6��"�C��`����ќ��˹@ݪ{bk�����M�g�yo|�ĥ�4�7��Ȼ�����~�1^���(x�}��W�ÇT�L�rD�w���ح��b@��{�Fg����֍�\Ge�C�j��
U �nV�X��|Jw"ϖ+��
�c�l��RQ$Rn4�zt�=�1����Ij�"��R��V_�if����oZf��cis������E��H�+�u�utR\�C�_��+$��A%�6��A��l>�;���ŀ�8W{$XI<'������B�l�:J67�r!4�VO�ܙ�z�R�D.X�����W��S
�TK����~e�{�����BL�z@�ny�V	��o��OÉFl��|��p��Q{�)Ts'��B����?�2���l����;�g�\�j�-�N/,��JL[�`�r��9�`X�k�I�H�ԥ��;i)�q�PP:7պF��`�Q�`�����DUtQ�H��*��7���d�(_L5���l������y�?q�O�qtXt2db��+L���]���Ɠ�)�XR9�BP��T��b�y��4GP��R�����e+^�j�mKs񨦼΁E��[��;�M"�����+���S1�ƌ�?���Sn�3������C����Ik���`��.b��gr���B�A��<��4���L��TG��P IP<ӥ����1F�jDi�K&懫�#��̝zR�Lgzo��*Ά�>+�%�B��q���-U�Hs[aҍb|HC���ۜQu5,:2���B��|����c ��?�x3��L�y�a�^�� �Tx�/�B�ҵ~ک���.������X��f��+�:o8n§9v�ݟ� >�];} ����}������=*�˜�y~�W5��ݭ��&י�6~h���8J�W�a��%��� 9z�l$H�h&`�npE�̧�g�|����=��l9'���i_?��r��b��އD>#)��T��E{tL���ڧ)[] �hs��"�P�_���@�:t���3�X �)+:K�X��S�_�rL��ǝ�}����e�+���g{�u��ei�U۴]D��W�w���?��A�?u"�8��@c$�������v^Ş�k��+�X�R���U��K?��?0��oH#&�J�*�;���\��^h^�څ�읝x�zƭ��LN�w���n��}�W:4��L�: ��B~ Q��$��ݏّƞo��ju=3��3&���{�qӍN�p"�3�>$r�J��	�Ə�c �9��XʤqX�x p���츝.yS̆�B�nGw�a��
�Э�#��f�����M<#�ɑ��b�b��§�؉qH�dZ�?�ao�l08��w�5Y��Y&
#vG� I�z�܌]��+�|�b�5��[�lla����=Bs�>W��*cY͊���Pm�*�kT��6g�L!�L�T�� ��b���ij�D'�Db+?�@�ܰ�8�M�B��'ͱ*��x�|��4l��V2����P�Xf�7$��nWdQ�_��x�j�_R���f��ԍ���'Q_��l�'"�u>:������A��L@&
k.3���X)���gf��P_'�U��x����ɛ;��~C�a�؟	�8�S�n���rL�	�G��<Z�^��GH�p���*�?�J C�m̱�N�,�C������$'�����A�ϻ�守Y�Y�L�V�U�%�|"zO�`��*�&J)���p�Y�Rw��F�B۞��-s_��x+��&�˶pd��F�����b`���@�'�}�"�6c��9P�^ġ�]f%D���X�_�ai|!���p����s��$�e�l~=5���Y���>aUF]A����6`B����Q����a�sE�:��;�̚�݌�XCə:[�*���f�dI���'��Ή�㟘��7��ӿi��r���| zDĿ�pcN���&	����)���={��}�55�࿯��4���'#|��s�/Gp�[*�܁�E~}��Q����Cʣ8�$E��ys�B��5�fb�������i�Q7.+�L�Q�	�8u:��,,�$����`��!��T��s�=�R��h#�yUV�FY �d���Ġ6��x�M�
BZ3|��])��l3�6y�?@���c%x}�ѻ2�)�v����S�V� ���N��>�h� ����Y:����S@-؂T]W�ڒ���6�r_�'79��%]ܨ�-ԩI+{z'��j=k��Ǝ �d�rNop|"_`Hف���>��)u؝����<�!Sakw�a.����~�QH�������o�3e՜�l�G��"�l��0�Rd,��/��-���̦����Q�A��=�_��OT٦�a~�Cu�Y��Rmh)�<�:�.$䤪��ȨF�/s^"]E2�&��^�T7�k�M��k��6��JT��W�Q9�˟��ڡ����1k�0���nCF��9�� M��"`�`r�]�?�O	�-d���D����wE�|�Ie&�^��1�g?QF�s�B8�����ۙr~�D���ho$/�b��+������^˰n'�4쏞��0�u���'ũ1�%&�Ψ�����H��	�+Q����d!�8��w�5���ֿ*��E�Ӵkk�� Ye���Jj�h����,����A�3/PjG�����X�Z���S�����߲�Զ�~�}��y�ڌM���Qeuj���Rz�,$a�_��E�#bY2������-���]��t���OF��/�xW@�}˷Ԩ��<Ј�ƹ3����|'����!�K%����&��r��_���]�BY�R�r�ȄU���� \���.-��uy�۸	���|�y�#��=�y�wHs���7�`�ylK�^#����oqm$����TG�N�B/��G?��Ft��3�{VW���`{���!��)dn��ldx4�����A���v�"������s_"�����ľ-��R�J�ԮK�"�C5x.��m1H�����1�p�aAP�O!��y|T�Ӈ��3D��p��g�	��}O��R_&��TP�D����H/��1J���}̷x�6�)�
���?N'�BY�Pp��?Tl�`���0}���o��$e�]���X�!�و�%�+ojj��^z�����"���}< �����Kj��
�=�2����4�_J�V��(��NM��6zB.-{`p�aW�O"��gU$i��AtD�%�E|t��V\NxkӐ�c��ّN�-��ۼS�Xǚ�S�.(�VO���4�.{�8��;�-�,!��s�UD�"��?�'���q��+Vx�C������o"3^p?�W�g�)�n�-1��{�ۨ��m��_�aȦD��{�>o�b�j�i��:6_��G��.e�H׸���M�D(� ���(3�5��-\�K�U��ZoU!�9���l�#�e��Sq�fIx)��bR��l�`砋���IB�E��ْ�Qဒ҉�ّY�`!ZW�j3y��]�]}�zS�VF��������K����W�Kk�~�y�e��_�Ɋًr�0I`�j%U���p���?a�'�[|1p1�Q>���G4A7|��6�8T��Q��A�ފ����W����H���>F�kH��9<�+�}ah��)ɼ�pQ��=���?�/{�f*�McЯϑCs1�l�Fi
��B�F�@�?�XG� ��7(�-�� ����`�5SLڣ�nӫ��r�"g	�]v�����7|k��Msͅg�zX�J���(I�ySX�j2',��/c �[�j���0�e��}���D���1�3 "A$��P��Kmg��r=m�۶T�`2?Nǣp�6t2a�«2<U��Q�ّL����kO�Tɿe�&��d���Ў������L%���S<F3+z1�oFY�r(���\}i�&��������x���n%�#h�
,�R[j�{v��ν�(�����\�ǀ�N��«���[�w�>e�Q���1��.+3:E��&���xF��7�:�V[σajn��=[ܳ����=��Q��j[3uZ�;��#p�v!��n\���Ev���*I-*� �I��߅��.wNo���{r�6��\�?�5i}tG��`K�KJm߯&u鄇��s���ۦJ���*���9�Xŷe^$�������-ʛg�Uէ��>&G��+��6l�|�KTj�՜���c;Q8��V��֏�K��F�^��Vr�ۇ� �{VQ�̉Bi� ��S�D���QM�/F� 8��3ƎIcȔq�E�IK`�M�<���ÿV)G�]O��C��5.Ѐ?C C�<`�����"�C#���<t&@�ڳ�z��-�;��]���-��O�.n�U/��V����� ;�L6�&��e^"}�'����э���魓#�#�;9^w�q�Jbvr�h�+��?���Í�\�Nx&�o�Nۘ7͈����L�*�)F�V/��_���3Ey�
�k����܏��Y������F�қ�8�x�|)���+����	GO��\�)0�Q�Zr������]C9�@cTF\_�)��41ۀ��B;�|�̿�hP:�S���2�}lxG!KW�������@�Y��|�X$x�l�Lu#���ҏ�g/�Y�.��&�2�A��U��D�+@��*sd�9l�����zoOܶ�����A���ϼ�a����=Nͯ�l�d?^���Rkv���~(�Бʭ�������/�j&y�;��L;TC�h X� �Iճ<�	_��H���:Z<?����6=��'�,���M���5�)�58�2gL��Ι?6�HLwi@=Z�AKA���
��3oA��T�[�)�d�� ���57��ă�(���<�B$b]�~;�rÛMI_�'q���޷��>01�+䎛O	9)I���~�"tҐ���z�|e�1�mL�2Ăr�	9�d�"����ݦ�׵(�MPg��z���z�v3T��űl�k���k�Wb��w2q'ɿY�G~�GZ�dûw�A��>�??�7�3(.HtS�E�Y����%_V2� ��jv��De�� x�	�� ���,U5��܁Bt`�x��:~�lx���<2�36�Te�B�Pw.���
3o>����t���V�n0|c)Vğ$���׋����fElf�%�]�x�@�;�2�}X��ҍ�m��ޚv[��9-6
dڎf]�Ā��,����9+�(O�M-��h��� ��7f� (�q;�v�26 Pm�OEh�G������lؽK��])2&��$��J��F��K�|��S�Ht��F��<:S�
�e?�JS��
�10ٰ\g����ZUYgϡ�Q�\�N|/�Y���YN���/������b��"��ʵ�OG:S�x(���L[���=����ӽ�f��h(U [�S/�:t�����~]	����0h굡�����SR��T�E9�sˈ��`����L���n���݇�E�1h�'&���7���5�g|�4�7��s,~IF�"�Jqrg�|�e��_��v�w��z���L����R�M@hF(�뙟��SjoX*���$G�ֿ	¥�^8oD��/vjel���%��C��&�o!i�v����� ��e����|��E��Ρ�G��V��+L;z�;ߩ>wT��u�x��u {�0+�w�����ƫ�M��m����&͞�ِQ�]��/�~i�cUP��Ցmp��п�ʶ�VRs�ƪqj�܉�Óq��9>`2Imylm��;�Iu��1ۗ&����o�fkc���x��C����[�o�5�\!�a�������������k븳�~]�X�<�Ȅ
��pI�;8wi�7ڤgf��A��*UI�������~e�k����Ӗ?q8H.��U���pޕ��+A�y�mXh��Xv�b�[~�D��4���؀��m,s�(���9�_�nxRmC��D�Ľu�ho��s�ӄ�U�&��U�/�G���>` !h����ÿ�X���pd7-�F�#����X�&�3�� 7�4�*�^�F�d7���!�b�7v��J�#���'5���}�w�cQ���<�3/G�*Ć�M�7\�7�_�_	�"����-ҋ����:�Tj`���2A	�,����c�ވ�[z�4Dhx��Ⱦb�=��&�Xd2R��a���>V�����AX /Hڜ5��~�&<{]����f�S,"����9ťBoN��|��s�!,v�� !F�gD�������n����G������1M5��5m����@�R�֣0�S���o~�a����bfe���ff���Xs�M��Y#f!�/���Y8�Jʐ�R��NT.|��P}��H:	���u�ʒ⢕N3Q���K*��k��<�iڱ"ѥzB�ē�ֈl��-3��0�A�~1U��w����������h��2�dL�\)�������-FG2c���b�:s�G��5%���Lp�J�V�`aDJ����!�:Ԉ2����K{y��jfI��#a�A�:5A��3г֬�x�ý��&��_t2M�ޖd�rCJ�ox������B�#L�y^ͻ�ܷ����t�7�*X�����9ː����\|!%�bXz�+	��{�/OQ��ȃA������,��Ri���@+�{�"s�I� ��&�Xu�r�m��C����&̭�54�������p�1�E%�O�~�%V~OϣfڰfD�chu�k�#�H��]�>�����(N�T�����	�jS5�����l1	�ʈ�F_o��x����_�7�����7�S `����R�"�7��k{���A"���\��cZM!Y.ĞҒ�r~-���1(ef*+�? 61�0N>��;�Ԫ�z��=���b�����!�e�eU��<rtҔKw ��5�@����9~Ĥ����3t*7u*��0y��f,��aua}�,1�8�$<���%˝�?a~�o;���'�ʎ^��U	���,�����f���6\�b�I��AjF^�{r E�آ�y�Τ���X�Y$� E�G�y?
�1Xt[3B �.��!I�S��Ѻ��Q�2����@�m�$��m�׋z� Q*�}c�_�	�Q/����&@���BR���|/k}��Z�8"R?z�R��Ak�
5�v�����)}A��V���3��S���f�,sv�/~��p,��?��d<�H1��k�%h[�,�+��O�YD��L1s����\�-��U��k�+��g�@�j��d���!���0�v�3���d'7`��BY��)�Q�����O��$��x�����k�؀��W�7�H���k��(":o����W�9����{���߶�$`#(u	1�r����ÝOXƴ/F�朝p��y
�9S��蝞{��	Q�- !�ml�}�a����j)����p��2!��!{+\�"����v���a=���}�79W�FL�O�NO�_�^n��p�N�r_P����7���q8�����	�1���̄8�U@��C�F�݂a��� �xک�M��[�0hllų_z���*������5���l��Y��C�ˎ +[,���C)wMWٷݧQ�*�t ̪p|�m"9�"�gφ�ϕi��c�<��(��f|L�[Wf�+��ظ�
�u։'��3C����v9O��*�C�c�/���)v�q.(D�
W��RE>�����|J˟�ޗ#�袿�G�~؎�� �.`鑦ҁl����k��MO�1z�u���eu�aEZ�"���w"�i���v+�;A�}�J�Rg~BF' _��g�Td6����,�WB53��d�L�4"�����
t��
3�ƞ^�zӜ{��H���o�fs�s�cO���]X��/t��Ω?6R���
�D-��8�y��1�Nԋ����'"��"�z^;q�~ů)��,(¡�W����>�9QI� bO��zL�Қ���g�#�*��b����'0��g'��#PBM�e��J��yY���`�
�w�'6��D;il�����/	���	�M�5�44��?3/D��E;�k����>�z3�1Ë�����#Z���!��}�4)^���80$yʌ��j�\��Vl���'�8z������4:��wWZ�ʽ���&as��R��� �h[9X�D*cl9�\&�-k�g��MT!wD!�?n4�����74�N?^g�v@z�{#Ψ�$���!JY��i��z�5�rq!/"n�T5�Qv����zc�>%:�O��c9����0֙g�E�PDś��0��re�����w!�X1��"���v�*�c�͌�G��5��K2C#����1����(���͗d1}H����J��۩�\��eY%�i]��8�ޝ��i���=�:�zK�!��j�"3��X<z2����q����$��Օ��B�4�h`mi�`b��[Ņ`�P�#*�:c�3CW��B����K�;�:��.ayJ��+Td0��U�1�A"�"&k�U2sp�Ѿq�yQ .U��$��4��oSL�N#�мf���3Q$�M���	e�́dì�@j=B0�F|��o�YCy�?�ilU�31���!LH'm�U.�����3��*�JN�����R�Ԩ�u�Al6�f��ѭ�g�YH����$�T�ڌ�(k�7�&���K�>��7�=w^K�<�����a%,��9V�g7���w_W�v�;��7t{J�	v[t'�žpeϥ��ީ3�,jL �ڎ�����P��1�C������Aٺ��Ќ��$/z�=�O~��.X6��*������u�,�3��+p��\1>��W���V���M�G�~������<�c͏�v�b�8?��6謾���1`*]p��iO��� ik��v�� ��������/�cz�oFTԌ@i�5,΢W�9�仼S����lW0�Z�Kv�����T��	�.�n*�[7�v07R@�94Hn�"�A�o�Ia�	Ɇԋ~�e���
��/+�����
4ஸ�Xa&=�y�����ꅆ�A���M�v�!EE�s��d6f�����j��#��';�0����Ρ�S�	P/��/����]���=q'c\g���3x��*�n41 �|�����p�}��D �T�����R�m9!��i��S��x�)�L�l�s���V<��+i��,q�-����о�R�g���z@\�sTx��M���礂�`��t}�.(nI?�O6M��!�xxx���'�^��zoz��> Wy�f5�� ��H�Ҍ����J
���������0�%����,�h�@� CZ�e��6����d�&t�|b3�����Ym�Qj�J3�>F�V��e�}y����? Lt��s����R���%�H@���V��Tmu���PC�W�(y����a0�n)��ww~U���@y(�.���Ú���;A�^~�G�`q�k6�i�:�����#	}m��%2E��"�T��n�����A�(�	����޽�u�D��+_X˯�X�"��":/��,�*�'�������(�T/r|M�T}�_��{�1����ϛ~��b�aOl���1ͅ>��Cm�*�����dW�?�@$Q�ҤC2�@�b���a�!��u�x���.a{s��Z\C�X�}��t�D�>&"�F����5M[3�X)ke��!3�>p;��#{0��Kj�2�m���;_�@ٚc왝5Y�qϙ� ����]��q�1ˤ<����[���N��P!��[�Ն%N��-H�]��V�0�GuE=~��2�'�����\y�!tg�{��y?dc�2�X���C3��͢��S=r�����V�{u�b'�琛5r��+�����b��p�{Cմ�mw��|��!⧨��Ď�o�tG�hPf����ehO|�5�@��3IL�g:���ޅ��v?X�eb�Th@�?+R��࿵���CH���lrM�WncIۑ��~Q��º���5)a�B�S�4�7W�S��jt�Z<���\e�!n-IųM�I�0���d/�)k�ׯJ��@M�:,��	Ü�`z��d(�L���	� �i�Z����ʗ抛K{�(ϔ��"��u�+鼸�,�q89"	fd��Y���#Y��A���OnL�����]��pub�h<����E�v>&C�]�6�2
��tn�5DF�6Ȃc�y�veh��	�\�F����ߐ��et�B��$Zm�Z��K����9+�2����x�G�H
������R�Ү
 �^���t+��8C���:㶧��zc���8�nx8z`��a��R8T?�v�@���kӠ�����GK����I���˃�n���m���z�C�n0%�j����ST�-����/�Rv��*��)���c��o�q��F �����xϼ٣(٧��l,
�� tjk�la O컟�W%��G��f��e/�i�[�/k��/��̦�(Io30#�D6�8�]�Y��o������"���,h���!�$xo�2������-�t��(*�N��<O.i_k�o]RZC��nm���2�����VO~4���v~���̴�M�$�f]'�~�x���Urb�ϝ�R6ՠ����4������JK�
0�a�+wj�mEp�p�2�cYL��+!��BZ���$.�I��tO%����&����U�>�mln�]�`��N^��hED��"�en�3�ʙU79���W��5ْ�=�)US�˩o9h`5�CA�%'���x���Cz�xJ-�Ȍ>� �{�Q���`;���ؠB�Æ%��wƳ�����"�e;h_"�j�[�ź���66($�/���	��.ln�')�ͱ�jSF�V"�[g&uS3��>�ޛ��X�,e@s��T'W[�e.�O�/�mL����b^�umR%k��;%,�PVV�����Ů*}����Z�q�2X6��q�=F�������72���O�e��I�zPh�~���׀�B�s�^5�\ IH��8`�0���ka�1D���F+�̦�%נ�� orv����@3��*)���A5��a�jw�E�C�HM6�J>�@k�w��3��:F'f�N�[�#S+������C�$���%�{��� �<�1�M�;�@~FU ���;E��6d�
Ō<��pp�
��p�`����	0����h�ЊzyyH)�෍�g��mr�[w�č�O>�����B�%�]�����6�W���Ubz��w;���O�2a����fg؛��C�d� ޾Iȼ�2�Ε��9�$ϑ	���qVZ��f��N:z�b�I����}��+!{�
5|a�u�~�4��z���xI��q"�QZ���6Lf�� ڽ�]X�R�&c�'6�^PYUr��MAƏ��u)��+�>`u=�6g4W�c�ո��%R.�G��Z/Z���ChF*$n�t�A��'�Ai(̐y9�47b9
�j�.�
k:���Ď�vs�t&�{D/-���9���]��B���ƿ4��RUr!����UCq�]_bR���&1vۈ$gDr�Z��k�0VZ4hďs�C�ւBs+g�e��q7,<��R� �< ���ݷthi��x [�s�7K(��_��K	t��+�g575�;��e�g�:����\��� &� �{Ü:�-WE"o��1_w�	}K�
H৤����h����1�;�H���V��B���b�0ܯp�x��-I{�֛���ZU��.���3��D�(��D�l��`HqO�L/`NJ#P++��.\�	�������=;F���}�Ծ�Z�EU��m�,��|Uv><G�~��2��$��t�mU})8�|�Ɯ�[��J|��E�e�u5��m��~)JR���!,o���u?��N���Ty�q5���Y�h�/jty���hC�� R2,��c�\*���M��i�F忙���T1~����9���)��+�^���1�LթW��@�M�ew���$:4�(�k�Җ0}Fo3K��B��o�W��n�.N�ϾhֵzMlE����ǯTqf�v�"�@W4+��"_�1�`ae�Rc|lY����喝IT�^�?��w�W ?����w93�v�8������9R�'����\�[V`�����։z����y�kD�����,b��n��#(��^�|b��_�7�EB���>1�9̣ZY�(F��ɉ�1��g�Ϛh���oϽ�������ww@��`�n6N�������08y-̶��X��-�R�����1���P]�QT��\yYS�~e;WX5�_q��iU�R;������0�ȈSj�&X�;�=*e��b��Y,:Z���r�M��TrLP��Y�[}n��K�g3�J���3i�0�Z�b�cMNJF6���r���M�����#ߩ����`�B{5�OZ$�V35�GQc�l�:L�����St�=aң]��%P('�J�F���K��'{�?Z�"�`�`�)�Y��'!��	�h�+n�U=G%���H�Ԯ���Sw~̠	�����0��铠��r��iί��4�AE%�/ō�
x�c�o��i��#)A��?���O��AV,f�ǐw�
[� ���=����Bռ@��i��N��D�<E߬ްK��jM{��F0�)���{v��4qAu���=���Ƙ3��&��l��*����{�⁇���l����(�>(	�d�![�Q�d�G��W���bPI*֪Z��`<@��78�㢦�"�hr8��%n��Ml|�n��h�Jȣ2d�$�x+�c<IvJ[	�1��-
I��\6[<RRUM}��s��o�`�h&�]߽�f��S�k�Q�]�����XĠ7�fb*ѳ�-��+Y�!�f1sj��+�`�	OI�m�
���z����K.�ΰ]���@ޕkk%���i�h������e��:	d��W�CqI�{��ՐΆ-���o}�7���������w� a�lo��/��C8�f=
����h��r\�Z<�L�Ȋ����!7����j��tC~�K�)b�l�0���T�?��aq�W7({���{j%�;�D�CI��0�Ĥ��8]������ῩE:F��	;�I��p2��;%WCL߹r(h3�y��)�v�| ��s ���c����;�`�ۢaz2�-��GTPۖY����(	�{���u �u$��sF��+Z��^�\��\ݛ��B�MЦz_������T쒵��ƴ��+���k��H�\�Y�'1�JE^)�	ԤԪ�r ���_.����y���e,>7-6 #s����fn�:5m�� t�2����l:^���وa�d�G��/�)�pA�C���Dd3i�B�_v�.�g���76e��C�i�那i*���۞��y<`�nTS�Y��j/��:���{gPC/)@>YΟ{=o�z�To2D��?�Bށ��!Đ
�ٲ���:w@͋��BS"�`�XkA�{�>�e�B�j#��%3Y�W��d�n��.�T�O1�k���BA���J�S��6W�W��g�l�UL��A `撸����1��(�I����%���ME�d[A�C�Ƹ��~/�2���P��8���Q4�W&�z{�)�e(8����@�K==
O?_B)�ͤ���1;�'F�0��Sw=`O �a��@%���-p��Yv�9�H#���x4kƆ���%�_,��������I��z��_�Pk���c�G6m��P�T�~Q��X1q�����!8�{�q�vwth�Tv�kj'�����
*}D"�!鰴!�(k�Av�'��J��&L�)6��׷n����/��(睎豲�+���H
F����p;K�9;�WbHc���s/z����w�)��ӻ�dHe�ļ�6��yj6�8"�z��2�TC��Ay�6�X�>�ȭq��3w[$�����#�9ƿ2��9qĀW*��V�䣶iᖖ��'��k�A���r����oҊ��I��pM���0�sR���/\e��v�X?��gb�'~l�����&�� Q>���/��(	��gb|N�]�;ף�a��5��H��R����=6�!��Y]�u^y�]����E�Q�'�9]�'�Yt�"�-i�ŞbB���O���*�|�V��)��NJݕ�Q��
U�pS��Ӱ�yh�����b��y��s SNм���Y0���f
}�3����7�-�ao��LL�c�{O��\�4�ҕS +��xVNlA+������M�� ��T�j��}::��v>�� �"'(��F�Q�f���U��u�	˵O�eF��!�����H�aL�ɖ�xʬ*�
j��nɦ��N?CBL��bu�e�;�D��a%5o�	m�ك띸����\�����4�1f�%и�.	��u��=���U�0,_#�~�y�����ʀpkA���������tI�Y��B`���aO64��t2���W��WXㆣ�@E�l[�ϭ@�����P��і�2S ;�>����癋�"6F�L�45ǚA�~��u�M�)���h:���{�9_��� �m<���%����^%���b����t ���@p/C3�9n�|V\�^7G	
��gl8p�:GU�0^`�[�%
2vͳl7����M`�-�qK�\�t����nE��&=��r>���C����؜�W:����.4��^�����oc"D�x@|������Z����G�����~�7�����r���ݔ�@����̢/�yRJ�=�A�8�ׇ�����"�HK�w��'�᧸p���Pj��A���ێ�_+�K_�G�ڹq��(KpW�F@�XK���J��ՈA8�{o	���Fvta���.�����5��/~׵ӫE(nEO��P����H31��B��ry�M��e���=��@P�GB��?W]��ct��"Vx��A�z��y'&7�9WC���VV,5�J1m%��9M&���+6��YL�z�CC�{ �a7�s̒bk~a�*��Q�-nؽ��~�я��Ӵ5"H��!�D\-�T��2֪(�qlL��nv$N���F�����Y�5buaR@����	e<�hZk�Lg�f\/<�����i��{ۻ������T�J��_��2"��BL��\��"�͡�Iq7��kTg�򳺍��Z�`<c�|��VƇl��E')_H�lX񞜾���O�����)���Z:���GR�乢�����aݪKڌBe�]�/�V�{����/�a�,��3�@ �Է{ޥ���#tuE��`u���7P�y�,r�:�#2�G>2��]qF���r��HNL'���&9Yn���xa��6�ǝ}!(-$��'�0{�N�Vg���WQ�c�*�O�
�T�룰_OF}��p�7"q��{�����?Ъ�Q�u?Iy�B�ȫ���R>JX|��d��՗�l���G���������YDC�×�N��gB��;!h�xE�1joJ;�1C�-QJ��G�t(���+Eq���r�a:~@}�q�e6�ؾ?T����g�"[��J(�)��j�A:�ВUZ�ϔ�Q7���XW�Z�W�G��~�#���A���+�L�=�,�N���9�+%y��g,d���ema<X���uz�����- �.�e^�%(ԫ��Έ ��a-DY2��`H�����<����r��%�u��K��ThZ�jB��Yǜ� C��tS��[��ct٨
�A�{���rA�'9�ækVbqIu�t���c%��8D�S
axU�}Y��"Ec!�6�G ���"��`��\e���kcO��}��I��MsD�Y$9V�>��H\镤;֑?�=D���M<��%��CK�.�Y����*T�*��gs[{H��#�
��F����PA���>��ܴ/�������� ���ZC�r�U��#OR�;wh�W�w/�O��K(��A(���n��@�
�4ۥw��D�cO����n�B?WC5����)`4����}R+��̸(�|�%�q紤)U�U�K&�"L}\w�_�䀻����yd�°j��8F�aDUl��=jcM�Ѽf��L֮~�	��V�'������̞)Ҳ�`3�3�R�"�����<V���/��3��+DL��[���r{����a	�z�b�5��b�L�<C�Ԡ�(l�"F�+��@���>�C&B�?	\DF?ӁB�*��a
&�u����HK|��8�}�	�$�l*#��M͎@�9���(��>ѕ��g���h����Cqys2"����`�t�FiY�꥕�3<�Z@��3E�N7�!����'�
�0��tC��|k��ë�L�|�w�����\��9��
u����q:�)X� ��.:��@��P>IU)�]+B��(�lY5��܋b���MT7��_K5$Lk�nM�Y�z�!2΃���4��]�]<�Y_VT��NV�������ꅾ���x�f�w"�Ď0�K����7��
�@F�����^9��!���e%6�w�ZI���`�r�oQ��8�Ѵ�%~�޷R��C�*�\[L�1��Ҭtg���������a�&~�~��:/j�8��#�Zi���cҫ�� ���>�jT�p�[�
H_����,�\X��l�xK�n�E�>	S��@Cr*���$�f���{u�L��c>^���%��*�CV���������ie+ϋ���V7W�Ճt�#xڽ�	���`D]�Tbs��f_�H�5�m
F�Y-�y,�XK��mvW/�yJ�� ;I���Дպ���2]����a�y��n�@��H2^�^Yy�.�㟞���Jݽ
9�c���AV1�	�= m��P�z�k�`�Ȑ"�!	6�V�ut	hY����XeR^��� N��[��!_hf7�(ƾd\���͡�H_�LqxF]5� ?�69�]-&��ْԥg����� �
 `����k"L�(�r���%[]0ꯘ�Z��Qyy}b�D{��~��ճ����ozgډk~�sS����f�CI%=��: p�|,켴"m����齃�V���xRh�ъ+��X�����W�q��� z�?B��l$a�^ΰ�����q��L�R`�Y<�a��r�0O�-��\E��:�m+�5�#[�"�9"t��菺 �ρČ��B�����l�)�(_>��%��MCv�4 ���<5O3�܈�VZ���k�����DփLгq�����L�h��ⴭ��ہ���E��(I�@��}��",`��]|W�J��9B��������&"W_�ȘZ�$�{�_x`إA3��
.�֏����B7�b5?����E	�I�*��,���*Y��P�\T����F���-9(R\j~��k�扈~�)x�VbaMl�$�o�e�scRV� 2�����z���u�.?�&�wW‍��0������
W���N�q]��B����ڠ6DXI��[�~�{3W7r��`Tс�܆l�`�E7�'/'����z�|'A}�l@�hh��J���8c����U�1���A8�]������  /dµ��k����	KP[bKc�)�_(4�2��S��$��ӻ���䉕�H�Ь�{�d�*���Q盱f�4�KZs�1X�'62��tt�8�^l��8h�`���:sG�.�xO\��}x-1l�9�2X*⃫.̉ka�w����D�}<�l�v=h�7�{ʇu啀���\D����7�5�����$A�(�*�g��P�)��S��p��~�'7��SO���F3푒^�M��o���K]�l�q����d]�U��쾼T��~2)`�+�Z�̽a�z�[o�nAn��t?�A�_00O��r�9p��y.bb}��crM�����������e�>;Q�U�I���RGIg5��D&\� �?vbX���Fv������Jp����M����Y �'444+����"z�|ϋlY��idk��ۭ�Ѽ0�� {F�X��h�rI �_�5�q�Nk0Et������Y�Ǫ���Y���`ؚ���3�Ӯ�Q�w�+c�k��Y�@�=��)yz�f�"����Ѯ'I�ݛ���R>,N�J~@4g)��n%�+�1T~ڬk�FbX7wX����;-fc8��+N��;
&F�m�~'%�wT���l�$��c��p6�{�ؕ��쌳���VR�b!=�	�yD�&O6�i�)�Me��}B�d>��ˍM�h�SO:B��i<�PZ�rPbP���5!�Ш�J�� Q8���i|�E*C�r�֮�(���!\����2A�[O/�S��u@����q j'����W�|�9� 0A� 1b���)N�������!�@�N�ރ=���f��E<�*�h��Q9�{�hC)�`��}���^����`�I|������=�*+%�M
n�t�N��j���,'���4�����#�x����=��>��"�����i��f
.dF�3[!�|`�O��v���#�O����S�0)Կ�7�d�y+,�O2��.m���v�Ga�uM֠f̄E�ht�n����p=�Ƅ�<})2��J�0�	��p�F7.�`��Y:s!��L�w	�<���e���6�b��&]����+,[��?JM���:� V9|bnO�H5��Q~���4��`N_U[㙖�1b[o73��OHCt��r�a$�K�E�.Uq��o�Cg8�yb�W���h~&��{{�Z86��\��dJY�s�X����E����+���.�]h��˷ ��YGʡ��8��g����L�]/���\�j�߄�i�����~[�֜=%jn�!i_3s5~5�V5���C��.���Fg�z9�d�ζ�鵙�IB�����X�N�qc�*H�F?HE<��gF�ŕ���H�E�0��gx���B�.A7���[i�zڦE�L�˚v>,�'�Ep��F
!�bv�O>��h�TFϝ����a�M�#�hX&o�<X�?�k���6��eN���n~1%�m�b�Ik�g��e&�� 7�)a�I�_�s�b3����e��/]|{J�A�9 �-��������0�}E�1��B��IC�=��[�C�I�
�ώݐ�g�:��u`�i���ocO�rƛ�Ĉ��w��!ݿC��1�Omt�Ҝ�5����i�:��
���y|���T%B�jT�)$�Ma@	y/��j�G4O�Y�?�R$�\�mQl,K�������A���<��`K���Dg��n�T�`��2�*���'������F�+��_���}�PL�F��>�sU�ô���嚪�O�xdt<�K��1��le[K�k�!1�
K��X�ĵ�1.�塩����_�Qܳ���~6�]�		8�˼���b�.u�W_������Vӓ��ھ�De:��~2Z�&�iL�� ;���[��!SmVϿ��z��+EZZe��,�����
��g�7V�'�Y*��b�c�x�r@l�d�qN51�D�i������v�{t�u癉U�YdJ~�L��Q��ۮ=�bT��n��B�+�9Uf�APu��Qx3Ah�ԓ��+���F/!�����>�O��P�ǳ1�)O��z�o��K���F����g)uM��*�_�q�*�{�����,&xX�[�b0�J���q\A���q�F��.�V' �]<_�*b�A@+ 1�_چ��C5+u��p��-����C�q^¦lSl�B0=�S�Bǆ�UM)���U���)dIb)�����v���nu��dg�З.�3�QGP��:�<K�M��o�J��'�����4�a��	0~� �* #��>��W��+
H͜���E���1�=R%���kٹ���\X���rH1Ū:���)}��Ȳ����wp��٫�����M��
��e:r
�uԛ���$x�GuU�$y �qq֢�ɀ�yi�^��I���̒h�:�ǫ_B�n��v�F��>���-'}�Җ��o�a�c��L�̰�JB��z��U�q���`i���߂�wV��t�9�8�ì('���+�i6@]��j%�Օ���m�&�>��a��n%�w� �P)��n �d��Xާ�b����W)��(T����\�I$�PZ��X>�们4_��9��x���}�R��_��dT��5�.*^��5_����FA.�q�!>�?�Zu'<�u)_>`�^óTtnl�	� �U������+�b�a��~��W�ڊ5�#u��l�c��5���b'�u�SD�C��~�ת�%2	n�э*��:k�p}؄w븶��X�l*9����~fxd���fs$�;�օ�)��_�yz�y1���S�:����J�U��p����F�
�	F����1� ��DA��x ���g��ر��34�(����K�T��Dmn����\�w���KҰ(��D�\���>E�5��q9��g5; 9�d1�H��u�o�����O���f>�/'�5K�ǣ-�(��D�s�d���a��XժgA$]�;��X�0�c�n!T���.O���w�ҋ���k��v��aq�M%i���t�O��P����I��o[�,�^�9U�;g3�`U��J����Jr��N}:�l�Փ���pmf�L�mo$���q�5�E޾��J�r�%ϪV��NS����}׎q���7hA�����ޛѻE_���i�}��AP}�����+�p�1�W}�7)G��ׯ��ѰC<	��q�`Ы|��Bюf�������*��#W/���	���k�gP��k��Y��0��q�]�.�/.���ǎ���Ko�Ѭ���
�����.��S[>�tةQ{I&o M/�V+�A��ڮ�����\���3F9��8��3�+A��ӡ¹����_a�ٟ���8��1Y��D�E��E	����!2g6_�$�|��᠍�Ҹ�����/�ͬz�����Y��M���.�96��fl���X���a�O?�9�C��d��DM��/e S��>�)zF^�P�S`x]���k��uN��G��%R��@rW�t^� @����W=�i�e�6��`���,t�M�\z�<<���h��ti�
(�1&E�Pe'(�����߫�`Q�kv��{����z��_Ur#r�U �%�ө�x:hV_��v�K��� �l���Q)\��hO`!�m�K����Zy����M�D�i�mf'~�v�@����x�^Z���"kdP�V5�f�����\g^g�<g�f991	$�O��wx��$�W�*������	�M-�+��a�YUc��M�T��}벹�,=hn�B� �9^G��F��;���S���[|��~���Nh�{%�g�G.hp�.�-
ׇ�=��Ἀ����ao�br�p�똫KV|ZфQ
�q��Þ$̩��u�Fd_u�XZz��LV��P�V�&-+�Z�ҾA��fsߚ��\���mJ�釰�6H�!'�	�Ӄbt��̏6��)i??���!����ȣ*�7���T�Q�����UML�J�8����BS/FH�k��˒q�?�ƿ���~x��� �/��Y��BR*S�y������.��A�*�c�v�mW�ܪQ LW�@{ɳ�ߔLz��x�Z�L�Q��vK�ؓω��-���1��5B�����
��''�C��� ���-%&��|)ƃ�u����4���d(X̒gKD�aߡ5�VӝCB��/�QX(\�s�kSNTZg�?�(� ΃��V.�H��T�rWQtl��R:��1tL�&o/������,�w�l�ɸ�vu�2��|�?���@��5� �ƖdDra �;/�F�N�Ӥ�1���\�-b1]�wr�!������2��oQ(Q,e=�]�b�D_��f*,C"]t���6^qfUL�F�� �\��aN�٩�k�W�Cg1-.�R��Pj �� {���w�޿�	���o�8s�G��c�w�b�ֵ�i��|������K�����FC�7��n#���$-oF
[��rq"��N\�"�6�,H8���_�.CV�$ie�e�f˻��u�'@R��7ɴM��O&x"�C�m�=���r�j�$|{ְB��?N1 �8��z�6J(;���:���՛��J�:�S�Шrhι���T�^ՒK��ca��5K,�F�G/�Q&NQ���k�hF���z18�H�����h0*,��g�NAP�^if��|�G�S�����소���
��p���$���.r���0���Y�H>&������+:Q	�����S�t���{L�o%`J`;RD\u.o�O���O�'ü*U������m?�xJ��cF��{� �g&���Cu;5�X�_g��:���+01��Z��������bhޭ-�I��)o���8�Ewu-��ݲ�GA��#�pF��i�5 W����mw@'��Bס��ih'����A� ��Ȧ�B<��Pv�D4)1�p� R�K~ӹ�����%g��=.�ѭ�r�!�	"�$��"tp
|Z���h1��p��}�(���<�Yw���F��AG�$��X�=}TN��{hE��n����	(�pcy�ʺO9�4��F�Z?���0�J^ǵ��>�[��,� .�I||��������]��+2|�qK�b�s	��Vj)�_ˇM1ۜ���fC|Ԃ�b]���.�=�ri����Q��x]�hM+]���1���-6#�.��KGVk��&�Ġ��<�c}
�,�m P��l�K�g؇BV�ΕM4c�kԾ_���H��\�"����\�6�/�:�mס S)�@�o�Fq��65��l#�R�+f,�C�3���)Hf>E�ю=�-�@�6C�������(��vJ��x/��2	���t�����*w�F�(JÁJ6
̥��̓΢��'&�j3����R��wi���
q�h]Rx�z9���x�� ���p��.VU�8%%��A�jB��٦��]�^���2�S�&/ob�$i亭�D����Vh����At�c���C,��g���������i���m�7�r����r�
��ܻ��
�y��߂j��,	;�I޻�E�pk\
n�0�d=Ɗ�]iNM
	X�ǋrfK.5R�#��I��`�r�t��w�+d���V{�K��А��c��~�/�f7v��$�/� �@�[��!�u�=/M>�L��a�A��dʯȥO��u��/ݙp]�7��Sv��6�6�1@�Z�Bs*�5ɈY�r3�#�+%��\.�~���Tqdpp�����Խ>!�����iT�j�}T+=�^��<tj<TX���%�M�F�h+�b��������d�[��NSpO@@����*0��Ո`#��5�wE%z��Ŷ)�[��%�n�����D��:��>Uʇsz
gf��:�O.�PV4�KE|�����o���bE2�ͧ�NF��{��F��n:�I%����a*v _:�J5?�}R j�;�x#n�,�{�D�d�ܠr��|��Z
�h �cP8�S�V��7t�G�x=�(5;����GjV������Wj�%]�/p�y��G�0�Xl`�<��R��w�,w�����6d��m&���/T�苝o�W|T?1�>'ȝ�e*����k+�T0}�>$b��m��i;"9K-��!t�#��<��JѦLGB�ӽ��x�޶�J���t�NP�a}�9]Yާ��α�R�m������iIKzp{����3ׇ��$��>�O�Ax�V]�I���R���L4'���˜�~t��v�$`�S����B���&]yl���9��_E�m%��}c6�h,^#���gt�J��N�l�z�V��"�^����_�twLՊ$�7���o�#x3��^"��h
�M�#9��L�孫䔮��.��R[��C �cUbj4E�u������;�
D�y�6�H���X���>�A
�h��(��h����������K��>�^�m�����o�}-��T6N6j�|���'p'��aOG����B��E3�D�v�II47Y�����[��|{�� s�[%��H�h�R)V��Rcp`��a��1^�q�gO����\j����|�M6~�\����ho�+�&��*��PWYz��6�p�M����&���'
��^�����`��4N>?RK[�b3dO��w'��YT�2��;Cڃͷb�D�G��yw�����07h�1�k2�2�0 �VY��<����aS0�Ml���6x-��c�e=�5+}E� ��]ۓ/p�/��>�,�6��F���8A�� Q����4��؂�ۅ�/hƱR�Q"��{�<e��au�����pcf{�}��Y�ؔ��U����<���q\���10�(Qn+ ��ä�^;�?K�����b��Ļ4��e��m�8����U�R���E[قk�;�������'����8�����8��f�p�\����S��_׷�2�3f\��� ��!Q�wB<���($���8U[nJh9���'7[__�3��Ɍ�"��'��k�1�ؿs�s��N�m��C�Q[�Y��s�Ngl����kC�f�|���MqQ�
�*��ϑ�p[���bm4sz�]J��=N_cfH:n��>$� ���{���d�{�3�FBt@y����W�4N8����M�zbN8�(���6�0�� �����)�v;�ҭ�W4a.ib=��#���5����d��8�QN�Y��G��+ K�n���V�(0���'�TY���q�
��%dy#jfwt�D}��8t���C\-�3>�o�$�j��8
��Dn#k�G�Ê����)F�B�LM��'GR;[ d/����g�F�J&�R��G;̪���S��>⦒$(X���-�Д�ǽ�Q��@�"�5֡`�:I�ك@���n��*$�]�N�˘_9�*���Lo�hB���09�s�|:��3;��q����t�$�s�<>,q�&�(,ݯ�G/.x�yF1^S�s�z]��Y<F��ڇS��+4�l�;���W;
��	�d.��� �'�ЀF+�bq?����x���NHp�R�D�3�Aϝg��$O�Y+�G��h��1=">2��]�����͝�X�G�߰V/�!�cۺ�/��ܛX�g��|�\������~^#����O<�,���%^P!�����z�b}�V��H9���щll�c�6�]DIkX 6��:9��f8�ߋ����}�.�"$|������χY�q�7e�g�?Cġ�$���6��fځ�U�Be���GX���� H�Y���������̼���h�}�@<�;�b�ф\������gAt.���ڻ�n���g9�$rF��$Ϗ��!����]Az�d�N���x��k��d��0}Y��g��jp���ͶN�13��(��a�\��TZ��-��6���W�	z�'�Q���3��-��1V�0�!��g5pk(w��z�l��0�����������B"8�/���ݨ&Y�I����p8u�9K,�S���#�j�Z��H�mU1p|�cV�w������=[�^��������:��������tCޢV�����[g����x���y���N�`u��������E}W�|h޲D�>cqc�:�)P�[LG�����_�5U���|TZ��q��w0s����͡��s�jw�[Ӣ|+�7�����՞�%|��^�����ԍ�>�bΐ��39Pr�e��`&ྀGm1�s�hZ>*�$���1{�r�,�A3�%�%p�f*�(h���)7Ig
]
����a�1����\i���g�N2s��DM�K:Ġ�ۿ�
���B��np,gs�7��e�\d}@�T*�!���ֈ��r-p�Ys�W�$j^�/��q��Xd��QQ�K�[h �si�J~��/�����q6���������;��=-Q$���7b��&�0Ж娃W&8�z6n4?��tL3n���ž��ȃ�ɕo
/ݰ`�	&��K���Uj�=M�$�7�3'� �L	�7��˥�*�3�b!B�tP��
6��g�z�y�d0�C�+�.����9�����դ��"ߚő�I/2>���Y���we�Z��Ӎ�0̐�)i�}�v���`�rʱӎe�%?EH�Z��À!we��G��/�؈�HL])	�)�a�q ��@5cS��&� a������h�te�[����3K�R�5it^ �_jH��)9��r�A�Z��i��Dڠ#J!������^.�	���v���h,-b�Ѭ���ڿ��B[����|t ����,1� )�4��u/��KX�N��9s;��p���,�(*h�H\;��E��>|6����@(d$[�ۧs�B�ٞs���gZ��|�Hn��`y�A?�>�9M_��ES7^C��ߑe���5Q��n\�U:���+��՚�/�~�;�  0�'2b@PK	����H��a�~b�M"[��J�/ ��r�%������&;|$�{��(qi�+ԏ��F�[���C���5�3V�4	SF�㑭������"�>��P��'�q}��7i\p���W6%��(7b����FƓxeg��W���c�ru���
�x��%�~�2v��5#,S���l��+�����n���i�8���_�G[B*'�GS��KU��:02�iBfv�e�?�O�J2���^��H��N�i�6������h�;l�g�LtY��Y�����]�%�3�Ʉ�qG˹Ii�(�]o����;�+�u�� U���H�M�?�Q��_�U�.���:�S�4���&��Q���!d�¾.vz�*A^�#Y[��H�j�ߩMp��1��e�BAMP����w�5��I�]\�OB��|���#q�O�p6'�~��"f}���$fuy�h������2
i�I(�Ӭ�7���2�
�|W?ԭ��G7A1��^�Sp�P�H��ǘ8X�V}Gu�5��`��\�E-AI����tC��'�i�@Q8�:t�+���	�ኲ�^N��î��0���+- �oY=x��x]����&��Ð$r�Ew˥ GA.Cč۬V��0B�j1�AV�O��d(�p~�������_R�ǌ�+�Jz(���.û�7���ޚ��aZ�����Pe�1vBO�r���[0��j��	��У��e���֮-�p�ɐ$}<��|�S���d���G��+-j��bq�� O���L��3�Bq�p�n��_��lOR��4F?��R�N��}�o��%<��`�S�ē�DKƋ��X^��n��M����ғ�+(EE��lu{ `}���G��a�!u�͂R%HȲ��~ �����Vl�˸Y[��1 ��NٴYfV�Z����(�j�e�=/!z�}��z�Fo�bI�@c�]~��m�kN�yj���<*��6`?f��	�\��|z����)���m\����⩞��s��t5U�}�v����,~1t!�3o۷321(�����8�mt���*U�Gw"��G�=_=�h7(�� <qyb<��q����<_p$%��'l�l�)��m��쐪)%Zy�[0��91X1?"S�����*S�!���+-��r8Rɪ��#rB��F$��!5�̰��E��,k�L6���t,1�R�Y�N�1z�$M!��p�� ���4���ijzrA��}D��?<��Gfs1��� �$�~*r��?M;���(���g��/��o�7�x�Z���v��7���/���t��ڡ:MҼ������I�&U�z��k̑GT'���ZL�g����6��Ĉ�Ӊ��`:#�ɦoH�K�cx��S������X���g ���:C��I���>OFR�|:��$$	ɁK�/�|��7{�{�K���:���{��x� �b7��KS�*�)oV�xm��úW):􆯚�7��i�Y��"��r'V0fDQj.�Ok�c��0q� -&?G>�\�0�����M���s�=f�M)��e��� 1�I�1#�щA����i3�T��83�N��x;S��ԅǔ<s�p&Q�$�ܙI����/`������e����vZ����Fec5��Dr�m3.��˸ܖ�в��<[��YR���jz>�_V9��a^U�̿�t��»'X�G?Ly	�M�4-s�_�+�$2lAW��)a��c7�Tyo�NHSv(6��B/�!�U�pe��� 	Gi�2GC\-^��XL�h������r�P�;.������G�+C}G裦�|]�ј�ky%KzBqk3w��io#��aJu��&�sP�.���Sl^�[����oު� )Hn�,} n��.L��k\����1ʨ�FVUsNK&M�&V0 ��9/Vm^���!y�],=A�Ͱ~ܧ4
۳��p�m1H}dk���N��s�]����]����O�k8�t?�-xVx�P�+�@kl�e&�32��Z��z� KV1:��L/;�i~�ܑ��nU�'.u0�Hi±�����`n��i"{dhpp(H�;���M�Z-� �۔�=hjFH�m턬�V;9/���E^o��?�����Hۢ>p�o��+�p�+�ߟYu<���@KGk�B���ɰ�@��zN^vϠ ���\�k�2i��Ʀ�Z �����ԍ�{�á��iz����ĩ��!�~@�gQ:�i�Pa��s�i)�\)c�1�ж�ޮ�M+�.+�a��T<K�z���V���.�A���'wE�f5�R�U=;FYI�'��s��-��u�\b�����exs��3ZH��_}�R5�I�&�푄;�C"u�NC�r�B����})��p%r�F�@K�۟˰�'qpO�m�3G%����^J�sM��ê�h��Z���������9;Q�vbL1�z>�%���%>�\���-@���V�F�Y�{p�9�8��%P�yM�N���%[3S�9m2չ��/�B$K���l�`$b^@8]e�G^�m���+�k����b��|���d:~��qtt���ga�mS�9M+��� �� ��}���v�l⹝���+�]�8x�F���Uq����b��<	�e�gK$�ל\؁����'�c��C����l�����������u�/���k�nas������$�fz!�6!Wx�y��5�>ӻ�Ep�Vo
�C(P�mm���ފQC����jBD$G�ĩ?��RFZ���˒)�|s�K}Pm�#g���4ts��Ѯ�tUkfA���O�]Cg�t�Qk��C̀��ϣfz4��t ��Iw�y��V=�}�)����>��M�T55�ԡK'� �f3�L�]#� ?"|K0�{���#���bv����jƩ�q�DQګ�:-B"�r|���&�TJ՛�_��Ԯ��rá��R����N���h4�®��]4�:|�Q'�+����A�by:a
��(2�jH>�o�3�-� �sҫL ]��)"X�7�x1<�ɉT���l��bn��4��b�����I;�m�۠ $��B�;��q�;���T\�t>v��"�gSí��� �A��zϡ�g�ld����x8��N��&9>��W0+%��S��(5IA#x߮K_�2d�.��JW�c��djt�p\f,Z���jfO<�@���8ď���������as	��Ќz6��V-~��\��<.@u"�����
Pz%���"c�ׇ..�!S�!�Ǌ�AO���2e)Xو��2{����ht���c7�yp�6���Y&�:T�2���2�M{~/��|Q�q���4��ow�Q��0Q�H�{�x@�P>���_7>�2�����	�d��)��k-`�H�_c�?��� �.3��f���X����|Z<��g>MRl� �t2X,�hK�)���x+�GU$�����zo@w�Б����m:�t���x�~ ��[`���X`b��߄�H$��}��r'��oRk1n���jAǷOʿ��Ų���拫*qUD��Tfޚ[�L��屋���I]�#�ѱw���؄ƹ���Ҽ]���+�7����st�~���f,�����l�V7oiBgPj�Ӭ�؉�5�ˈ���q�|Gֲ�>�{Q�����P�wŋRa�Γa?A��_��+T���mV��m3ǟ�a��\�:���?]"I�}& ��$�w����htW%֯k��C�&��n�׭\����Q��������TӮ����|��R�{d�#����f�jd!i��vfL=F$yQ�	>�I,�|�N�Y!Ch�� d�l���Uw�k���eb�~H$8�.K&�\�-9�A3�w�K�]'�R���l��,�v;��> yW���s�Ӿ mƘ	ІǞ<a9Y�(0HU�$�6� w~8�`N���m�#Zf�Oe�:�c��E�Ȥ�[����u ��u�OQ�`R#5<t3;Q�M*,�+/�%C�p���K��b>�,�޿ٌ:D��Ks�Z9��z��������P,_����F��̡����=YY]0��/=�!t�F|��h�G-������D�S<DG�L*���B`�#��$��oc�:���-�;�9ȗ�#BV���� J!�@�K\M�VX�#10��,�&�I�ﭫ!�t1�� YoЪU��։�X}]� ݊/��(K$yf�tB� ��M�%�{j����;1~83���Ӱ�qF~Jh��drG����`��Y�Z�v���X�K��p����A~7ofPP ��#T�ˁ0n�'�+��\(揲�w����&g��"�����w�]��b|����}�������6������
�Q�E�YT.��4;�T���O\�~Vh�
WO|^4��7u�-�NA�(Ai���)Eb�	�BW�k�7�����`���4C�bA�%��g��iHK9Y�S�q#^��Qv� �'h����B�A�J
5�j���-�qgp��f�U�wHiao�bM�_�S4�}��)G��^�@�{��i�tO�z��0�ZϠ�Rԕ�	���R}u�
Tu$���/�X̫8�s	�Op�m�~��*JF1��g�e�N�6�ڸ�b4�6�ۄ�\Ġ�����^���K�Q�2��oL�J���mX�����G�<!��)�-�L����E槴G��D�ޯ=k�@��X���#|p���0�ED�lڧ"���<�y��dZ��a*����JcI��ܥ3�UA���t��' �E�3�9�}4�mB�5����,��|�X&S5��, ��ǉ���y�4%��M�_6���^��<,�0�1u���'�K8�`.z�q:����ὰ�8��].Ώ~ۼu��.A��s�&�N�"��=�7R�9ێ���h�Բ��7��Õ�gC.|l,����%ā����5ß�K�Qt{�GJ}ж���������.�v�m<�S�
�~*���Sx3�Ұ#�d�
sim"���aA�i��Y
�n��;�ƵJ&fM��6J¿�@w�ɪ����p���
�0��!��P�����X �����]d�.�֧�N��5:�v�:���%�sB�m!=5����5�y�ԞTMٓJ	>���4S��N#!FNS�h@|��c��gP���$�~�躊}��޸'�bl����/�~a�������;�%N�6�����P���Mh&�����*��]�����z���VX�U](�ǣ!,�҆�K1-!���3�F0���e��釼��0�����ű�,�`ʂq���64�7�8��!v�?e�!n���|����p�}��j÷�EAw_(��^�RCB���Lu-E��8U��{�#�=�@�"N�X~��7�C��C����f�G�Y�%��;y�*z���&9p�p.1os��
�\ǅ�)<9��!�E?z���y;1��Ao�Cv�OY �.b�@�r���B�Ԋ�1�mUb5�dX���yKi�܃�Tn�ƚ����U��aO�n=���9�Z�v�08���i���:vye�0oZ��LpYu�D�(��֡�h0<�0OG�(^�F�t�N&��D�	���KsR�7�r>��	�[RB��(>+����m�M�l�y-H��D͎�N`h0�eo�����I-xg��j�5W��Gp=ʄ{s�B71�I�"�Jn6��&��0;�\Efݐb�D1>N�4=��=hgW�1)zn�� ߓdS��RdkUp��2�@�{�v��>�^K<M�'&�N�_��Vd�Va%6��lKY�,�� !�{K��}�ރ��
����V	�L���-�'�)����,��>=::(�i�bh�[J��Z3�(� �ڌ����m����S4F[Q�eЗ�N���񷖑�=� �7J�,�Wu��~}���?�T�����m���/z�.��6�yNl����(���礛f���ԳDGO�<pC۾>n�rA��)��жt֒l[��7vt7@���SY����0.n�=�|i����X��Y�$�RqL>��=�7�8&q�7fc�����Nd��ۋ%��^����m��w��P���z�6�o��fGϛ˿�^�E"�� �o���(���##ϊ�(����fZ���W�M����xY�EİIL�����Vo]���Z
|�����݇��U�x�c�a���I�������s/��L�Osb�yi�zT��b	��n��Յ���.��8ք��n��Q�vg�H}l)�5w.Q4�v9��A��sl���ѧ�#�?'��'���(R�����9펭�{��H÷�)CP����f�y��Cs�Q\(���^�<�B�P�<Uyeٶ�o?]cDVJ�KY 4�.�2�K��Wx΀S
�Y�Y�8��R����M�w-�(я+[>{�0K�<�E�e�,pj��)��#���1�2���R�"8��:!.M�q�� �����O^~��zO
j¹��'ҥ����.����*�T@�a�XJ�9����캥Um���H������];s���C��w)�2�floWD����i�W^���%�)�(����%bԡ|y�N!��R5P�T5�x��R�ɧ���~�PG�ה&�D�e��E�zy�Z#�u�(�}�o(�#fj��Q8a;"תz%����b�In��ѹѻ��� �w�����z^��[������LR�2+�	3�� wu��!�Y�RD#�̞�G��H��y�j�۝6�:��mo�Z3��P��\�6�ղĒ�K�Yę��d17�ob�,NQ��ԭ��Gb�g)������0bQ�dKY!�nZ/�Q��c�X�w����U�><�i�z�޲O|	���j�u�������'+e��ۮ�>\K��v�I�<��l���)Th�2�^W�����hyB�c/g�E������O��5�HR�YL*hG��OP���n1�bME�J �J$�=����{f�>��_�!Tq���]�:$�%�9~W�;�������~fq�!��+d�<������8�����Q�?���?a��\��P�6��ӻK��a�-�U����7A�f'X�X��z9BN�B�hj���:L��H����H���N��s�R��>
�/2����p������ׁ���ޏ�c����[�y$󧩴FRlq3�M��V������u��0b+vIY�-lDnr�ɕ-7_H�pg���NƗ�P��{k��:��/}hLM�"uIj-;����� �c�S�5lЯ�hD��Tgx�
I����l�6�et\#��Ue�h�xT�֠Z}��^w)ӷ3�g��������z�>�����Q)�udfc7���,�ez攨2�5��7���b��ٕC*�P��|�TU�M�U���ֈ��C27�	~��~��tFX6���7@���+zM���p@��%����j�vM?nŏ��<9�T�g�ߍI� U�TZ�{(�VSB��RǦ����G)�13�>���慮��
Ǔ5R���$ǊE��M�b�lsoq�E���i	wd�X�$��-E(��۞�A۫p�rl�?	�����sl7o6+��Gߓ/�����D�"�J|�U��d~�1�z�b��DZ����e2�z�+��m+L#ä6�ր(�]~	��u�A��)h�q$H@K3�,��F0�����Y��73�g��|�YV2[���l�Ko2]�>k��L{��9Ts�H�x]������M8"�V� �_rPoE_� �c�oݒ#�Z�v�����'GJG�lv�?dh�@����g�m�jW� �j���Q��=��li��Zj��
��Bv��Zp�J&G\>�����2�2c��<u���k�ү`��ʑ�,[����.�e;K-�X<r���Ou
U���u��6_7��4�1U�D5]�N9O�ѷ���ӊ*-��G��<��(��2}���%�1FD��~U��� ��'�p&c�89vON��H��n���o�2���B:�$+�ˀ*-h�z|�О��(Z�
]�G֐5�
E�������il/����aV􉩔�"��0A),+{�d!*j���q�#�͊�
)�X���	[��b��*ߞ3�t��iT��c��KrMUx���*����G�ܼX�
JW܏}_}=W��!��R�a��iU9�t0�x� d���ޟ�?������7Aw���������kP��ju5D'��q�b��En�f��]h\F�j��������{��y�)��aEb>9;����\!ߍԌ�&_cW|�û�E��w0fG����{���	KV=i�F���H19�_'�����f"9�.�Jo�Q�3j�P�SO���Z�Rti"�%� jK�80�X]�c�C�/ $E��.Y:�i;n��V_����k*y�@"~��*Ǉ�/@��"�%���c����%��`=��Dd͉|(�䉪��v�UYp��k����T6�-��v#�Z�Z���1�q�����1�]i��S,�ρ�=�*�F���lB���NT�Α۬��֯�1Ohs��85���-�6�8 ��A*l�9����6��-�;S�	��F0#�>��]��j��KV��H��X��5f�,��)�Xb\a���F�0`,�G��gͩ7G�}P ��$�
�� ����@�A�SV���/�H���5:�)Z�B�r�:�Ia/� YX:��7l��$zR��u�=3\�ד8��(M������~�i*y/���"�N��B��{�ŕ��U���2 ���ax:Y���_u�B]]&K���B�a�������̵ϩu���·a�̪�Z��yE $�*�7��ޜ���������D�^���c��2�{��Jk�.��~��3u�L/�D�f��{��*9D��w����V'u��'*[%��N�8���K�F(WAI���ab�hE70���5�U�A@��M��s
'�;������$�C�J�N�?AF�"<�#�9�H��'r��j��t��2ژ},��k��嚺o�t���mHb����
K���m���ݩGI�iAm��o[3J�t.�d�d7��;H���|�FUG-8�])"c/G���v<�n
��>3�kn�����iO��je6ǁO3�˩~���h;���1�Ȓ%x�ug6��"i�Z]>�̉��  i*_�C������,;[z��H���}�����&��:)��J�ǰXv�qp����(��b�=��(?.�l�f��!�qS���:$Xs�ڱ��XQG*[-�N����L�����Q�j����}��:�J�3�<��%q��d��1�؟?�#�R	��^ќ�!_���&�vR��a��M<XDs�
� ����"[h0��e�A2U�-�w�šs�X���a�>V����^��A�)�X�0vW7w:�E�S;d�A*,��:m��q4n㷽5���� �O({�:m��D�8���֝�M����(;Tw)<�V6m��
gl�1��~_�������s�Ȓ6�/�C�AZ=U��>
�P�ؐ&���n�3�(�#y��S,uMM�J��F���o��?�w6o��8f}��LG���+k�
�
,�0v�yE�"��qjB�	n�dq�w�獱�a��4'��Z?��DYƺ�(DG�r��	I�h_5u��)�⊫7l��+��h���^�f65��S�3��̭�x79��O��x,��e����LA4�@]�ɷE��au��oɜ|�sx0�lÅ����	��뤿4l�M{���A�.qPL�!�T����_S�]f�5�g/,0<�� ��!��&�	1l�I�� 8X]�U��� �y�3;zF�$�S�<6i��&V��h/�Y|\�T�A�թ�v�-�b�p���.$=��c(x�i`m��t�K1�",�� ��%h-{O	Z1_-$3�\	��6K�	�<<_K j�)���3ǵ���P���&nS� �=���˄���<�])��lr���q���f���r`^b����\�o��_C2��q���F�}�h:�%�*^��A���V�@Xg�8X�0m0�ѕךp���~��;��Pѕ_�:��lK�����0U<{�/��� ��M�^X����\탏8#�ގ���w��X��q�۷ 옞ܡ��''ѵ�f�ޘ|Q����lW8,�e	�`�
��d /B6]�#�J��m "2�:�CC-�$��ه��:�,�X�H�0}����86	�$A�������}CQ'�#6�f�h��:9��%gp��9/�4�_Ғ~}��=ϊ�|�����`[��Y%y����S��ka=|�lmX�f*��@�������[�
x��INy�]q�4�U+�����qrC��(f
ԅ���C�VJpWҡ�G�|<΍(� 5v1���H6S̿��]7���+�K/z0!@����J����&�4��i�r�f�ǳT˧@s,�;�(ۈf�8����Y� }�k�9Cc��6���vd�q�Ǧ/������a~]���`g:��ڌR]guɘ3�&����V; �����ҷm���'�-����� ��0�?	�Lh�ܕ�����xq���vy��J����7��%��ܾ��"}+z �<:�H���% O�~w�`�5`�6�rlH��D�%��駄� B��~���>0���_�����R�"���~��,	�&p�B��ګ�������8�iZ�C�j�,
k�9Kv8�S�*j2AO��E��s�t"lpIdP���<�� ��:8�C�M��j�g���PI�k�z��� i�p@�V���@�(���� ͚X)b��o��u#w��2a����*B�!Fq^��˦��
�_�I>f����ٖ�,��@܆�����W�hƵW��(�����}��!
T�
����ɞ�JbW}YU�S�5��7ҧ�,�:=�X&�-�����3����ys�0��}(��B�3n|�2�h��Qj�f�qT�&��Β�;����[��/S��?��Z"�"��p����O�:7���9t��jH�*���������ɫ:u�[hX}\�]g�`Sb����լΔ��Wb)���o.p�Hr�]�.�^I/�\�sM�$�2�4~G7$w��&�L-*2�a�<�%A���VY��_�٣��j(�/�q[���v�3_.�����0��Ɍ�"C��H��q���(�Šp�d����oCŜ(�NYk�^�Ht����d���a���Cdw3-�Hy2ʺ=O�;b�ZNJ�{�/�r.iI|�jSx��,f�B`�/.S�1��V���h�8!����y�ˡA1M��� 4��e��q�jp�-榸9R%0���|�E���j�C����~C�����`��Mdj�l� ��˱[OR��֫$#�#(�-~���ٽ�7I�#A��\�<$�=�2���A��M��כ*O�v�;$�?ƥ�3{-9_=!voj]`��P�pL	�_��t\�\=���tCt$ng�@{���7�hiw�RܼA D$m1��Ol�v���M�}������]7@�&�q��(����_�d�f����2�V�A}8��,�����"P����/��������ǗO�y;�K^>
^��k�x��Dt���X�	�Z���T�0$�]� \ ��Ǝ�6Q%�=�և�U�E(��s�
TΛ{#�!V7���
����958���]p�d�y�@����9���Y�%���<���].,KX��Ǝ��-aN �"�_l��i�E�>w1�O^Ր �d�-��E��cS<S=�,4f:v'��f��X<}o����n��HA�P{��jubIUS�;k���^X�3��4���L���}��E�4�l��h�7*�D����x-�܊����xT%:�v���Ǝ=j�l.ۅ�p��'Zu�����_i��D�"h.Y�Z'��h0��_1� �Sa�����oa��Kmmv���5J{!�z2	P��E�Ce��:6�3�ҴC�Sہp�@���%��T5��$*�խ�$��ȴ�%�N���{V�:�����O��j>g���^�Nm�V�$�B���؃;��e����ej@��C�ة�2�����ϥrJɓX2�y�q��]��&���ewr���T�M;��L�􀰸ίڗ�kP<��p���J��җw_�w�y
%�EI��Y¸�m	���'�ۭ���S�Et�]���"�m1�ן�jf�M�ۂK��3�҅���(cǡ:��,�n���\h��I�T��ǅ+(���';�0Ix_��%�ha��s�S�R�*�F�`/F��\��/�U�W��*��8-9zmݍ�7��t4Y��yJl?,�yk��o3H8N=>��PHF?�M�/*��Ⱦk�o�(읊М����^	�r+(�z�K�ݢ�m66[&�bSd��[�N���Z��Fn8�ح-����s}Ai;~ߟ{<�bʊ�l=
Y"��1�`n�(���+�mS�~kw�q���˺�e�x����.��A� ~�&W�����'�Y�=�>�=�����p���<��&�G�S¸�kC�����V�&��i��$s6RCmzޓ���x��@��E.w�s�r���B��Uw�b��A�Y����s�IK�b�%�����c�{����8���u_���٠�eJI���'Ǽ}!�˅��#jbڈ��,r�&�x�Yl�t'O4S�N��V���k��,��h7�SCح-4�8�[�5������%E7A?u�l�Ϩ�G�kU�6��4[&{�2{M�?�ؓ�9�� ��E\���3l�T�t������׷6�T@1��}�rܾ#D�Fj^[I������ܺ�Ɏ+�FZ���q؆�>���a�B�.��AxY5��zڂzY����"��^�=Nh`������vw�a{��H��{5Q��W��9�%�^���R�
7%�ЉT�-�ݓk� v\\<���K�]�V�4O�pcĊ	�"�0�i���g��<��0&ʈ�)� �� ,��I��kG/#������9=�e�(���KU7ʻ�p�5��g���9jw�, ��9j@���n>Q���(6w�
�J��$� Z�������8�j�oTjj=6�g�}k�Q���e	�����׀�̄��n^���Qhm]yf3�fb1�),���z4�PɍBu�j##��q��j9�.`�|��k�l�[�'�۹���#|�V�������s�XPgeL.��a¸��=ͱW��O��>eш_(/t�CX�w��yܳ�L�!ۄ��R~�j�@QT�ȯ(���5��gh�E�od�!���3h���aiҡ+~aă?�J��n�����Au6����� ��������*���d���.��\�*�rE�8z^=�
�´��df��h
s{�{�9N�n�
�/|��ba99�b\Q���y�C2�9Xl�  ��y	6��;���Nn (6$�z�K2���6���,��Q%M�;t�n���gr⬳���i�.���&���K�\2�XQ��p�V�$m�.�,<+��%�4h���9���R�΁�"Z��_��2aP�zP������ٌ���-�A�[����+���	�k�.��y=z�Ŵ>bPP�τ�\�t�������h1����:�tO��2��Ҟ�����}�39G0���j ��)͔wTɁ�q��h�h���񃟠Y�,~�gd6ɖ��eF��D�'j�-��r^?[�pT��f���A�-�AK�"��A���4������θs�t�]�$p,`ŔZ �X���!E��ܺ-.H���"�S
��g��(l�i_����v��	H��ݱh�RG�ȥچ�p���rЗ��N.��8:~��<!��]h7u�Ø��˖��76���7���x��5W�Fw�����s|S� ���bߒq�T%�O���ך&?*o��k��C�N9�5��\�\�b�/P�s�3���?�Y�a瑁v������;����~1�;�MG'^�� � jp ˵v�8۫���A�����m�d��k�4"�=��1�g�Ʒ6�_���y�$���X�8�·�L�hL��V�;K{�>dZL� 
�4M�о��s$�@F���Z�"""�l��Ti\p�~����O�	Y�>>�`� �<�Zױ<���(��'bB�'����������[W���*����a�١���B�<�Ƴ0d؟X����K�6��$As4V�}��G�D�a˿�|���k�
b6j�[=���As���ײ^O*WI�`h �Y��X�FsĦJX�T���x���9a�+F&H���v�=�d���)�u[�*� �qA<n�(o���=���Au]6h�h���/0����HZ��dV����w��a�����"q����
��~��L��}=�[V�FF }6x�-S$%^_O��ښ?���IV�Q1�v�09�u!��x��>�CvWJ[Tdr�*[�}}��o�9e����{���M�5�����D�D,C�7��Q�5��G�6yte:����­�Js��\���mS=Y��wc��5��?~�/ɋOߓX�4L�~P0`�I|��t7���37�n�)P��zԞ	��h�����Y0)s˙��]���G랰�$���TYo���uTa���>[U�*�j���m)	��hj-E�()ujޗ	)�XX�uQ/���?��72l���2\�za��,���t�S�n�/y&�e��ԜL[��)B�1�L��� @#���S��m���rXP����G,7t%��kR0ͭ�$@�T@ \�U�8�me3q�I[��~dUi¶��E��R�+��������Y���[�or����{���"���i����*�U���7_{�U>�A��ҙt����C�Wn��x!��>6GΧ�ߝdG)��̩�l�}f|I��2�p�y<�5�Z���.Lq��b��	���#��E� (Wي�t-A����ex� l{�4�Np,�Nz8ߟE�g�"o���L��{�X����`�p��U�d�q�)�/���ܿ�ԏ���l��R?� ����B��r{S@́�ə>�t��{a��8M�L1��$�\�х�8�c�at��e�� ��mZ�ݕ�����ݾ���D��.h!�/$��#y&ʿ����Ԅ=V<��i��R��W�c/
�H-W�#�8�����s~]�z~���`;ø��[� 닩�rb�/��" 5�S[@jm,���5���`u.��x���&`u-tY�n���ǳ���ηg����Bt�"�m	u3�PΜ�Qf�%�]%�:,d�nBRw�vj�g�Cn��=ͯ����:�g��*%2eb�߿���}��
6�;Ӭ�uȻ�b����=��DP������a\ξs]����X�G3�wAe)~J�lt71���l�uab�V�������84h`��L�.�w������~_5��ő�Q��ݢ&i}�L4{�P����"���I�-#�k}��4�ț�������e����z��)�p�qs	{�J7�1����5��9���_�Y�?ԛ��!���J��k4�3^Y�T@�vCu/[�N��U�_�`џl�س���0E�����&~o#��C�Û�3[�]�#��d�(�:�H�k�w�v��>�tgLM�n�C��v���rښ�3o�^��ɍvS�����=Y�����᫄�Ď��4�7Eq��e��b8�o+-�b,>97�+Ю7�sY@��f�m����u�T/�V��d������BjSz(v ;1�3ّ6�0�v�D���_��4����S-�T�w��6#�<HŞGE>M�������W�Iq"x����r(���	�<���q�����D cvR�h>3o,��q9�����%��MY{qv'|[[�'���_��� ��|`o�>ъf��}^�z��/�֒���>*y�V�%/[J�1ޣ?dT��1���:TA�jP��t��j��gKL�di&s,�v�bXƚ,�L²a�As]h�b���䇍�����m[sb<����yd�����L��܏���KX¢���l|��'�������,*� �2KT���[l����x�ݿ�N\�n�+V�X����5�a%���֎���_����É͡���RVm�Wpv]�D�wm�~s�VYSy��zߧ��aþB�_�2��Q��q����r�;�M�t|)`9�f��Z��K�ؖB���)ڨ�.P�9�xTLj���m��؅@pRװ�R�( ��&�x`�d���	�.�>g`N���q6��Ϳ��Y^ѱӽW���n�z����]�D�|��K��kۙ��5����`(�����`�<����'��^��O���/
�9�1��Mŷ,��D��tW9�$��P��¤�>r.�D �M6� �/>����f��b��vp8/�Z������+��n�h��!U��^O��� �̱u����;Ud�4霗�4P�G�>v1ٙ�K?�*�:�������QB�R������0j�ե�<æ�k!�p?��C�rQ�Lf� /{���+�s"5]�rѱ�����tpS9�J<����A��#�ەZفc�\��d��{���+0��9Kd�Q���62�r�w0���zk@]q�R��#���]+l�a�C4�R1�@��H���7��8�/�W�>�W������(���:�zvþ#�!�OAH1
�����Pj�� C��lJ}a��A�U�\�в[��dּG����ḱb��|f��ȸ���~cE�\�]X�3�x�G�kpi(�� ����Y���B}p[̒����Aw�y�/"�$`�ߢ0P���N
�����A���?3�b*�C��5�+El�����?�R��84z�A@�Y(����O��������K ������C�{c`,����-��ޮ�(���;(i<�g�<��>��+��ujmBE��{;�mQ|��{\F������Ds#?V[��(Ք*���E&�=�^��}�9Q����DVO'u���u���@<���N,x�*FS-����`��k� �u�(O�	�A�&�l��E�t����>�d�	D�ED_4���޲��]@��d�3_�Ԁ&�!�#^�h������`Rd�CIy$)�r�S����+�k=�I�p��^=Թ��f�GP.�դ�	!��0��x~�J�Ծ�V����4@�<�a�;��<d♓h�Em��iC��i����̙0P�J��?p�b�	��4zz��ư���K��-�)㮅�"-ǰw]� ;�11��;q�����f����^_=����_7���@W�����^NS��;	z��������%�Q�ęX1��ѷ}�[BYJ�)�
��c��U���C���7�m1�Q����~ǜe#A�f�lk�
+��M�̈E�gY8���Wٳ�~�/��S����Z�G&�V{ٸ���_���8Vկ�	�¬�U��pu���xL|���%i��$�w�]��Ѡ�>~�mu�r.#Κg��l�fڛ��ǚ)�|���!m7���XEBM.�͕~Щ��}w
ؤ�*>@�o:B����\�(��|�^P�{�/�w���=�'�����9��C}
Y��ٰ�x��t�_�N�o�n�B�D@��
,rd}���OO1��o�U�Y��3�7��Rc/D�� ��;�6��̉8E��,ߖ)��@�Ր��*xg	��a�rL�"l�rп �0�О������h֨��O��*�N]��y>�_�ʚX�����;c�������2Ȫq���%����Θ�.�8�0=�v���5n�4�g:~ *gd�sc�Q�<Uk�:!�ty���"�1n�� ʞD��� ��/bǁ"�$�&�-�M�ty�i���m}i[�4���x��A��w]g� �|c
���5O��YI ��n�u�^=�K&���s=����A�T�%�X/?��#��u�v����Kq)��k�CPγ���42;�F�@��6A��B9�B� V�H�����8f�P�a��ӵ���6r�s6�Ff��YhԪ�*�0�B~#z��N�F2�^#�~������E�����pg��mR��@I��W֋�0�"O\�t�Q�ۜ+vyƧX�c�*/��W�J�s��a7��P�����p�~I�]b��.��_i�W��d�%�C*�A���>Օ;��+Ts��ޅ�ҕXF2�нP���Ӣצ4ֳ<
��Ly}�ǗRd,��]�����a�C����g*vE�oީ�t�	\[��� ��*@�a���PJ��ćW�UWG�&k��B�C�mpCGIJxՉ|y�L�|��2r��VV�S�c00[`����D��H���d�j��ơ�=��C"$�1�y{�w����^��յ����&�Xl4����0{� �sɷ����K���Rl�e�3���9[�{춄��(��2ʾ�J��Z�x���<7���ɢ����!m���˗�҇�_!��Bl���Bݓk���贜�]���O��/װ0�0Q(}o��P\�Ϊ������y��
������� n������͝i��{F���ǆV�s�%Ui
�y�yq��N���E���s��$��gb]�+<%7b��A���zszp�yo��E�,Ա��d�EL�մ�I���e���m�o*�(<s�!��QɋEFQ���2{M^����-_��9��?�q��P�A~]X�96��n�!iCTo(����⿴���<�pfT�oy7D�@[��ڝ�_��q$�/�Ȥ���?�UȦ�8H�h맜������*�e-�d��:Y��$���&L�5�%;؂�{��h��_:�y._k��t�y��
0yҔ�REΜ�vr7�z���%���Q�������Ӭe3A{�Ke9r�o�x�[?��>�lre�(�ӌh�_�#���q0h_U ��"��\�ε-)��p O����]�LJ]M�Pl%>�|/6��ʯ�@�s4QW�ܙ�d�oq��]�S�W��;?����.�b����,�$�1������ G��UD�Q����s?ᨧ�q�wͪ!��Rj,`�5�_��n�τF==���B�c��?��Y�=!%��gĠ�\}����:�U��*L@6��/��'�� �18-��ϸ+ݓ��2X����1�^��������#Q�Rc��\�8fY�V�3m)jԹӳ*�Br4D��m0�hC�̨IK"�A��d�����{�F9o��]�!�&�������ġ4�@�Бx�����q=<PҢ���ڗ5���\|n�:�;��h*:���RD������bL�%�t#����)]D�o^i��wL��/�Q��oNuZP�*B�r�����4��Vb���Mcw��(����ֿ�	���
s�V�<�BK!HwW��.8\;l��i7���,���e�K1�"��l��#W=|[�����Iq���V�޲m���4 �E�5�������U��{%�G�����ST*G�1�b�T-��I��K|�[�I7�9���18N���w�`f���ra�D�߿�4�fL����JD���Q��Q;�!�|����`M�n���L�"A)��֐�nR�KQ�1U�:X�Q�E��讟m����4�g��ġ��t9x�����v3?3���_�\�)�	��o�-��������I,��uZzt|Cx�F��<ޟ�c@UOzs7Eb]Zc���w�E��$2�o�*��\?_'&��v쏖 �n�S������A3qT 5����uD`��z�Y*���1PL�r��P�jM��^Ο��^�92�dSw��Sk��+,*B�"/�1E��{�2���`�o#��g�0"����i��7���OYx8���6 ���J�Q����7md�Ne�X½;�E�\��HûV����GV5Q�:�&��ņ�ͻ���� �-/_6���:�7�����B���0�[ϭ��Z�dpP�0�����C�/��9R�u��L@��y�����d�w���A�1� ��>�b޿�g �/�	�y�X���(WqHf�U�i��4,�C��m�Z�����V��������nΥ}�H�Kܦ��L��p�W!ȆM|/߬وI��>���s��C�+3��U�0Pn}���"96��T!�!�����O���й������wT�Q��f�F�'�a�z�S�
/���r��6�ɖ2
INé��#�u:��y_�$��Ǵ��\����Hrc�K5�S�?�S���{��bm#�����6�.��/׏�����?k�/�B��No�x��}n���[j�G�)�T�k������x��Y*V��>d���m�������(��V��A���%����n�#V�^o`iJd�LO����&�4yI,���ՙ�j��߅>�lɈS+��F��X��]�h�t�ґP2;�����"����6���y�6U�|��������5���g@}B��]
���h���.���ZuG�?4�c�E(VC�FB���9���#+��Ж(й��Ɖ<f<lM�s+eR⢠�p��<�j��Ӄ��k���c'S�Ϭ֩���Բ�%2��"�B8'���y��~` "Ic��[�h������;2����� �Ǩ��ҝ�?��g��墳ڑ5����qCF=L�X:��IIW#���G8n���j������I� i�R��#,+�쟨�~��D�~ �.VЋr��<�^l����4d��E	�Q��8����czg7��r#�W���A�SЗ_�8a</�jMҾ*�W]�1�9U�C3���o�nh�eڪg��H�т�;Fx$��k[�Cƈ8��Es9p*eϏ[����DP%SDǋJ�&��qLhW]�W�@
����v��:�m">�B<��tl'"%�F��n���G�Y];�X0f6�v�:���\�A���t���Lԓ0>Kt� ��JՖ3��Y�ᰀ�(k�w�-/as:��#��8(�Q���~�q���e��d���|)o�6	w�N�4W�[�ƁVM�L��x-@����xD�
�Kb��0M���TquQM����F���c���'���v�a��]���e*�ʐ���p&s���O�S=.�ˤ+��[q�Uv5�Ĉ�5�<��X� ���������EH`�)�眷A���ځ�^�Z(�`ﾐ�/�CU�b�T��'9�`�2�x "2~��)�7�
�� K����zh��d}�d�M՗�8�g�t�./�Ú+���bf6Xy���1�z�]�'s�O�a���8fxu?"Q�-�/i���&H6cʎV�Tf���Ob&CK��+���Xi�.�9�pT���O��	@1���_�ͷ�Oh"J���B�����kR3Q��x*PCCa�3�s��j-fY �J�GdyEn�p�W����q�O2��_pt� 5ٌ='Hj�p�uׂZ�~H4Q6��a��0�dLД:�6q�hLo�nҧ�<��8q�$���&l��4])��K�jT�Q��Q	�z9��.�}���0`�$1�eE��c�+��DPa#��f���NA	L�&~�I	�NV�����s�z�������"3"H���F���w-QaXY@�@��w���Tj��SJ�!�����C͛ �CW�s2&T�v3�Ş��������/�a�P�~��5A]	O|��ц������<r.ڙU0��D�J7�ۄ�u�
�	�� ����T���dw7�'���1�zQ`!�7��a�	��e��K�����G2�x��^E�oX�
�Hj���Tٸ�A���2Y���M{)<�@j�n�l����	F���A����h�.�����:t$#b�zay�P�h�*���)`�`�߆�D
5)��^�Il�.�-{ş~7����j���\�)z#}V�\�8ܿ���Oe��z㈌��!��̩Ï�TLL��B�\a�����=���z+�g�色C���k�t�=��oz w�4����X����W��§4�U,3lL���w��2T�v��O'e��a����E�Qǁ��U��CE8�`��s����J����*���)'Ν ��$+"��5�J�f�s7u`Otf�����(�r��A�|Es���i�T[Ϩgz.5Fv�O^Y��O�����WV6�b?h�Ag��b����|~�%�����'��p�����(t����o�`�c��� ������է_k5$mGB�2���K+H��$�n�$�
k�؂��y"�o!�6c-�b��Ckg�D���������%����j�O������+nKO��A���ٺ�������H�*4������rk��,}�r!����\���g!�]J��j�"����*8ŝx���1�vɝ1?�u��H�kk�iL�8�D5�g5З^��bdt,z���=nx��h���� pEb�����{`
dP|��+U��po��^<ȁ��8��-DW��mi]�u]a4�����^�/�*�D�>�֖ʎ9}ˇcB��Υt�j��*/Y���`;��d� �w�&LK��x:����=(��V����2�
�L�1x6�""!��񥙎A�ݿ� T���q[���!zo���B�?�E-
��Y�Dig�u� �'6��w351j��	4x$�r�s�B�r�6cw垭����x�7ud�K�꿻M��sj2���D�p_ء�n_��)O�e��H�X�`&��\<���t��*��;ը�r[Q��2xm�	J�[Ğ1�5@�3�b���2A|tC���$Y� 0�bxS$��x��z��/S�F�� 1�5�My(�d[��?�sBd]Ş���ǰ�TL�]��]��t�l��;e������ǃ3;|v�������ݗÊ�AXJ
���{�{���j�{�ۣw��ԩ�0~��if��c3'&����^|>�����9�za�^'��t��Z�90Dp'2�i$�y�@썸�E�@>Ϻ��� �6o�A�Uz9��LQ=<�U@DC��ˏ�'��Qe滹t#������U�����	,m�u�N&�ge$��Wt~�����x2��O7�(zD5���c~"���ɐ/�A������%=�Fk����:]n$i�:���Vc ����|��Mnޖ�(0D��2�-\�1��1C^U�a�=�E�TR�ӠJ��CR�s��1�J-����j��<ߓz�X{�6�-�e���&��z*�YnLw&Ϩ��C\������-f�*�x�Sp��,҂x����f ��3?cA?�!o�r��9�n�{�/���J,5s}�*�ts��L@����j�������܍��5��Lf6ߔ�8�5�Rt?=��$0* O��:P0~��,��́*����ZNL���!,?��N�B n�v�l0J�O�]s{�m+"��Q,�B����g�t �����r����� �e&fT*���4�cJM�^!��_�7��I�]DŠ&<���#j�m�DLe����>����z0}�se9]sǤJ�?+�3�X%%�"j!�R1���A�?A^��X��H,g(P�M~HzЧ���¢2a �? ��p�и[���z���՞��#[���Q�oE����NA)m�r"�F� :~k^���K[)��3���T��W9Tln�|� ��wU��`9��Ӡ���UѶ\Fp�������W��)2��U����Z��7Z?�m��*<#Du�Dߊ�a�
x+>���Ǚ���`-1�T��r�yg��ʳ�V��C}D�(,k�̈́G�~�Rs�PE���m&���4@5�PTw͔|b�Gi?>�HMYnh@oe{'��I%�+��U>_T���3R�<�\R�����t���(�Vx.��x�$�e��&�л���`0�]�Ua�v����H�|���C}�ǧ{@.ƫ*�o�����xKU��T�Jp��É"G(_�vɏ���UDi
��(��Tm\,~'A�ںr��A��QJ��I����T�+ �	I�Pq�:���?h/V[�&0��F�`-q�P�yu����������a�)�z����0�A�u�F0e#�L� �E��P�œ������ÿ�YX�2nQ��Sj���7B|�Z>��P��J�I
�� N��K�^p��Tul�L�qe3�ɵ��Eܿ`�=퐇h�s�S�d���{1�>�@���º���|4�\�=z|�s�r\��:��-�I��
�����N��6��G�Vb�=��1��'����'2���R�OR�b]���>c�U��H�z�h�0�wn��ur��[]��5k�6)
��������av��v��9�
��t,������=֊�?�;q�8S��I�o�$��c��=u ��_�Q�M�;��� ��9kP
�����zJ��;�-Z��Pq���$]ӥ��<[1�N%�|%��I?l�����Z��o�(�r�W
�=��V9�՗�-�B[d�*�<r��';����	fၤ�Jqc��5������G����A(��HM�������8�nJ��l
G�94�W�;	��nD����L|�L��^0����.7��\��B��n~b���
Cp�m	w� �vZ�/4��S�5��o�&�c5�f:� e.���ݞk!fA�(�x`��54'�FP���69��R"�7b����B����=,K�8ZEx�8� ���?lʗ�=�ٜ2���M��ī������P�9ʒ��Ι3A2�b�� �g#/Y�O��9�EK�Xo9P�J���N�xؽ�ιo4�B���r�6>��m�����n��e�gI��_�Q�M����C� =[J@�'c�Q��d[�WȀ�.�i.�\�lG����*"N%>�m����3�'���3֤xf��G/�[�J���|Q�@�����3���t�8�ˤ�0�i��ť�D[��������=f|����`�B�E��t?�iq�`�S��3m�[��&Ħl�D��^T0sH��ΛE�t�$y[-;��]HuUv�˺I��6HNB_��^]S�r���kc��7�7�����N<�����zu��T�v 0}#u�Jw��D748YS@�aS���85z�΂D����e�ӆ'��~��y���X��)J��ܶY0|` S�%%b
[��K�Ut�TI�e� �G'I���ik �tJջ"ޝe��~��D�c��#����6�8$̩�sr��k{սj�T�dp�F��ظgN� ������f�@���n��/0�T1���
�TTGc뻷Nij�[��FͼM}�Rƅ��rdڸ�#��j�<J�((�2(�(�R�8��q,/c��Sޱ�/�jd�VG��a���v��t�sϏ�<�D.��][���g�w]ޱ��5)M�h9�h��4Sq��^
��}�/�{�����Ik*���\���P�ېC�L��0��YoTTÏ/���9YԘ�@�fw�|�4��[�K��*��fF��ln�9���,?��2��k\�_�����)���HTS��0J�wk�Q�R2"�;����5�-V� ��BNg���˺�~e#l;�n� %�Ȩ0�0������[��
U�$x��>M�V$�p��fBG���F\�n��y��w}����5��ӆ�����z{�Q�Q��/m�	o)���D=�f٠[k0�-s�k�F|���T2��Ȅ��gE5�	��ِ�6�F��Z���-siJJ�|����~%	l��;�2�ԴY݇~�Zz~�v=���<�\k�!�&���rA���I"�~Fs~Z�v��M+�_�@R[[�bu��YL$]4�x���u8�E�Cc�Y�g.@=�C�ºO'�\��v��J���o>>��'�`-���;�2>BY��ާd��\Zk-�S=ƟI�|�� �B%ف�ҍC䒗,$���9�nY"�\��.���X
��".���z��$+k�h��O�c*$@��2I���P<���R.�����(��3J�["�eU�*X�h;��D�[�����-k%�k�abː�TMHDx[^$V\�[:>��{_&v�&&_��>2Q��)̳rr�4fs�A�Tj���5X��K���L�4������7�m�^��(�˫��3�LȨ���u:x����䛀k�½ǬIz��B^W��y̤�U��ֱp�DдEBnV؇A{�l+L>����2��������&㛵�r�|�bF�^���O�;e�-_D��i ��,9k֩�f�$U}\r��0���3�$0�%��[[�\/ar����0����)'jJsӃ�J�r�}��VĲ5'�}}a%�1�y�7�V&�:~a����̹G��Q?�W�V'����x��,��Q���~�C�[J&|��Lò����O�)�Yd,m����0��i��1f�K<�t���T��J�FL�2�J��\��m�*�)=y�π}x��'
'p��$�	�����4��<�Z��J@_@��h�'?j�$��t�-*��Q�{p����/Ƥ��^�����������<��E�2V=�FMC	t�w+�����#��I_�����N&3פG�M�G��y����϶����r+Ro��d^}�%?����j(���Tn�Wk�f'�=�]"5���Lؼ]�/-��a�S�B �4H�9)�LS���!@���|P��4c�>�}�������?	����z�׆�K��a���1N-�W��wu#N��.�nm1a��ҡ/����`�hD�1���ӥX��W�'�&�j����+ ������f��,<�n�4]쐩@��ӨE�}L�#�����gD���vk������G��l�r$�_D��R��i>�ƫ����0,�c��l:vz4��ѷ5�.u�Q��/>`���8	/T��U��B����=_<w-m�=���t!�	�5s��`4���:�P��&�X�#�Ix���mZ+�P�?96��\س*Q�1T�˷����H��{/���P��o׎��z
:G���7qKl��$o�P�B�(8�p�^X��}�t�=KŚw���6��v��c�U��������!�݋H���Ռv�U ��r:�SV`����m_�*�A�I�
�����r����9w��A��`��+{n�y���"�<$�{�y�xh!��`�YX���Z�?��:�y��x6������Z=ϳB��/BoM���߭�_�t�������v�~�k�V����E91(�{�<���Q
�ݶ8H�k���ʍ(|�Q	���z'��cH���7a�ړ55Ҏ�<ȝ�[`��Q�� a���21��5"]��Xv7P�y[HI��j�@V ���^���� /NK��!�dw��v Mɕ�D���U'.ܝ�O�7�	�A6�˚:~�U�oLȝ���E�uGN�OF�"�n���u|�z��_���Y��(�l�.���U=�\}�.��"�D��O�{�y�nf�w�YV]�o	���@��:���g�����;�)� ������֒Q������x5!MX>��6�������l��S�(ϟ�B{?o��h��	s�C섀�0���رAߒ�7�>\��ji���Mքw�n��o��,[�Pt��|������@GJ��V{jo��k�i�p�,���(��!�8K�s���%����GF����(wh��v-� !�����*���\�PW�ť�?(���'�J�U��'��{�� �暵/����D����͓ߎ $xl=��2���C�H������ .����������e�f���BS�f��y�I|�C��u���S�$���O`�Q�Qb�#ћ@;����-�G�#U��߾�U��V���Sڴ/���4����.����-����ĭ����Z�R�j�w�,a��9���Aw1 I�۹s�_�Ɉ�_�q�2N��2��炂��	��[D�����&����2��l��O��B��n��t���R�V~��G�Y(�ɖ�����P����,ҭ%/~���cH���%g�IF��:y�Z6����S��s��k}�_#}{c>���R��I��<�D�D��1dч�m�C��R�:�b.3'~N�� ��ّ��?��h��,q5��ҳ`��&){�� �jn& w���Ixѱ���o�&��"�W�\���s\6�`���Z�
�/�N_ɪ�L��z��[���1[��ЉP�<�i�C�����Id�ܹ5�#�E��������{���omr���9���gH}��v	����mw�şT������/'��h��R�
��H��=ȡ�z���青D*7p��E����\�ӊ�e9�3�Ô���<@��|�1u��N4|�	�;�ch\��N�0_m��R!|1x�hU�aJ:���X���}�1��"��X��"�|��L���:~�2�oN��U+�-F�U᱅?E E�Ŀ��.$�{�j�hN�~���(PD4M>C�iG�Te���N��@|�u{�H?v�sV�J��~!2��.��i�X�aN�'�$Tg�7Ψ��%��!���X���@��DQ����e��t���~�SuЕSVU���Ԩ������}^�X���d%�!�C7�c����ܡkR�E�iq�ves�+��L8gąz��:�ABW�*�G�I�����:$Q�/b~����b�=O��P��;
]f�8y�r�(D����y��Łi����0(�;���3[[hy���� >���S�a��&���5<�D~�T��h��-�)��d�;�k�(�*���٣j�G+�f�SB�wQ���x�Ƞ3�,�?�;Y�(h�}t8��2K��_�2ݹf{���܁ѦZ���nع���l� ��~�QW͊.�oCj@s�t+�Nf�"l[h��X�:�"i�ˑe@k5$��U����'���i��k��Q�͆J���4���~��\s�-͟�:�B,�7�Z��f�Aq��.Vɷ��z5��@��#� �+*å� ��D�� PG���+6�b�Ŗ~�lV�$�2��y1I7�ז��iÔ�j��^p�Ijan��M����<��0d�f���X$�x|�'���%
��� �8�c�i�!����4F��˻�����\�V �����&f��w�*:�C�V������ ���k�-�ho�čj�6q��4�b�v-��o�ǈ�:�O'�vZ���0ǈJ����_���LK�Hi7�Р��b�l1H�7F�!ӛ�lǾ�b�t�b�mH�j5�ji���m��'v���nI�6�dh�U�u�E�m��"��i}�y����m$�����d9��~���hM��?�m�l����ĭ�0�R^����M0��T�QW:�fh>�L[�e4��@X�@V���'Y�F]���\�sC�K���-��D����$��Mv�	�(�@�̟l����	�n�X�;G��⋢S����HӴ�h�����{�eM ��k�#gE_ܑ��#o���f�g}�*B0��2���<ʴvI�t�K�8c�z�i7Ժ�ߓ����D��"V�sKü������lK��1uK��#�f]q���lR�����h0G#��<�t�"Nh�<.R ���^9��V�"�Y��8x���b'������65�n"O=\�M�=﨔�{)�s�ƍm�L�fM���	�/����+H�l UN�(�Mh��cO<�>l�v41�|��pK��[k�(��E��P���,c�%!Q5�����#�y�6�`�S��p�>5�[�N��螠�G7Bʧ��rT��Vd�Sa�?8��^�ך�ꡍqș�BI}� 7����a:�9���;���(�\��;<�d��t&�d:*tfi���X$��"Y����9���ݻ
E��/BD/���y����%��vɏ/�`q_p2P33�9�zU��c@
'�sr���`Y�L�r�|+�=1f3B�����uÞ.���8+�BNF��
ݬ��i����txI��F�=�ŊVS��,R�l�h�%r�I��@��k����}]�`_�<��+�Fy�{�^©�sJ�YBWh��6���>H� K���b���B�E�U|8�Y^���JL5g�ZU���Ѿ��}#�I9U����BK��-�#����GH�\�ᕄ(WԬ�����+WP3�;8"����)�����}�h4IP��� JW��4���]w�V �罇&�C�m!{T<L�W�7i�')��f3����v�*?����`������B����>Л*����6L��������P~�MQt�y���-��e`^P�S�h ���5V�!8�B���W� g�Z��˪�����X�����������h}��f��4�QdтM��>�1���B�=�xY���d�4�tU�y}֜짘f�� }><��>~��oف
���F'(~�Wf�,�#�cO��w�iJ��B�pa.�X��P4�Ց�S�ݲ�T���D�e�����pN�fmVc��#�C�*mLe~<�}� bS�;w継mG��U#���${�-
Ք�K����b+@����x�m�bj�Y5��*2�H�����Sm^�8ȓÆ\Kl�̒�@3]"ȅ18�ţKJ����sx4pg u^m��?��#�ׁ���L/�>�ɈI����eH����$��+�jJAwARm�/��3��������T�L�0��J�l�S_n���B�i1�i�$���:�f�ř����y+[R
�O�}蔫a����Q�H λ����+�,��1�sd%q"���B���DAn�Q$�E��#�K��2�� �"��K	 � d�:%cɫᴍ1��[�攽/ݛ���'{��[�Y8.ߐW��C��T|8�Į��d��%d#t��/���ځ:SX�^T�l�Y@���vZ8�Z���<F%�_��%����u�4��`�De��00 �Mݎb�k��,��gd�i�����]QUVh �J]�����Ď�'��R),!3�� C�yH-�W�g�����?����8/�Uz�{Z�Z���9���cG!�׼���!�ɜ�2��mY'|�?��JB핵��	�E$,RQ�ڏe
��cr�f��D*&s����F�;�8���y��nU�y]�9�U�"K���j�P��������΍��;-G�|>!��6��;���8�F,����0K��b��aD�d���
���6�9;�@Y�q�\~�:��R���A�Lv�2�u��⾃����[m� {1�Ҥ��3BO]�[��Lӂ�v����9�ℂ��Cei��TM�x��`Йg��H�R��lw��hp\��D
p�D��L�@����X=�����D㶐]��=���(aUV��t[��>�Tz"e�1WK������V�����tSn
�l@�&���׸ς�)���;��z(�)\��%�>1�k�;+l*�3&j����Љڋyꚣ�Eu��4F��<[��I�?�5֜�#�jGB爴�R\!yA��"��th��ժ��u)Gu
3
�:W%����X�q��(�
q� �*z�kr17Ƭ?���
�厣�x,4��|�t��,$@�Q;�����P*\B��H�|���A�X=I�Rvg�2oH�\?D�����(���#����T�}DI�T�=$�_��1�>��R:0B�@�vݨ'T��|��&<\�B�Z���Oł3�p��ISsi�Y��H[T��1�Q� �� ������*�\^&3�@�݌�6^	д�Z��P��x�z���@�~7�!C��j㗀�V��'m���vwJI?o`��Z@	�W �VU�> _�y�+�I'�+�#�"xW���{lp��z#ļ\ϩ�჌H�7^��hvKN(ϡP���w"��5���~(�$T����(�wl=��C��F�E�Q��:N�|����}=�$ �g؜	��b
��:�=����|�;���g	2ps�EwGS�,��'g��������7&�$-�$d��9
��#
��1fZ"�;Db+Ӕ볂,��Ί�	=�������Ң�L8��G����.�J=Bß��YV�yp%g�����&�]����ݔ�o�j�A��b}k�N�>v"�cf��ηbPLa_��P��װDj��p(yk�
_>�
Tޒ#�xn��4�_H��D��#1tƿa7r(ݯ�]a,A0'K����e�TNO�;l������w<���Kc�c���˦�C8e$��`�H�ţ����ت5T�~Z)ёv��Wۏ��������lUU0E�M����9d�F�h[�8�,2�#CM���&;�~�<~X��;)�.�}�yOaAv& C^��QG��a�?:�����|V�F�7�Z��a�%U(\���|[�cڑʭێ4��SF��7�Y�����_M^\��gH���3�p2A�$��)��{g`����嚩c(�����$@��"�҄elTD�J\M�t��!;T���7�z��#Ґ�wm�(��x[ɐ��_e�C\�j'��52Y�E5vE�x����>9Pcx"�r����1}��]�+�9���b�z�3,O� ����AdC�N2�Պ�St�1KrV./�DɔF�i�JƱ?��]�R�?/�5>bع��!�8��s��?��9�|5Ug�]ưʺ�
'�@U��R�N3�)��_sA�	�r4�x�<'T�a +2cZ��^RL"8]�G�;?7��>_�L�sw��[�BE��P���p��$=z���d�#20	�qD�N Ļ3�� Yg�6������MS��g��U��%c��m����"yo͚�S/+y)�@�vK�ms}@�1Z��^#�b�����r���ճ�]Fl�h&pM
�z��pB���[�y�p���/�6x,Mm��2��tK�I���vd�Y�~P�E�o���T#Z(��wKO�"�����̥�Z�8)�-,���mM�j��t[7���v_�A4a%?q��j��>ۘ����:cLn�|q��@����xP��T9��s՟����aQ+������㦆�@$S��	C�ѱ��V`N�ϛ�WR����
����R#�5_N�J��ov��
/ʯYG�߇�tu'ߝ>��m��$Ciz8�;�7��v�!�Ob�y����~�i�Q!ġ�'n.����3����$�@�����l���I�ނ-���0s�[a������Bb� ��d=C4	l��/`�z{C�*�z�[��QEǉ��&��zp�Dmֹ�Vd�,�xL��5$Z��R�`�F��blu�4]���3:�s��R��k��%��v�Db
�$D�G;S�[g~�k�*R�»�(�c��XP.��ݙ�J���]�FpQj��Jx1�s[�)���J/����靁̔�aRHu���q8�� k��׶˷#���ؘ��Fj?fvZ�XFC�r�G��Cl¡$���iO�LW��X�~�3��텏����l>�9��Gw�X%��P<f�q��)�����Rg:���'�,���)�z�F1~�}�MU��$\@z7צ�F #�6s����b6/v�$:T�N���-6�x��NAƬ2ճ����ǖa}��x�� �c�{? �w���#����C&�h��N�3��+u�{'�1�/�Y W~��k�i�<l?dq ���k��X����\N�zf�pQM 5>r��S�w�ָ��.�71���>�5��vrmH��`V�/Zp�n��ys&�L7�@��	��u����z�
Qk�A�CW�ysGU�6�'����?�	u�\:�T�]F�'��!L��b'�����X�s����(b��;�~m��W�XT�I��я�V:zw�5uj1E��i��d���;Y�D�Q��t�,�	7�0N�ˮrB1B�c5�N���D���q��8��Tl5r��f�/y�qx��/^��/\':�e�pP �������4��Z�p�ۣFz~�N�o�B�J�|��������&G.����3�^����l=�0[�ʴ^���4��(��L�Uv}��8���RP�-�yn%��n�� �EI4Seb�� z�ŏ���jd�|Y�+��%��D�⎂(���R\���]Dq�E��5�"�zv�S�X��L�� T�Q��O�5�H|�UT�>��o`��ڗ��k°�K�@ �J	���lڸ�P*a+�M�Z�Hn��.Ϫ�v:C��=�J���pa�0!	k���_�d/���^JQ��2�,��k����e��؅���!^��0|Td��6s�>���ei�@rO!�R�D��}J�>�{�b2�}7L�S1^����i�~8\��a�N�wn���q��Z����w�k�:p'�J��&ђ��6�|��������{OP� f5*Nt��i,�@	�o13�n[;�F*f!�f�y�S�A��2�b�ƀn��bc�I�l�������+*Jo<�^�
\�39���)�e��K��xž8㪄���h����|��p�T�&`iW�����=�@[ĀX^g],u�r�:���GL�5dB��I�m�����,��]���5yĸ��m�߱��5�R�c�jEf�L�7��Œ�� ݶ�N��C��£ª�v5��vߪ��VA�K솤�9rG�I:��/}�����Ml>�I�|�O���R �jsؽ���?�A K�T��؋|&��l�N2`���]W��h}S���X��(=��A���]�EIAF�F¿F��8`�J+�U�Ɓ��� ޡ|�:\����y.̀�d'_e�����s����ʜ�:� )!��R��=�A�F_-{�������Ԯ3~y��������3*��6�w���'�&}PQ�J�=2�i��+ p���"M`$�d/�����[	�:'��ҭP	,Ti:a3�0Y~v�>���	ο�� d�D�,����%a���髡�������L�Uٔ���S�qW���G�5a���d���q�J�&_޻����	%gB6�U
��;�P����7���[zs/�F�	�^��=���	�6,��}�j)�I#)ĀaS��kZ*���;)�D��b"RQ��,Fg	SPRXY�ڰ��Ɯ�w������ ���x��,Vu�6���=�����|�S��`�@G-7�P�Z��m��ɏ�o��Z�J���q�γt��@w�_:���{h��ױ�G+3����:���U�ͧw#��:��0^!�n`��"��tТ�����o/�-� �"�KF�
ܶ_�Z�>�0s�m�K ���'��y��k���3���袐a���Xq�`ڑ�{z$!���P��_8(~�+;�l�,¹$k�&4�A�3^l_�u��kYjAZ
M��^M�^���U���ۮ¦���`sR��U=.�]���[ׇ��0M0չK<h�g'뵏Dو�t)���2����_�_7�4=��P���#EL����ڧ6�|�]2J�����  w� z�o�BߔɗmA���^КX��dA��h1��j�ZZ2�7k� ���F�{8�&]����*W���ҍH�(�|���-��+�z8�:6�ͧy�p}���:ö��%Ւ�� }l�/����(I����S�u��H�_�b�-ǽ��żH�|��HH%ً�g_?�*�G-򋇭���JT�XH�>���g�3��3��|���l��n[���?����SF��1K,��/� x�{�l��Wu���a�*9
�����j;�'m8[![',�∞�/�rq��F﹙��P��w���ϡP�e
��~����k^����
�ɥ[��{��F�]-�����r��o�n,ܟ��z�Lw�C�$1�,Z��@x=^=�͘��78���L ����0�_9_����c���0��)��,�CV��S4n�XhLz�T}*�'+u`qk�����)� 02~� �>�ݕ�/X4W�;Ru��
-2�C�w����bm:�g�os�P�.[�#��E���� #<���Q����$2RX�P*�-	SE��[�01�Cp�u.� �-�-x{��f�W��Z�Ğ��(�qa\-����d8��9A�3w�Q+���I.��
�ר_��7u��Y�RՃ���Q}ݳ!:�^T���G���0�$>j�si2!	J/)"H鄉)�gҷ`B��E8T��m���a�^��a�y�-����R�������"����O��)Ρ������.o�P�|�YWuz���%�:�l����G�&dG�X����ڜ�޸Pl���uh� ��2�<B<����G�ф�QY?\�݄�ؠXQo�<�5���-f,�e�̟�'��(S1yA��=s<ɫ]�����G�꾽$yg��8�A�pcؤ�5R�*.���t|��Y&���.�~5Yo�)��e|m���fi�L�Ԉ�=���Q�2��5p�/:0����k�uݵ�H|�D�,�����_
�a.�Y		�u<�~#��͇�K��<���]:/�/,�`5ɏE��f�ΐ4��"���F6��֌ո��M�V)�p�z-@	������`��Rj�]3�J��͏J���z���LM�_j2�3� �L��[ }]��,����\Jxq	E�]��)?	�L��Z���n��S��d;ĜF�c��Dyl�/�f�t$m��0o���/ӱ'P�J~�KU�OG��^HB;K7	5Ɏ��~q)�X[�!��)$����Px���s�c�[�n>/NDC����U�Ʒ�}1�dU��S���^G~Ț���1Q*�A1+{��-�fNU�޻��l���B�I:�D�TL��8�x��Ը�b����(�y+���;��0	V�FT.cA�NƸ��DJ�fv�,C��t��	uD�e�z.�/7:��R�����%a.B�a3 �d#w�Ι�SBan�V���i�v<��b���]~����Y�~\{�� q"',�"��*�1|�"ai�|�V����(���ғޠ{F�O�3t�-?6�X	�����o�iImkB��#�Nrby���w��Sк��w���X ��.��}!#�e��aN�_=�T�@��ɖ��"��%ϊ5VQ0/��"��᪤nWy��&�/;{�z��B����/똩s��L��5t=z=��X��uBc}2i��F���g|����9��f��Ɖ��.�FO�@Ӹ���!8B�z��m�+WzᅘdU;��F�Ԃ'�Q��6���?QMw�;��xyh��i';�H���j�,����|5�g�x49aPX���{�q35r�ç��n�� l>�"�"&�#5����Ԝ��i X�/�:�2��·��9@E
�̷DB����S&��W�7�y��s�<+^_�1�^��yIy� ܊����O�D%>�lH��_uū���P>���&�v*�b��ه�Ct"	҇��]�ʮ6��<ŉc_� e������)),4"���x�Y)� ��i�e�2yׯt�AĎŖe�N��^fˑ�e�=$=�hY8�6��+�)�E�6;nN��o��gM]ymJ��pf�p��N~���Dp:m����_t�o�,���S�����J(d���_�N�5HgL��q�0y�+>��:��(�R����:Le�N;B�#��Ǣ�"�F��%r�r)K����j�-9ѽ����B�w�����=�x��>�0!t/�	�s�ɹ��t�X:[���"b0\���xn�|%���YQOJ50Q��\�E�w������e�+7�-c����</.a��!��[��o�'��_�,1uz��x`_{5ǯӗw~�{ᖉ2pz����@s�mg�GUԶ@��Q��P�Bs�q]հ���C+�|g^iӳ7�g�1�`�m3�
�C,���:*�Ak�	Qm4���L�&�qk��`��i�b'$ԁ�s\����)�G�B����^���{��̃mI�����w�|+4S�6S_� gvQ�����d{_�%�t4/�����d��dOeˋ5����r���1%���OBG�8¤
�~|1�"oe�%ĿC(.rRQ$���c�i/�c��v\;{$	�C[�X��E��_,��dk*#��Ű1ɣpv��9�M�ǈ�M��ƶ�ڣ����rH���H pG��j�UJSf��e��@��d����@U���܀A��V������g��nP:����d�g��@�g���jZ��S�g�'�ѝ�i�0�T{.����F\�v&J3=���b"?�iWv߾S�l�_�TGn��֌�����q�zcH�H�4c�yU�^&ض'Y�����6{�}u���[���_����yMhs�,�y0@��-} e��?W	d裿�$�`4����2Mɖ���'\3�����I.����h�o���h���4XUT2�a[$�%��mr%u��n\�>*������$𦒠n����Ţ;s�O� ї��r�d
ѿ��"�)�ٿ�S��Ey�Ct�H5\�U�򾘂���\I���9ć���<��Ӹ ������=�AV,0�m��9����9QFq����Y�[���a�?{��a�Z�V��i�fU�� ���ߟ�#r u�]%�`2K.���=/��8Wf��o2HQ�H.���o�����=0�\%ܜ�w����t[~2{(vÛ����丩<��ѻ��+��h8 �B���%�Cg}�ek>tMn=��o4���:?��✵>@���jJ�(~%���l5A*+ �&�ͥ+����5�bަ��F�Ӆ�m6�V�w��HbԔ������ǽ������?I��S�j3�dԃ4K/��w}>�	�6�t�P$#�ߜ4?hi2�����R>|x\Gt������<0��Q�A��T]�w����R�p^ח �����2mCr袋�UX2�Q��L�t^��#��H˳x�X[���L(u�[��Z�D������Y8t_N	I�^=�	1e���%zrް�1� x�H����y��MV:hK,���7\�M8���͓P�$���D�N��!F���Vg��S�?4���*m�F�
�n\�#cU(�J����w����P��� K��'{9Qo����A��!Q�O�'W��#�< u:��t���Nm�[��Q�b�rx���)!�cOkJ
\��k�$�sV��]��y�Y�pb�{��_��}�!��kt6�)�欥�_��@�S��+d�K���z�Y��)hƮ�p��!�t �i�L��fo��Ǻ�W�_���j%8UB7.�_���3vz����e�a"�4+��E�d3)��=U�6��1��ӱ�Gɩ#�M�;"dӿա)��*�;�zN]��M��I��]��r���$y^���+ai�숌j�K;���L����X?�)�������,wgbc�(�s�I���S=��3��?+����&]���kT�V��ѵ�Z-����������3���p��0:�E���2���
����'Qh��h^ܝ;W�5e6�lL1IcYyx�|�B��!���:.+�ހ9�'W��W�vI�E���M,E#wC�%�)5f��G ��dS�d�H �5�09�;�c�~6��\���e=2�L�Wg��D!Nl��w�bA|W�	�)���^�w=1v3�?h�~�*|8�5.�.�c�8~���	6ă���;�S������@F&ҩ����cw5 ��Hީ�%�'��}j[�3g[��J9
vTs���ۮr��%�^�#���w�`�����:Cd��"�= �]���X�� ��п�O2�;�3"�!�M"�<E%�׆*�9F�x
p����
��ҋ��7+FRJ�Y8AJxTp��a,���O���	y~:�^N������W�}Q��n�3���ه��������M���y��X���/Z�L�;^6��a����*B�2g&��%HL��$v�W�.7|���l2����+���J۩Z�G���&7�'{p
��6^J���ID~���J$� ppm���H�H��q'�&����M��f"A�O�䘼��F6���f�� ���/���'�߭��?���X��F�`��y���.�W�1�Q����0}6�%V�^�i\�g�.g��B�Ԣ5n��L��;F�*�;�����5D��<AD�;1���G�	�/Ĵ������$�[�:+G��'Z��*(���+=aWg�*gj2S5�332b���F�4��
���������4�j�z)m�3v�IG�~�2�B�0z�S��ͱە��x�j�cU�e{3M���Lٷz�3��.g���5�����ƄU�V^`��P�Yv���Cr��.�)�Y3��`��[�zP".��U�ھ�s2��f`@����@����)�m��� �-2 ;j8n��2�Q˰*"⣒A�)u����aSH����ۚ�������`҉f*�}B�?��׏�(���o�����v6i���H��bqP�r"�T�����Y���+d��}�\�q�u�X'� �E~|�L��A3�,�P
�^w)���0n�.�_�.9�*O�w�_��ߝ��X��z�Jfs�drQc�����H֕�i~���t�����K�QR���n`�&���X4����u���h��d�B���⯱ي�k~MΕH���E^ݕTd�2��J��tΡ�� T�*��Y}�握�Uh�bl)J�#��k�@�E++���bn(�{��ї���D���x�2yG�ck%,.�wg�t*�}�c3}�P�$8渀���]\���El_�<Vnr5�(,x4{�S� -W��JRS��eq%�vo���h  nF���<����u�)�ه����W��Ej[{D�M'�a{��d�ikO]['�l��~��O�˜�p���\V�W���.�$��N�Fq.n>Z�W�����E.�l�ƙDY����k�O�����{" Q��������H���l����,my��0y&�)U��7Z��9Ɔzߎ��kP{�57��hJ#��9��l�^�����T�������ha[�.{6����{IP�f�)�p��N&SH@��|��9��O0�l��[�l�`#,��	y�Iڋ��U��/�Y�y�_n	�꽗; �ӝ	[�~����:�1���7#��x�A��A����z�.s}f������Ҡv�Šd �������(*��B�;3=+�O(k	c}�_�<��kVq�K�X7�Lz� u���i[o$��5�4�n9~�p@'S��%����4ص{�|���-.��z~��n�0��e�6�P]�	�����Y�A��������� �/R��Z�`t�!�4����2�{���[��N�Fl���ec���	�3���50`��o��ϯN���f�riѷ3��hK��O"T�1
X��0���P�% ��0ԙ�F$&^d�~v����Q�TE�}
_�:0�a��蘧����cu�g���lJ��zl��X�&�������(��C
�&�0�����=R.v#`u�E�G��r�������r*sd��7?5F�0��L4���\��"#�w9Ֆ�A7K���<Z��q��#�bN�#��Bh2���TX�?[Tn6��q_�T�*g-E����63-w*�£W[a!��"~1�@2�ˌ*��G��[}�m�Ԕ1���wq�%�u'g��Ҭ���c�s򷥾)�B	t�r,�,�]CÍ�קŃ{Fn%t�o�ֵ�2l �F�$�i,:gz����.���@1i��!����e�S}`�ȵ�N��.�$zj����	�v&8��_�F���1�ը_ٰolp}����b���<�j�	)�A������]�/�F�)x�a$+տ���"��YI��"�r�]��%�D��2��`�  �@��3�o#��9H7?��<	M�6��rXOO��I��<z��[rDو"i���2�����D�/����{����ag�n99�NxSK�wU�1�;`t����d`v[.o+��f�cr(�,q�V�o1]�Y
���ȏ�l��>�Z9�n�2�Iv��Ne��CI;TU�B�ڧ������v��P��E��nb1��L�v�XsX�I��-���'/.*�؄�b?�Pw0o�o,�:E��1Bؠ�)�����Y}E�w7���a�։sR��> D^��l�����Y�k�����e��>��3A��@>P��}�8j�MΕ,�
d)�^�/zxا[�I�������Yk�S�u�d�ڸ=_����U��������ī$��wE��0�xo+Y2�����Dč��n�=�(B
i��e��&�t; �3�������Dy��eF6�S+�Y�a������=�!Bb��6�7O'�F|8��OA\?#EȤ���x�J�C����sc<�>�rvk��bV�k$Zǂ��m��:>�[n�Q/�V"4Ac�`�����[�_�IO�JIBs�ؘNc�Uz~##7t�BHЛ�eX8K+>�t��ݴ���O��Ȓބ��QY��c��u:�
S�۬po�aE'i����p��.�5��<@�.%���=��@JH�~�������z�䗘|[�)H�_P���k̝�o!�"̚-[Ac-���&[d�%����w��9�Ì���ǔ0�R�^k�{[�
e�^*����Pz�iг����Y�	l:�r��r"�\'��|���7�0�{�Vd�f[���f�����g��T��~���/�˶�::��[����%�Ƥ�@*�8+���������¸p�
�|�-���;֡�l_Ψb�Y������-T[�
w�|�خ�ӓ�V{ų�FR��l�T��
Y��eEȲ}jR��R�ϳ��!�'����h��P�$#��t�C�X��b��m��A_�6`����W$L;ӹ���=��g���/�
7�V橺[h���8T���O��ʺ\k�ޞ�A��KWMV���B[�TElf�V�R�A��u�`�|�{��J��S��Q���\�v#;�ͫ��N0+�d��س�h����բ�h䶝
�㎱19�sj.�o�P(A?i]�L��>an���p��
��V�^[�[ظ����g n���WX/&Q���C��}�O^�4�D��+�)?������K�gy��)!��3����?A p�{�&�91�3���R4�18��C���Tgm��[�_S�E��u����xZ���YG@ւ����������ر�U��E����䐛��� ���6�?��@{��O��g��Җ���D�(/-�AlP֊-D�l�E�dj���F|h.ۄ���%�C#���x�˫n�$]�,d�!��o��dc��ݲ�U��@��P ���:Wq#��1��vA�SQ�w*�BόB@�w1Eb�Oߝ�R�t�g���x�܌�O|c���y��n�FyI�O���UFL�,��x�m�}e��r�~��.��hYW���	��~n�%>��U���	�`Yp"aE�o�w_/9D)$�UŊ�D���4��f+����|����2�x��: ��e�O9ou���aQ��yl�#��	��G��6Y5q�������
�,۫��ڞy�Zh�;��H��g_�F
���Aa�VٟD�c�4a",�N�����;p���~��ɕ�'o���u�lNI��dZB�����7�M�S�{��D��x� 'W����c-�N�5�C�(+��-_���1��:+�'�vJ[L���Lo��tz2�\
U��=�!x�	������Wފ �8��<�uA�(&��pH���|X��zx��"�V�E�H�����	�jӤQ��\aW<=X�	j6����0���1J�;����������z&9�v�����اt䏊���9�aJ��؜꽀�� [�Ё� ��i	%Ǐ�%�c:���lfR�ل�u�E'����t���C���x�s�0r783B�J-�0>s�TTK{<y�#���ú2z�Dx�Gy~�sbQ���|���줾�\��ku��	 ���QK�n�pA��csT��q��b�|��♫�터s�3M����⸞����c)��"�ʢ�!�o�m�bd�]}��:�4��_ Xz�0����W�D�.��-.�Dތ�NM>s~z����u�+m� �h4�i���-O�wut*R�j�+S�&!�ć�P� �:�M�Zt�Qg#���ht�:l��������8��i�U��V�;��ӏ�Q{`�3"7s���r:HO��5��og�Z)66��5(#������Ūk-��kT?2G�ps�T��s[��ꬿ����,/���T���)6p�zg���Ģ*IxuVZ�.�w2��qW�x���tP�	T���R5�BX�T(�R��!�� �&�p�|�֭2:�óU/����ܮ�"|)��)��PA�X �*��f�0���=
���J�ȯr�v����~Yd��`$MFr7̌�\F�f+-@[V4�hD���=4F>���<�*�`?�<�0����
FY|���1���ς�I�U�dGe��r[�&p6ZƘme�W��>fA��ץ���:�W{8	DS���Md�.3�	�3�K��#<	�J#�^.D�� 0G���PB��`&9��47�D?,�c6~8K�����"�baMU|�_�%�=��hS�Rrfu@|d�Ν�%*wч�Q/Zͫh�d@5AzW���+B
��}]��plvS�I��"A�ۄ��5�O*�����4�������(��=�Y~z PY��-[ uʐf�क|I�
$0��&����W���i��"�����hViR���86���&��K�I�-y,6�C9�1L��^�,ul���AM��jL�(�/�*����:D�~�j{��R0�I�\֝���D��5���Y�_烙�p�nh�9tJ�J<���A^0A�Sp}Lk� ?��Rb8����c(���W�1V8���]�A,���W@~��Q�1Esj�s+�Y��-�͉��[ε+�"e�$������������!k�&7YP�������V{�]��R�Ss�0 �9z+�M��"�%Ϙ}�Ec����������[^o]0=����zg-M�8:�s�I�/$�y,���U,�������,X)[z�kX�(, /�2� VE��@��2��m�Ws�Ό�����Z6�L��vճ��ws�U��ug;J��lp��$(��2�b'o��Cml�ל�5 z21��9�c�q{��,�g��3�/�XX���U�)δ_a]>R����9\x�ː�]��{y2{Jzc������a�7�5O�~�"[c��-�F����:����9}W�$`t��u!?��ݦޥ��
�DzkE���#@���]t|s�-#��5D�!�s���I~��{U�?������iO���l_bFb�`��D�-�#�:o�2�<��×�O��v�i�[���$�!��� 8�1� l_S\��gQ=},���z՛�����@͌��&"a�����)��ǋD�Y v��n�d:%�p6�)�šM�ϊt�1���T�I�f�m��5M�H^�e��9�4N��	s��GT�\���gg_��J�V�klQ&?a`9�FY�-B�ѵt�z���d`�:��~m�FI�ʔe)x��(q��j��Rp�\z���ŮI�]�pdҸ�l��m��i�<�iO$�mΌ'+^t��G%�s);aFL��z6|�{�sEEܜe.!�S��%�;�ג1��l����Q&�,=�Z*67�<B��1�N�ʔX���ɁQ�Gk����?&�6��R�J���'����&��qİ��9��$;���ʳ�o{�l���ۻ� �N�_2/�Zc|�i���?Ft8�b��Ϡ�!�7��Zi����mC�z��v�#�iN���D�ն�'w����I�	��� `-�}PH3�����o"�`� p
h��s�7J�������m#�!=��w��-���W�E�A��s�e'��Q�q��O0�C��}]���J1��.�dԖ��B%�3��w>'D��[�b~*�$Q��l�Y�		.����㯄��E6�{Q�oG��ݴ��Q�ri�B�ڀۏ�!��VM�4l1���XL��Tn]�����I���f/�OP�t��/���"5��~B��Z�Ӎ�X % ������v���lx���+�2�c�S���a~`oRk��P�xSsxwI0oR0��Xzx�y��������r	8S6^>�|�|�"y��P�ƵhKE�ش��O���ʄ��ѝ�qr~歏����ɩ�+�S�&զO�U�s�#3�A�,7w�"����%���t�Q�@K�ޒ�;q>x��y���pF����pdRy�e˖���)�/o�	'���/�#nx�9Ijǀ������hޥ@#G��a�O- �wΖ�j����|}L���ʮ����B/U��E"��J]���O�vr���z���eW鷞����E��Z89�SH>�4�y�g��H\y�|���'y��q��_��	�lU��v	g&���3��E������H����7{ϩ%Oes��Yj Q�,����ҍ���q�l� ��4�?�c�c�" &��OG���qr��7�(`��YK��e���x�t�������0i��·�"�:�l�s���1�S��#����0e��,Y�c�~V�C��7��os��/�T?� SFʍ�2����ش��Mx�v˳��M"̡��6?A>�w��TZ��_:r�)�;�K�}��#y�k�K��
�DL�||��@u�_ɚG��Q�-�k�<P��$yUoY�Q�8�������e����fZ�W���8��vj�\'�	kĉ@7��"�����3���L�(cuq��;k�`�v��]0V��%�2k��'}9{Fu�� �m��=����a�D���k���^���r�'�w�'���	��Ią&ܶ���ŉ\�wPpx�nE�K���y7֭�Y��Ҍe��,�1{p����`�m��uZ�}$.����~'���"��L�d]#�B�'��x)�.�)�^]m�eK۳e�����DSz9!"ߏ�4|8�-�Q#afi} go�l"�����'|�<涪t3pHtӻB&��1��T6Z�IS\�Z7-����	2!|6n�$�;���  �L��ߋaM]z@��Ύu}vu�Ҋ�
�t��X�^'Tnk֞{0���:��BD���I��# ����U�41�=zv�Hh�k���Y��5pRP�-�#�r�e~O�.������mu��a#	���a 0iAL��|J�K�:�9�4Z���kk�g�eKcL��ҧ�h&�+P��N��6.0�lgp��W���4�c��,���t�փ+oD���~�N^�OJ��t�w7F���z$�D@G�K�v�ěvx:��&@�Q�Ď�m�� ׬��u�E�T���[�^�(HkX�Y{yt���T�9MKa�j�f�.LR��uj#�2������4Y���R~�� ���Q`i�B��wYi|+9千ko���`WtOA��-�\1��X�Y�b�:Yh����!ɱ�O�K����4阂pjS�I���\]����a�[^�RqX=�M��#n�bE��)�J�t��9���W��ز|�� 61֫��B��H��n���Z_~�4^����wwܺ*�ߑ�c����l0��?� J
)B8	�v���TW��ʩ{)�֣rHD�<B%l���_r�Y=$�5Ω-՛�w�
��~�)ݦߐ�`��?ѬO�����cdt���~wD���@�%��'T��;���F��!�����V���������+��@J�YI��|�C�Y��_�J��K�Y�#���?��E���b���L��j&�I@b�y'��3��ۜ(h!w�rL����J��T��6�U##�ܷ��rLw�~Čx������w�����ːE�����ב�t9����C��QQ��'l��Rt���d%�V�9y2d��yߡo������@H�SV+u7�À���$h]��ތ��//�\H!���ᓿ��֗�~l��d\G�6���ˑ�(��aD/�ݒ�(:KH���〸~F��翬ee����dR]��|@t��.���$Q�����;֔��@O�c{���X{�ա{o7��V�C�+�� $������Ctߑ�q ���/��*
�W45ƕ�|FDq�"��)����ߋ�>>�۷�`���x�֞����3�h(�d��.'���3���DMp	��%��^� N쟂�lVkx�>��2�q�#�����ڝ i����P�$^��F�n��m�T����Ǳ{3n+e��R8�*��`�H��O�o���#�]�J���c��O���/�Yhq��X��sSd,�{2�# �vzR �����n�Ն���X�ql����JK͜��S�E\q0O<P��|��V�Ni�t`8��*ԈaQ44#[K�i��όʔ����l9�e����4�d���,$���S�8ݙ:vHɆ! w�����9'���� \X��ݸ��F��ަf˓u(�e/yV�.
��PN@Q���%�����>�OH���D��ې�E�"��v���Q�7%��g�hUNɬ��Fң�rePh�5��MV�u�3����6��)�i���3ҡi����Y�}�I�[O��hE�O��5
IH����oOUBj���p�wbYO_�}�M��Y˖J�Mlor*��*9�q������ J�?;�N�ሎ��$Om����P�~��}�?�(�O��izc%��5���М�d�6�z9�gw�SA�!���������=��9����q�_య#��T^���/��P��V~@d��g��㇥����P�XJ��mq��1�Z0� ��#���_q�u�;�I�eDuKN����Ͽ,�5t��;i����oͥ��䄺3���C����ua�c��&а[��Q�#0������6��OC�Н�.{g҉�nĢ���eȼ<
��=g3��޺���\�͂����7RV��;��o�[^ͫF��&�X��S�u���>����dG��� ��:���#⿤��Q:M@�Qh��F��a� ��Q��H��o�y�m8]�R�83�F`�ہu+���:�S�����ٲ%0˱�@Xbv�w~Y�b�n��ԴCO�s�To�Sa����f5��F�I�x���s^������m�\����U�W��ŕ�F�w������Z�6��A�J�(W���4����5
����M/� � ��O7��������U��1ԁtOe��X0�^q�x`j;@��ej�e��q.^���������#�u�È;J�篙!�/��� 'V���XPB3��g�,�O$T8a�sw�ږEW҈�e9��vf����J�9�ꒉ�"A�X�e�*߇�!3����^R����zM�z��>�^Jե���-�vb[�%�=���DA�=-s�k� W����6P�����0(w_�b�"����)����/4�l`�jc��֚�
��6��PE�v��˯����.�.�
h|�)��'}���b�%����͟��a�����o��y:W��ް����y��o��]�Co?4�'%��{�������j�ZS�έ�̾��9	Nu��6\�y����S"i5|:����u��@���T��ϻ�EJ���oZ�u�]Qw�����������\5ݘH[��Ve�	���1���a�2r��ͣ<��p��?���DV"��	�E6F���&��A�̬���	(_*WJ��>�_%7��m}����m%���*EP�L�<�`��ҷ<�xvg�B���PrBBk���`9��mm�A"����&d�ݫf��^��gb��gD؁���FT	��� �.=��QO�i��g=���i�y�-:S'\,S�������p�t��}�������|Ĉ6��4F0f}0Oэ��l�o�� �"���.L�jzTT6,�*��v�T���H��*���%�ր$8�	T�%��qC(�O�[r�ݲ[.)[�Q��x�6��5F�q���:V!*ngr���9O^�0�mD�� :F��u��sDM&N�v��>��,�V�X`{g/�4s6��ŝ��t.�M���U��x��EV5�P�,�<�����[�I��:���9����)M��J# ���ViLG��,�e*�XRp���|㽂��xh�S�M��d^��oe�/n�_��+C��0��xi�_n��&��$n*���U��$�.	Ikk8��r��U�<��R������9�T�����
��'��o}����H���:
Uq�߭�O�B���	�p���I��c�UF˜Fri����1���y�J�X�5�Ϲ�)
nJ�<�p�����_���������됏�b&�����i�b�sݮ����E�W��	����:���hSlB��g�XR�%0#VQ�A��t?vշ2������Ծ�)�e7
��u�d��bR�dx������7������'��ХQ���{��#Q�r�	V�˪4���JA���y'CgVҥ�a&T�qM�e�&J�2�1.}����=��i�����ix-
|hh��2%!G���рRB���`�W�I��U�i������^F�V_�+�p`	G�F�U�ofG�����A���_���i��ճ��iy��{�m�ʢ�/���Ti���D	�
�= �P`��o����W��S����2�
�BǸ�2�y���;U%��H �Ow�������k+ y��E�i�m��Y)�M�Q�'���E�(\���t�WJ�
;�;!��J�����.�A�
:������:���y͖�4���>D��l AD�V�-���{���-X��6��/ �~@~���N��f`�5������.QG�D?���p볭��k�sՋ��y�4��M�7�������a�@��|%i����L�UW����gΞ�����;�������.���ѧ)��� ��@O��N����	]xMڱ�UV�e�;�K{�+*V�[��1�@ɀ?��{��X��Mr��7w;�z��rF��:�ThC3c�(��������U�Pc�lG�D7>���������A
�� �V�bډ4t2o)g�M	.�=Eb����{%k��ksd��'e
r��?r����U���o�Lc6��G��?�'����W8�+P��8ν\��Y|*vg@+�\�ײ���&�ܺ~��R���vkZŵ�>���"}Pwi�����ٸ��ҥg��H��6���{&_A���@}(p���D���9Ҥ�H%�����<\Qw	�+~_R~�N��5.Rs���36�ʩ4�f�eV�k�z��K���.�(T�S�k�iw�����3:�3t��j��Tʵ��A�e��)���%l���r;؍o����f��L6 8�dxń�pK�ٞ$�l�`�{�R�MU���u�8��apڜ��f���q��
/�a+����ɑye�䩁΁�i[\#�<��țL?�S���- ��h�{xP��t��`AU�������;�]� �!:ȭ�̹̐���x���>dbI_�x�!�lǚ�N��������X�D��V7F�-����*4�K�(�2l� ����E�q9�*�,�:�T�P���׸�+��dWWTQ�6k������%U>
һN��f�o���I�����p�sza_��Ч:��Vh�p8�B��T'(森~k�|���5	:��PM�:w,�k�b��k���M�,�|��_���G��qi��U��¼	tl�n��ٍ:��n*����eu�v�Z�~u=��P"�`��&���_J�Fy-�;tq�V��S^B'V��^Z�}��Eа�f-��&#3{3IzIf���ѼR1
-+*N�OG�p���^ԧ��G��z�\�~���T�0�r�<a>tn�_S�xu�s�?<\��	�#w�~�|V���2,�
��s���M��J�a�)�g3�H矂=�_E��D�6�mr�������ԟ�ʴϴގ�,u�Zs�Ȯ�C��٘^R@V�ۧ�Q� ���d�rQ%W�w��?� 4�k��+��F��M���z/%熐.��F��ޥ���?f�0��L!������']E̚�8$�)&}7^�D|�nfڮd����jh��ȱH�v4xi1�0N��J�� �5hz��ZO�Uk4Na�9柙��p�����Ӊ]�H2���zA*;���>��~sucS�\ǕԄ�5#�W�ᰀ�O.�8M�L*�R@�N=�/�>Ϙ���34 ݶ�ZK	�mP�H���B3�u "�T�ߦ�U[)�2�n��m��ztE$����a��w�޹�pJq�������`bq��6���?��na��-���m���ڿ����d2�l����^5��M�/O�[��)��ȹ��W-�.k�6�艋���-�0��B�[�_��D����\
o;Ub��҆I���}G��*��͋��k.�0���q���eRQw���x��y�1FO�^~��p+h�[F�؈m��%���oE�6I�|ǗLT�`�$I�`��{�s5�D��L����~l���'s&$zPSH��8��F������2n\;#�|���$� ؠ��u�l}[�]&�y�2<>�j���/�/��qQh���(�8C�I��Dx���I���A���/��h�<r�i�`q�I���&ŉO��mk�e�D@'JO5L<η�R��Ǜ�����,]���J>F���s�N`��: e�Z"�0�^��n�
Ǣ cM���N9I����,^���}`����ogF}�'����&o�o$o0��?m;�H���y���T$���"l��;CJ�\��1�%peL��0ӻ���EЖ�k�m��3E#�i�B��m	`j�����;xȾ콉x̹�ݖ�M������y�ˏψ�ɒ����\SZո�tC�	E�Y��/+�VOG"t���T����a:�:�n~�Dk��؂�H��[��b}��UW�?+7��h�Ӧ�~�>����@`�t���w�V�<XV�.Wݬ�"�8�����.��7g���U=����N9΍Nĺ��R���XH���~��4�Y��`��8����?�I��H�0��z�i�u�[�G/aդ�^�Qw�y�C�ߪ�Q�uƞ,A�py�R��7(��O!wå4�
��K���?��v�]~	2Ĥn !��ݡX�ߔ�dUH���O@D6nE�s�8ǟ��Ǵ��X�9,���K!DZ�,&|�˗�VP�}�������Mn�g5��Oַ��ǫ�����۲�~P;��q`��9�i=�HA�(�e�y2b�%4/ɕ�Xꈂ5f�?��ɓHp��s7��h�驾~Lg�L����|L�+�-�O�d4]��.\�|OZx��7��LyWr��b�-��܇�*���`�O���@���i'е�9�F�����S�|���?6R^�,�4	��#�z4�1~���@�<
ݑD�V"�!�������p#-���Ap�X-Ip��3E�5��#��_*y�#�K�'��؟V�S=���&�љհ�����w��䦱�&T�ϝ.!��h�`[ˡ��X����K�O��U[ⳮzx���G�r�_���Cⳟ��PJ|o�xUȫ%D.g�2�Γ�n1��Z�~���[��{��߶�����}v�3%Қc�?d	qeK�I.��-6�A�r@C���-`�#���J�@"�5F���dI�0��.�=��p:��^��i��Z��h!�#p1��BN�厱 �4���b�:�>���G�S��_VI%+v���jC�O��"zF��Y����/��HK >г*r.�>Yϕb���'��=m7?F:�iv��u�,�Rya�����W1Á��k燗���XʯH�-���c0n�Ƌ���(ܪ�+�<\��g�z㺭�x�i���|��3g�]P��Ҙ,��~h��,6����x����^�����	�z�$)���cq��g�X�l*_x;�H�:˶P���|;mg;1�a;i���dӤ�a�y�$@(7�35�Z��$�r������_�
TiDd����`���U�HyA�'�B**b�0r�U��҆�3�q�L�2`��.���6���E�����H�Rm|���zdXm�� �'*���[ i]�թ�Ϟ_��#;߾o�r��f�p��>��E�'�������$o�]��d;4Ri�Kg�9}�+�U������3��EÇM���[$�u�Ɋ6����R�4&���Q�'����Y����E�_��|���y���60��Ē)��GĬ�?�"�H��������s����������C_��%�,5%D�I���ޚ���&��'��\�5 �oUs�Uy�Tƞj��=&�غ������n2j�my8������Q�͵��C�#w����Ә��3#U8op��pK
=���~�S���t�ۙx�K�G�Ӻ�R����u�궲u@ڛ���`Q����i��R"�bg��Fs��'��xʐ?>v�҇�g�4������w���H�:䐕=#����~�C����hd� }���OzJ�M �&4��-�nW�w�Aa�i�H-��!g�H��ù�S�E�)�!���x=�胰��-*�ധ^��A*����{��9�̫�X�=P�*��,�[Z\٤�� ڿ��8�
|�ک�!�4��M��a>;⽍����M>�=]��i��F^�����~ø������v�Gp�brM�B��`T������ݞ�%ϵ�H�uc���j�� �۫\��1ߏ)�d'F��q�evI�th���j�U#m�:mI��'z���[��[3�7c�/��##���7����<����&a�p���zFh�����RS،�Y�\!x�J�� ����f$lq��d�Z]\�fw�$�Z_J!�g#�
�4�;����c�x�>W���y\ǖ�nc��=�b��J������S�a�a�sn��;�6��u�"��ē2�sz:�@��mق�g�H����xi ��}�F���)}�w�h%!{x���m�_U�ѥ�{;�R�ǆ���L�A�M!��Ԟ��kNG��D�����OQ�J�b�9/'��U/�O]ZIf���������y�L����q��1�����6n��+��"�(�� #�6��c��Jg��H�J��se!m���v��z���=�����g�? ���_[���Ie��QC�T������_�bO�+H+QT�Q�=ԓ3�*������e�.^���!�No�B��M����N)��6��p2��Oڈ��P?ī& �]� X�_�eh���� ��tgl�^ConTX��(��v��QHy	4Z���xt,hCOz|(�f��[C �+��8�f�%)��y���="��N��o���%�X�/����┎N�IZ���6�E�+������5��+�Y�����5���߇ $�;Tn�w������ۙ�(��S�"q&N3��������Di���y���� Z��^4ǣ�2IJ��ANw2cXD��_El�Sf%Gy�f�,Ũ#�R��$�傉�?Y씥5����d��w�����c  ���y8���tC��h�2��}$�F�gh"�7H0�Ԝ�Pn�0[�$�<��U���>���LJ�q�����a���yTD}�̼'���pv(� C�U*]൘g��z�T�Z\K�sz�~9�mY3��E��2\��TP�RSʾ���ۣ�-��'��	{���o���̈�yBA�()[q��i���
��	�t/�B@��ltj.q�{Z�k,��u[O�|���0iT?}�
���(���k��{T�b~V���d��L�{��*7���PL�r���O�g������|�VХ�e+aD���u�?0u�g�҉�g]�#�,x��+�A�ӟ��QXr�t�	k0\�q{���x�M��1Fف?��7��A�>M�r�ʎ���	<|��'k�D�m�� _L�[�SDy��4T���9��HG��d$[%^���C�X�����3�ސj�1��tu���j����*��fL�z��a��yN�!0�7�Ff,7]�y�Ef�6е��� MLG)s1#���>���Njz��@��ߤ5k�����u�.&���=w��(���n�̐ SN�K�'P]�@j�vm`@���w[���ݚ��y���8W��ӎ����6��0���S�R�n�5��D�yd��`�M�&�;�ڨ�Aؠ Z��0���V�!�b0�Z(t�F�
�e�%�RO��1rs	�]p9(^��6%(�;�Dan���*i����b�u6ߙe<<(��/lѴ�$�j]K�z��WoC�J<���#p����.��q�Ԫ���Y7?�m�D0�*{���҃��3�l�G|ڍp�0伯SQ���1ظ�1qz���R���ه\�J��v�9&��3�k� ߼�#�i�����gC#�tR,�N�k6[x@�wg�揓�%�%
�v̯���|���o�2D{΍a�ޑA>JO��H����?f02��49�b�/��АR$q�҈�O�_� R�d��|&�~:f�ר+$��q�wDٺ����?�
���z�/7�W�Ԗ)19�2C���!�d\2MH�U3<���1�94���p�V�j�R*���x�c�3��|��+�ɛʿ���m�(2L�����/#��+���E�P﯍!K�E�VD�b����+�����AT��nS|$Hi����
��\&"9�WB��<b�#]�<�_��$�x�na���!�Tt>C�nZ%�"�)Sr�q�<`���r�Mp�Jl��Q7r��8��v1i��'3^W
F�^x�Й٘�j�\2O����?a�q+�V�W�C��v*��cƜ������Qɸ����t�e.�@��Ws!��
C���"F������S�5�K"�M�l���؈�y�g1�Lac~
��Dm�\��2y���]�MW��@���d��B�_����J��X˱`���i)�����(��h���W2����z�x�)�p�Q�3 � ?l��WHǅ��$�g�2�z�[X�|�"�m<��K�;&s����K�g�w���C	�)�Ģ��gk�c��.�0��%���j$#n���o�ѵ�u@���E�&�˼���l�rt�j:0G�<�R��/b8>p8�n���r��UP3�OfSt ��f;晨�A��u��p!�-X���E�N@\z6!�+� -/f��r����#e9&M��7s|�vv٢d���D��tfg"y4������a6t��T9*Z���	m��H��
#��%!,	�x�j`��o2qK�)��6�_,MR���ݓ`vUь"=�3Q,H(0�ag;�PЂXΜ!�7�vu|��i�%�:����b_�)��i��M�D��3��7�����{��mࠩԟo��:�K�dȾ"������|�:M��m�k��6�'L]�����I&M��ØH�;�Ih�縷-�4Ke��j��Y\����o�@]2��,"[�;�
���37h� k�|��L;2�5"�Q��E�5�){��B�l������7Y�:W��P+�
Z�ڍ���=�K�<��c�ѱ��,�����d
o3�8��n�6J#�r�� "���Z��I�ͺ��]
���ʳղ����z�x�d��;�M�1�AȨpmKĄsL9����Q@p�H4�c*0"Ue��I�@LWcMA>!�.��z-^�	����B%���l.q�og�&/��`6�	4�� v��͡�E�������S����jD���/�����&�ih�T�M�vc�L�Nz��Y?���i��P{����8��g��?�.Yr�D�5�i�O}�m߉~�/
��,���d܊D&�q2�j�N����	:�)s��+v����Wb��s��N�'G��.�0!CY�8:�a�Has�^
@w��{���cb�]�c�S�r�4���_�3��f���hz��-|�A�0w�8 ˖��0h�9x)MH��=�mȫ!�y�,4&O�T�-Ռ
]{ݽn��ku����ʜ�K�=���~��?7T݊:	�Nj���6������^^�Fr,��EM�}�M�G�)�Q�S`��_����ӡ��#��o C�����[��ImJ �`}�JSe���Y jcW��
^�Z:��S�mY�]���ȻF���T?<�#�g�}�c7]�+�>6�f��,�$qi�.&��R��|�Žћ$$d^�aP
�qq�[��яę˲�_�5�.'��ц�ux@�܋����O�!"!��&ݬD��{x�t�QXwDC�4����	�h�W:b����'���K��
e�~��s����2@�%�����V�hs��uu8%����B����AX8��~���,��9��{����G�WE�ڨ�c���V�.{C ������r~N�8�볃'���-R����wf�gN�� }^u�+�i�i�:;_�Y�f[LD�	�[����߯��n�����|7τ?�=M����fb��4M�_ ��aTz��N�j�-c�`��D	���6��}�è��<�՚�߄6Z/�����4��%�UP��J�]0{���E؜<�Y� ;�(9JƏ�v��Fχ�����Hӑ(��`9=K�w�]�Wu��U�{���Q��D��hGQDb ��|1�ev���`j�je�+��*��B�R�î���@�����y8c����y+٣���\�[���H+���B�M6��"��}̱U�&����|U����Z�v&j�%	_Qy/ܟ̭N���S:��OK�J��5��c
'�d�,�4/���ڧf���$�t|۔F�*Ų�а�Ag����j'�`R����"����,�<I���6G$c ʵ\Q;_�R���^�j������3�qA��C��r)w�x˒��d�O� c}���X�������b�_
�u 1����w����Q(��轆�Xc�5Q����i�J|�%=����^�u<���s�0�����Q�|�B��$o�UR/$�ՊŠ�����i���ʵ���]w�@�@9�&7����P�h:%I�0Ҭ4_|3B���8��Č�k1�Z���i���r��n�֯F펆�D�S�IR	Bs�8u�<��\�,�0�������Uԭ �~�m�݈:�j�Eh�=H"��V>��bϼc�l����c�m.���?�ѐ���6;�Ȕ�-��}�&��G`R��6�Z�&hWKg1�z��t�i`<:G��3w�ݽ���g)�ϭ�j�}^���N_9����E<Ѣ����a�uNs�HG/�e��;���
�[^���r�<W��|=�ԗn9��h��3�H�e�m_	f�����g�ܫ�!ݖc21����^�J�9�u_���+E�xmS	Ӿj1��Woҙ�}ĺ6`=Ƿ�54�q�z�����@��.Uoxz���xs�uBh���}�N���D3ZU_χ�.!�WM�-<���ݨ/���?YZ
�o�YZ&S�f7������DN*ovwK���b�>%�h!�� �%�I�=>�x�!3l���􄑣�rQ�M�����B�A�H��D��N�$c>����	�VY�K�������h��)��ӓB���E�� O�,��*u�8��O2���A�腜�ٙ{6*��L�b�=1�;�/ã�M��ߨ��t�`��.��>��G���$8��Zx�����?o�
����U��>UQ@]Fu�>�P�k��g-a��Q�ʅ�Cp�O�@�I�d#���7h�����vΌȊ����Z��Xc����XQZ�M��/�<�x�%�#"���Qx����!حѼ���e�]v,���?e+���9a��v2�b.f*4��h/�_���h�_V[7m���w�L�rzgAV�><��k�"~9Vz������MN/l��@>AF�!3�=͢���X\���$/��U?m7��^����fC����ޮ��,�\|�cݨ)Ww��r�$�"-�X�{G.���>�jƨE�$����%wꦚS�&Y�����Z}�<���I���/�Xu6-��?��r���m�4�/�iPB�sر�W�h±F6��E!ʣC����d�k��"��
��?&��,G�zӫ��r� &��/���CT��\(�Թ}A��#v@R��mhߑO�<��迚O�D�2c�U��e�j�(W��g�9����[��\1ɝ�yM�c�$��>����ޅ�2�,�@�O�-�K�4tar�c V�w��A�1�|����<�=+���&�%\���@ 9����mH�M��?�]E����J�.�9�t�"����,M�dT���#���T#q,:��� 1��]X1���^j��{�-�?�_�:-��:��ﯱΎ���m7����7�[���_	��Ѿ�5vF��>��Y�_P7��=ĸ��9�ٝ��-.A{g���FB�e�G��V�A�[t�Qе�\ƍ�^]ݰ�.B��Yك�f��Y������}Aaļ+�Zq۹:hT��"~�����֮?��i��&k�\37𕻐��5���-��l�j�c�"&��_i��zE �Ǥ�rc��`]�~�]�K��8P=�WSwg9s�3���M��smkF֒u���#w�B�L��T:Կ�	ޗ�����B���3�$/�s��T���4��	_�[a���jh@��EK��b[4�{���2��$��8
c��z��E9���f����dL�	M�l*�T��.X�ƴ������KH�s�W����!=�S�4]�i�ӊD"#�M��x@;�XGb)8�^�g1&�w5��đ��Fk�Le���5�|rC�6�ÎP���B�2_�籏��Ǹ|Q���stj��Bb�8l�z���7��������.�c,��x�!b����0w^��10\$Pcr�%�@��1��:C�2=�q~��.�g�W|�X.�6N�>l�p%ZL5�2/ؒZJloZ^p��L�� ;��xeI~��,e;�o���v�O�y���㉉�7d������h�l+�r��t��Vr6��Ϟ���c����M����mJ!�.;ԏ��k�4�5��:��j�Z[�V�<6���M�N��݈�f����^�&�;B6s���/�e�SC��5EUaU���|�R�~=��tC;����������qx���3Yx�c-��7��O�UV��r����n�4@��!`(��S���a�f}�3�@�����\���M��7@��Q�ݙ�R����H�R8�l�c��OQ�� ���A ��!������^B���������U�T��ߗF@CIc���
�����s��_;t�v6��*=��m�b��9�xݝ�UuRr�L�2��9�����lq�+����XA*S�����qz�Z;��ܤ�X���xd������Q#�C�3U��<Xn�tE i=�+��a�8�Y�/O����*�O�K����2I����KC�`��'9
?�1gV6�<t�4WÖb	Q�B����*o�q�9������`P���m�p7-���wq�%Q��� Ro���"�T�%�П8�/c�A�2v�dO��>��Q.�rUx�yKaL�*��j�6i�k�Ľ�D���*�(PG�JQŴ�r��*Y�SP�V���t�krTzbe��Z�gWx���b*Yu:�?4-LGsT��k>?�9�AKo2�����R$l��a>�r���qjj�ʻ��C��a�	�_rW@�3����NN�Gm��
�`�Ȋ��q�*(Z�x5j(��l����:��h[�L �=.&uwY�1���k��N�>���p68
�Hs�9�ڍ���N�#��m8��LƁ�w��"�����+�4@<d��o��5�9�<h�.NҎZ�RȖϗ���qQ�3q{��3D,�\@}
=*�L����Z��U� )L��G5�SS�tRVa���W��X�u��v���}Q{��kf�X����R�M'<Z	��T�z�eZNpw��Ų��<zx��>��U�3b?�i�-����V�٩٩]����j�K�f�+��i�!�I���kՆOݒ[���\�����N=�� (�CZL���ye����A*:f3��ko䙟zW9B��"ͱ}�S��i�� �,���4t�ǆ 'v2�"@��/�]�7E8���u��h�W���c�TL�/U�HKܲ�5ɷ�jy��1��d$�D�`�B�A^���P�f��<$��()�^]y�G� ��p/'\
>� PR�Sjo�\��B7���+�_h������~T�\@��R>Sz_Ꮷ��(.eR������.4ƛ�Tcq�w���䈋��E�����O��X(;��~��|I�@C$�8Wb~��W�v�j�ϯ��������z�.mVe�{aL���*FX y� U��(��(vh���Q���g�/�ށ��v%|(�&l���	�mK�Q���_�5+��"�e������M"��"����a!P��c!�T3`���4��W��)�����!l��$�I�*��)��,�W�xg�l��r�Z�Vh��c��6hK���%�E�
�h��&g^���bιp��Ж���><�Z2Cv�ߏ��~o��q�>-,�6ם�h�7����e�F����Pv��G{^�gS>8?�<!T�W|���	�}���*�$޶{�g�@�njݛd�m[��- �;;O
���l9�Y����Gg�?�Y�� ���jd[���O������w���T���P�����7$m�0E�H�y��f��
��#�Og�7#_8�D����E\5iL�y�ط^ӝ{�`s�-���4W��Ѧ���N �^��Vf�T��7vLŞ���5���3�OT��A������T����g�0[�!+��zρ�lp��0�k�㖋k���I?�Ⱥ�l���vJ˅�����xds����,v�}��r�j�0��*fT��&>��ز~��i�6=\lUt���e �C�}p+Ք�A��['��ZP4H��y�[Z�@@��M�SW��ۘP 2p�r����'�?$�~`�k#�-2�cL�P�M[�-��s<Gk������p���>a�C�ɾ�����g�O#W0Z�\m�:�@Þ8ӹ�C���L��6�n��V���o6�|��.��Z�	3��Y4B����b�!�l�*������z��=�gw�.yFZV�?ot��ʽg�9,r_�|EQDn����H=)y4�TN�G���˃�к�}��!`BB˟8I�hg�'���.Ix��T�x���R�(��'F�[%ŏ�h`;��r�ӵx:A�Z\�,RÈ7���F��b��ǻ���^��¹����8�~p���.��6�-|�Gr���d��۸<�Mp�	���iSѦ���mA��{���9����rc���v�hg��o;�}�7���4���ڢ�Y<;y��՚��jkR��Eܞ�����3 U*�4�<D�����Q$����s��ՙ̤l���W�p���K�R�c��D�7��;)ªz��`p4��`�l.�܏aE�WQ�\q��\�ߎ��*{�Y�g!��Cڟ�F�,�=�����j�1B$M�D��.�'|��R�B�S ���4��H{lB1dSJ�dJ,B��ʱ� \�˅;���l�cR��exe��W�8`>���Z��z��W�v)�����̡;0��X��{�8��x��_�63J`[(m��-�(��ˀR��_�Yt?�Vy�#mr��sJۡG#���j�GX���vӥ#��/�Ӏh7�'oV��C��U�����by�(�J���@���ԏ>� D3"q/h�0����-�����҈�˚F�nMqfj��|[���Ӣ�K�x���^T(��U��zU�ʛ,��.bq�S���[��Cqx�� �^ɿ�����Ϥ��� ��lI-qh_�[`VI<qJԥ���c?��B �i|�%�ye�ۉ�{�*��4V���g�2���J��5.r�(!��z�ə��e�Ʉ2�F4�O^��7L҈�.:-��#>Km����M.vݎ�A�-��:�����J�]Tk������R`�	VQ���N3��������YU���:��h�	�~*#h����կ	�z2?���M̀S��>���H���n�L�������,��O������y=�����AC+U��1n�O%��C��M��sX�Q�pbp��PoP�`�Z��1{NY2��
�HH��}!k�r�y[��I��� n��U�e��L��f����[�_S�ꔤ�܅�Ӷ��Q�D1q&ŗ7�iDd�x-�%P�I��yQ>q�Ø����(�ϔ1)'��bТQ*���ؾLxqq��MB������[4�9�_����7��]z������"w�n?o \� �y,b��X�x���� S�#p�v5�7�o*o(:.�<�,"v+CD^��h[�3m���,X���?�8!�}xJ%��J~��i�!�,!�<�w��#pW�l�7	`Jc�S��T�u%L>?�z�F֙?�P2n
�P�Л5|�y��ڱu�-yi�X���'嫟����x�D��"�+G*�yZ(=&D]���YD���t�a��0�=�����ؿ%~�B�`LQ+��{���{�i�b�[�/-�z� �]�#*��v�����C7�,� )q��E�XΟC^��PNGA�[=��r&d�yVz#���Jq�\cD�w�Q ��E��(��l�$5Bd3�}��5	dv(Y�p*M ��:����A�D�R��������9!#`�-V񬵃D��p���`MZ�86u�
����	gc>܂:���n:|�ｯ�u�S\�v��Dɉ�]y2e�q�Yc;��0�bJ��..>)�1��R�%�*�o��tPQ[֎l0�����hy��8�$+~�T��q�<p�=�]��,I����c�`��ժ�����������'r۠��x�)ٙ%t��\H���%�#/<#���V�h��N[v�Ӭ�� ��	�zCh�{��jWQC�9k�6�z��X/���w\F֋��T(泄@�cYz�+�����{� u��4��'���&�mg�"����1;�����;(���"��!?�]s����T��]�T������o<�,1�#O��5�	js�j�?���{̬�.�7Ю).2��L�bXWW���<2�_,�~�S�2�N<�TF�g����ӣo�:�nÑ�z1���0�Y�^��G���e��t�ol2�>\毳S6K32=��cQ�v�D���ؒ�lĶ�&�N�L׋�B�E�#���� r�ͥ<��'`I����1�Ҟ�'c�'�BXxu�=�%��W���W
#Ր*_��f���":����75����vgګC<�Z���GRi�^7aO�+%��%��#�,����7có*j��TY�t��(Ņ��f�(�O}p�i64h�|\=�^ʺ��ˁ�,}(��S�O�=�0A�c���;��b�p���j^z� RG�ߗ;�����j׊Ed�=��B���ˌyO�.e*4#��&�K��N�(����(�3�+U� ]�Ԫ�h�Nz���9��i���o�T?���.�,�&j���G~VE#Փ� E��͠�75�e�mk%���$��Q�ဵU|��Ќ%U�X�&x��2�ڇ�
 ��6p��C:S�$\B�N� 	<6u*���q�T�1P��f:ϵr�ă	���ω��d����35����8�ۘ�C�H~N�ё��ڸp>�*�O.q!J�CaC\�� �F�S�iJ���BW���S_$ 
 t[��N��es�������#{�h]ת�U�"��T��B��Q� �X;g�u�_ژI�x�I�L��CO#�P���oU$břO
��FZ����2�� t��4��3��\�b�UpE�P ��c�w8�5*V��6��(�5f����%^d>���L�@d_V�a�B��0�� J�Z%%2<�Fv��ߗ��9(�c$�~���z� ����j";i��:a�̈�
���J�$E��L��1���z����e�G{	�9�J�ߏxU�QQ�t��ׁ�|����yF22U�,��X�T�&mkT�U�R[��VJVG-î���Q�*���x>�.1"x4�\���'\7��X?	ں�	"n�
�C�w���2',��b�7��7�@k�$�~t?H��v!Jh���?Dk�bZꛣ�]��u�cR�tؖ�僣O����p�}E��	�7����-�N
*��������Ȕ��W����E>�i-�m�d��w{t*�E_�厬+��Uuֵ�9��!�pa��*����GT'�G�>~�wZ�E	�<p����v$�\��Yd=՝8- |:;N!Rx�K�Lw&A��L�{�p՟-,�=W�}M�� �������˧A�L�:t�j��2���$W߭��-�����O~�܎��V��J�͗�|_ǣ����	���2�Zd���kw���s�V!����8"�G[;~��`�A �+�'�!>��J
�e������@�{����H%�xh$����E=���>��� �����
��[
Y��hF�ف'r�D�V�ν�XU6����B%���Y���u�Uʧ1;{/Z�⣵��cj�P�ϯ�'|{3���A�����Cd7kQk�a��T�9sB�"�K�5���v�z���X%;A�"��M69!}#�#�Li�"��r<6�Vq2��o��_ |����@ �������/�Tl�p��>�	��:�x�1����$d[�<�����9�	F7�����.�|4���p�B��2:�7l��K���M�����X��ԉ,����vݾ��(s���UV���q�(�=�D^Ck�b���˗zK��Bu��*��@WV��cf�L���	h~=��8��������T˛;_n�(���g�a���d�2�c�R�%�
~f����)!�VN��w��z��ܕ���fN1TKQ��y�B6r�¢�jg7��rq'�wyA��!�;T@\n��w1��s�����$��/!U_���z�+����oQ���N�&ލ��^*�EU�SKn�Hw)�H���sod�0��nQ�IR8�-��Y�EF���V�#�M.\�
F�B���?D?�1j��\9��)N� �j ��D�NwLSL?{�q��#�E��=P��2���('�� �(/�4��r�&2|R�H�*��:b�p��N�y�kY>x/C��(RM�$��D�.z��fÆA��ŢlE谛�&�Q8�l��[�Se���g/K�F�/�@#(,�a%W�&��t�;]Z�2�e�]#��lR�&6{§�4Q�M�[M�5N��R�8��j��׏T�:�:4�3�W�J��u�V6qDOB�_Ne���F�����*-�x�uI�q_��3��z����ݿsm��9�Z�S/�7f�v��'F1�q�`e��;BB�`&�&cT	��g|�	;[/�aN�TZ��
�yF�'��\ �X9[����k����|z�{�� �G���'�L�^�6�y7�}�B�X
t����l&�Br�c1]1�S�)p�k����4m�e���v&�
�t�*;��8ؐ��`ڇ��T�,��/���<dpttSI��w�Ӗuo�io\���<rf�^LC�z���f���X�3��%�VsZ�8`�I�$��ف������©��E��x ���!L�ݿ�Vs&�����|_U��w���c�xU��7��|\����"��z�N�X�v�a���1���S�7<���k�	jb=��X��ƍ�#�K��0s�4lűw�XW;}_}|C��E�-�\�#���ax=
t!�V��i�����D��Ը�ݝ�+/�6�L��< ;��b�1����_n�Z�ѕQ�RG����̕J��sg;D"�h�������u���~k�.n� 	*MU��ݻ-)��PI#��q�^��7���d����]3"���fʂ�`:�/�q�=�D�̬���0�2��rL�.齅���yI`l�}߼�۴�24��>ϓLr��?t������W*ܩ(������W-��m���<���3��Qp���usEK�D��_��t�&����bc��k~�CE�6��pi��Il� F$�F
#W���^Z���H	���L��Y�p� Ի�`�+�y�j��a=�$'���^�S����Dv(�'�Kф��|r[�ee�*��|�G����K>Ӵ��'���@���]f�R:��8�$G�ܨ5-�Z�&`^��c䎱"��F?��L	kw�|�ϧρX�2n�;ۇ���k�H��j�����"W����q�r����Ε�rN1Q�1!�A\�n�ٖ��m���V�v�e>���]y�Ig����!�X:�(�X@ؓu���',���,�W�g?j�Ű7+P����ř�lp�1��X%TG*�j��[��-����%*@j�y���-��6&9;p���ɗ��q�W�s2s�O�A�.3����	�M��<qE��Y��u�B�8�(1�y�����6��]; �jY�ԓM˿s�Bd ���ذV��?'����~Lg��RX�?	u͇� &<7}9u�5�0\o]�z�A&7���mq��fL��Ē�tr��oc��00�K	��鬕��^+�9׼iE̍���Y*�7|����GQk���������Â�x+e��a�z�j��;-�z���$�4v�i��]�1�قK=��)ms��k�C��-/NY��k�EwB�۱y�]	�|�"���j뗙� �Ta����l�q;4�E*5Q��5��6�fKْ�nf�S*�w��.i�		e$��]*i[Z�U�$R��'S�΄-s>���8����I$3.o��n4�W��A��sg��TWA۶X���B�a1oR�ɌN�*�+�L�h�TI��VSJ��mx�G��:�H�q��/cUjM��0�� �Mֳ���MC���/���	��d�`��v_}��aQu�S��c�����d.�p�s+h��im����J�3Ik���1t��􆚡�>*n��y�Z>'�B��*ڟ�z��Gi�0����
7�+`��9��.Mi~�V�M���W�MG^S�c|�EP#,GD��0~�ĕ⻿U�ͨWM�7�[�EPs����W`�r��	�=:c��0m��UW�R�:Ff�E�v���h���a���ܟ���d��#p���2�Ï��;�M�~:�_>��9~�G�< ��βq����&qͰkOAJѪ1=�ދ��|z�vB���5WH��ǠG�H3Ѻ�u������T���Z��?M���-�XHt���P���R'�s�M���`i{���������&��q>��L	�VS��>�}���1���3|�f!�H~�gMP�IY��@f�_}8)��>���DÝqd(~;����RZ��!�q��n�@-�P�{׭��@�?i�]]�b ��Ϟ#�q����vLֈl�g��䣋��� 4�O�����n��#v�\���[SY���y�י����!���U��*#8rZ�P��F�EZQ@�A� �ȹ�L����6��r�b�:�� �����p���aA��T������kn�b�Ҷp,c�zs�Sgh�X'�ޡ��j�dN��ު����i�&�|S���o�ab)�@�>�|�^H��-�Lɘ����1����;�0��_t��HV��"�g��]bh�� ��U�Q�T�s���{��:]�����e�2>�!&k�N�>�0�S3��iÁqXƶ�"����f��$:t��j�a��Ȕ�]%!�M�U%��c�j�oj�X�Pݗ��6c��L��Y�W%���YH�=�ش;�ŉ0��$���#�&�"����ں�Yh���q� rD�Rbs�.�w��m&m��|�C͈����֣�PiE)�^)'� 0�Gq1aH���U]����Z��N:�p��S�m`HDK����=�R�D9�ᾠZ��`�_g�:��4�ڛ,�?��<U�E*!��CI���\���r�%i�cW$;��m�t�Z.�벧4܍�V��5�ܗ���P8�&yCJ�{��̦إ��C�B5BR7��ƣ�`{����{q-��5��d���W,������)���g�+�\���ՠ��ea����1��T�(���Gl$C�K�&��x,g
}�oS�ʲZN�	.,���Aa��t���Y�մ���7�1n3Z�Khr�F��o�:���]�Ŧ�,�/�#�ľ�����x6}~V��=[L��%�b���Y���2/]�������֢��Z�.�Sޠ�s��c�V$L"�3���}X�u�2�9$b���D���	��m���GlW�;ÿO��c�9��j���6�rԲx>b:E6��1{�3h{@���7B?�,?�)��|j>ף��G����g�h'j�Ũ��g/9���9*Z��Ӄ8�,f�K�r����auD�ڸ�с����g'خ(Q���H���vl8x�X�q@��<#�H�%��.3(|��������_�&��v�y��a{c���+��{�d�
�~�TE6w����ҡ�`��i�Qu��gM��=��	)�������D�K������i��gIehq�� (n�!G�i��d
#V"�dg�� �lQA"�8�5�l�`�QZݗB$�/.�"n��C���l�%I�ㅢ�i�.��d��ǐ��EP���b9��֤�a������G^�����ؐ5���G���h���m%�e|M��L�ײf	Àd��S���6������~;���Ðz �k��I�־��y�;�wF���*�#��$���6RV.��O��Է�P�s6����h��px�A�uO�St cB�z�p�qt-J�Bx7�4"Zg1}���sA�+V�-km������kT�����)$D��	���i��z#�5��s�, �w��p�p��QW�Dx������/r��G�c{ � c�C#zV� �X^|�IOU/�̤]��	$�[)����k�V����p ��#r��c�;�zw�#D|�?�6�J�������{�=)s"�	pq=�$�U�k0*�,��h�S���dt�{�8{6�I�|���f̻�����R���X��͏r����n�q�-��	<�Q�J��.ݩW��%z�/�"��md�+B�pB��d}�m��f#�l��&�����<ɸy%���c�k�F���O��F���7�b&�w��UɏH9l�X��?�� ]�]M�m��*9>�F��@�w�r�.�9�C�h�/��[��>d[;+/&^�<��_�h��%֨7��ǺJ�uA�CTb�ۡj��x��}�.S�U��Mm�l��A�Y����,�?��o	�N?���0��෠��i�響7�'��=ݓ-sa����:3�K��{xQ
D��"�KieQ�L�����B��ޏoċ��HE� ����<$�+�W����������
�2ϧ�O��"�s�_\{l}��̡��KZ`�o��a�8(sg9��VR�1����^�_�P���jRb����
��Y�7]�+L��bC�α � �(=<\��tU`L�������1�}��p��I(n*vd�`�x�uq�T	3�P��(�ⰿ��P��(�p�jċ@�"���$��b�v}�d�5�����_D�w�T��_1Sη�ف�r;=�=<��afm��m��
8���b&��]�LF�UqIx7��Yg.�W� Bv�v��i�����d@D���w��<�2I��\ ry�ج�z6V�C5*�>�/'so��(n���R�]RVJr?`���wt�{�d^Hn���[J/n��ʑ\�f����3�q�//���Dt��V�z$�ͳݒ��E�,�f��M�t�Q#]�Z�c�A�K�Q��@0G�\~���T!1�\{gjhd̞�,�ɻ
��Nҥ����O��C�����@e�N{��"�ɷ� �a%�uPvA�+����䩾2�����'�K�Lrz�+�#H|W�NJ�����S����'w��F�czSB����7���\{�����)|s�*�z��f�;�w��	���Kv�Ґ���>�����cIJT<{0���c��N̅����|��\\5I2��n�^11?�'�h�������Vw��u�D��C����Z]d�'�sXK�|@h�mH,��_"�����Z�nO�������6���c���ɟ?H�A��~p.Oǫסq��ëd�����&8t��&��3���Gƨ��,���.�41��+j4큨ϟ�3��`���Z�
f�{x'a
�����ǧ)v���aq�Lpk9�O��}A6�k����{j_{.z��R(�ML{�4��Q;�؈�#��r�v��v�"m��O���{���-�e��w^Q������s����;\�ʺ*�%t��>�x<���H~���[��E���(4@��?,�v�:_��ɩ6԰���Si����	�hd�wg��C�I���.K�y���bg���'`:�u�q?�wd)��Եcw��b(���j}�=�S�����/�hIl��˚<��w�p�X]%��P�M
a�	".�Y�R�A�@PL�s=��^+��5#o�g�F�t�=@K
_���"�������ou
���:��R�;r�`�a_���{s���E"�L�l������pG�_HѰ��`���`ޕ1��a58I�!�	3�Ƽ_��A����.<2vF76����ђ��\���qhrFP��H�Iv�ࠤ�����RmP�J�ձ��>�ᖅ�U�aLL��~�KgK���4�|#7�U��zS���ê�_��B�Ÿ��<6�Cj�,d_�by��Oe�=����
�t, f����P]�q�x��X5���&������/�l�)9�{PQ�	�y]����t��e7���H�^W�F��$�*�n�H�|��p�?��;��zO�c�9j�����%Ĺ��s���Nj�.���z���Jee	�H7��u��n�P5FW��\���6%ض �w>��"S�-�̿�Vi�_��|>�%P�݅槄N+��)�t���Y�{�~B��1l���~�>9e�TU�"4���1�)2�Wz$y�cΑU���LQ���8��Q�AY�/3	f�|�Xʏ�E�Z�%8&xSl���A6:��dc��ӣ*�Ǳo�%[*:)�7���f�����Z�8X�s�*5{wj���V�b�?|a��`yY�`u��C_�L��K��`�Ua�P���d��{!=��텰����ER�-��ЀAE���0y�:�n�@�\tS|�-H)�u5�8�@��	�-���4��x?�t����}	3M����5��)y�4+��$��z�ͣ�=a!����b�|W`��^�j	��N`9�m^�@�+)��E����d	7SBQ��ǉW��$]��4)+���� �?���=���5;�_H!!c�}9���2�ȃ#���2G�"�g��E#?��yd�i
�����/U�犽�7^�����6tf�愎O��v��s(R��L�,�v��%�ø���C����4y�����CeK��Ä�&T��v���q�����(rM��dl�Y����YZ)��o:-�)La�V���7�wK��i��+V����ɶwK�+�<��+<����TO�k�D Gd`��w����(���3��h:Ik6q��C�~���=H3��l�-Af�c�]B�^�+=��M	u�W<-����;6>&�:�t�L���A�$�վd ��Dn�G��`
�]�����X�:�D����֩z�_�y.��p��m��ruj����&��X�����N����㋧�\��f��jZ��O���.3m���vYx�o�T3M�M�d�?�O��{�Z����j#If�$-�J�*�� ru�BFC�G�4��s��Ȓa{S�� UY��e$��l£4�����3X�d�&���=_��"Ǌ0�/?�a,��ٚW#WMy�j��"M�&�W�K�z��t���xðl,=���G�I���'��,�S�Nםk$d_�Ώ	a�yo�C1��_[�o9(���[�{�-�|�&�8��� �>Z�'��nО����US�	�s-I��]_ʀKz��M�q��j^�:�c���B���ۯdK} ����[�!IA�kl#�h���\ҿ�;	=����3�D�l�Z �?�F�x����.��!�����L�2ٿiA�|pu/�0aV�����&C�qYNK�y��(2폌*kq>��Q�0"�+�#`�Z~��.y�%�wX��톀ݷyj��{�P�3o���Hp�|��i�w���G����S��,���HBW���	�S�f�+�K��@���P�lW����^��	�k����42���u��[����`�뫊u�RPw�Q������J;;��nwǧ����x"�؟�qSnX�i%;V�%�T,%��&��Wz�UQ�k� �"�f9�p���ѷ@�����"�'-���yM)�Z~2K��(3�v#�H�C)L������� [�.Ń��|EAH�pιO	��`	@�^t@kq�{���}�wkx �6�R2{x�s���2_���}�ی*���7>KbD\�pz��ё�F�Ԩ��u`JE����[��:����K�R�����{�#�)3Cs�,hq�|}y��+zէ�m9��B{��u�z��#Ǿ���I�6��(�VdgSm��)W�Bt�Z3���\�F�A �w����y�q-�]�'���q
ҪQW#8X>��
�;+��㸷�0~�c��hGb��)����J �4������t���wC�N�������yd
�;+Wo>�(p����x�.�&���E`*8�8Aj�<6�a����{�܇G�:\�	R{�������M����J��)/�o�f�?�����a%3x���N��k���t�fte�q�`c�z�� ����1� �9��Ӓ�n	�����V��u�������,::���l_�W/Ms+�2"����Z���R| �aۂ0�G�J������I��h�Dʡ<}�t�3a��]l� �����4rM�����
���;)T����۱�y8&q�u�2�\��b�n�SG~�*��l�~n��-�CS@c��2�
<7��=nl�sG ]�j;!�jI�"�����Ni�yq$]�^g}c��Af@`!ga�*�f�&���lՙ�����Z����N����ؒ�ʨ̄*?H��te���&Ty���Pnv���Y�ގ"k̫p:�z�~R�{pq_j��*�3�b<I�)'���K����}�SG���`��.�5w>�߆����i�ں$���8Ʃn�53))�j�X��eע��.tj��2�G>˵n��,^�-Y,����TrTU�,:��_S@bD��O�4��M��yMxq+��N0����|��ǳv,ގFg���j$ub+z�s$*� �f���f����u�*�y:����"���?'ڼ(W<�(*X�%M#��Zß�}a�>���a�Ydh��g�+��s|@��~{�z @��k�{��t�9k~���qg�5��o�/r�>RԺ���=b��^���@�E
����ѓs�~��,��6�,��y�~�5��]yA@�þI~i�NAA�A�`��X���16n�r�{���W�o$�LEn}|"�H�u�n!z�}�8lA���ؤD�'��b��ĺ�"�(`8�jE'�V���$��k�ǥ��UIǱ�'E�{lԡ�6�}u#�B�ʇ_�IWd�X�/^0Q�.l�^����s����6�ݧ!�)+��6J����\���v}��b�Ɔ,���5_j�����O���D�&z9��� 0r+��\H��u	f�����L�@TIW6����2�@,!���WyR
��W��`)�޳Y�:�r��+H�r\.���8��2�l<'1U溦�w��"�0�t����0Y���S üM��"U���.ό
o����K`�?e�uE'�+�ܦ���{��R�ET?X�'�2�97�LfV�(�-��"�7iQ3>zT��ZOO���l�����&����n��ۨCJ�2�Wg����s����V�gAIO��~3`���^I�9 H������_	���G=�H?M+�	�gT�Ya��d��+E�����5�����׶�k�p��_X�b�������S�R��,�}�}�^e� �3�;'op��u���r�tQ�l�b`��5�e):;��֤�*� ������I�k^1r���� /��1Ҳ<LcE�Ts�2�i��z�ɺS-�PY
>+>:l���4��&��LՑ�ow� ʗF�F5�ReT�G��z{��hض����u� J�Z��W�x�j��8J�bʖ	����P%		~ɺ#y=�Z2:7�����h�F^�P�T�ȹ�Dd��2㬦P367jg��P�ඈϧ�"U���o߹)C�%V�]�s؝�5���[��6Dux��$��9��c��N-`���{��eIR(�-B/d�w��⪒e�	{�0�p���_/���4�#�ڟ9It�`���i�c���s��4�O��y�1�#"L�蛢|�ˢ䏿ǱL�"��@	|�t��F�;�S��:�9��nH!�Q�]�>6���*[looH��Exw`l&�}�n�)	��0�Fv�o��D��8i��B ��ops����d[I��	�Y��!P�|�fe�y�r�#��+�F��<������ߢ��t7N4tL�i�)Ʉ���jQ���Z�j3��8q{�*��[9�r���l�9H ������p�Ԥ�-7SD��U�c.�14��P(�=A�$��o��4]� ��� lv�u�L#�ݓ��t�2j7�)Y	���U��E�����$��
A.����v��I3����V��5�JA�Y��%V�oJ(�N���!��Xo�;�E�,�����rM�Z�Q3�jr/�fD�-�)CU�+`Ʌe�|��V,X�0�+�Zi�;p\0T��fA?���W?mmW�Y��tv�������d�R�ve
�,xAͿ��@
���<��dZO�U��j���R$�Ĳe���I����ؙs�,����,���I��;��$�&M�<S�#�Ph������l&� m��qmL�E
�m{�G����z��T��p9�u`q�_z�����> ���Q�u�]�O�pb`y�{%��GpQ���!�g⼽�(�:11�;K�F8�(
�A2�Rԓ!�w�ӉK�[��z�}����6|j�%'��S30�(��!���^���p�HV�u/�����6Ֆ\>h;ﵵ��P�E7�ܳ�5ʯ,��� >�5V2�k~����*[�t�;t��W]���R�����َ�`ŝ\K�W@5�I��$����v�Ȏ9e���]���S�/��c[�{�FÎ�1�lJ�.eG.ОҒ�=�yJB��(=�p�O9ŝ>�������>�U��鬽{�NP���;��Hz5`�����C���m�B�,���l�o����E�	I�v�������7�	�)P���<lw�Gg+1�z�E�q��v\��sVTP3 ��i�8��yKi=���\ ���Q4_�66�;����FI��s�ǖ��gb� ���Kq���l<Pf��M�#��A�sG�!����$�R^���>�[;�$���֟yئ(��gv7ɏuT�a7�w�/�<�OJ��4ˉ9=ף�"_����k^Kw̑"��)A�.kP-��fw��"����l���T蕯 n�;�F�D����`�`J�JrO"`,ً���!���,�Ѡw~S�qbc�9�lG�
dU��L|�_�8)�>0ܹ�c�i+ā��l}�1fy�R�cŞ~C�q�g�J�-�nFI�A�G!>}ȯ��Df.s^�DO1�h�[�3���d�=�iUD��s$�N��O��͛���ĵh�r�Ap�C���s�1n�ʨ�w&0�l�2�l4�;%�u��a��'�F�qՅʏ�YK]W��[¢�w�A�����������{�"HBQj�8!k8�"��Np����u�}qVB� �+���1k�� 	!Z��O5k?�!6QxM�8�{��"�h%�q����/�ay:'n������G���2_4��1'*i��y�D�&9���&-2WfY~ ��|	c�(9ub:�
���֞�J�i��S�r�Ln�0#��� �0���{Nc�F ��܋��3�;=<#M��,��rĶU�@V_e&�ڷN����w����硷��)�����0Lp� rɇ7�3!�O�m3�ˇM��8�Ls�vݎ2�w�)�ҕ�����~~�4�-����$.>��Yܿ�v�z*"�۾�he��ã-mV�6�	;���k�'�����4�@{	'��`��*L�1\}��~{�@��������L���7~�Q~��-��=sJ�^��U܍�Xd�����M�����RKsS:d�<4��!��S}��nB1O��L��郵u	� ��&��W�)�	�E-�>��/ݹ�=��qۇ�3�����p���"����J�%����]�͜j��ob�X���%����>_.��<��� ns���jo>��P�w����{���r`�����)���W:����7�L�~x���T/]��_jHw+�a�$��9e���{S�&��#!�����!���Jr�92�-�x��������5)?8k��6{�l��ǁ�D�����zw!��L���%�+��cgb��-n�p��Q v��ZX����8�U⤣��@�t��e��d�~���� ��k���ȗ����?Y���u��UA�Ã5�C�pն��]�T;�Q�0p�۵�F.��Ͻ����E��'�n��?�e�<���L/tN�&�/�	����ݗ��.:K����||��Q8Q��IDCپ����11g�P���Ofc=���X��v���ŘP��Qh�p9q2�ꪢ@�)�G�rl����J�S���S�iArI~���
��B�P\�3T�8{�6Q3ϥ�z�� �>�w`�ڣ�{>�1�R��%�������5K�q��?��Sv�Z��+����Zx�܈�ҍ2n����P p�ݣ�62�9)o3m�)��V�	<�j�3@z��ʔ����l������N��+�x�b�)�~@^�����O�7(G�I]���%���B~��Ln��[m&�����q���y��������egW_>�Q�(���{L�!K�!�7���A�	GJ���c��`���@<��.
�0'�L�R�o;�\m��*��S:��t���&^�J��[)�}0,���rcq��Ō�R��)�{k���D"��I��:���QA:�EM����(i�3�-S{��T�l�D1ژ��G_N���� ,*P��s�]Fbu�S�r��եꍧ�j-�_Q0��Τ�&�A��Y��^No?G�R"iĈ��A�������#�����W%�-HO�V�{_5�.�eO3����Η�n��w��Y��7�I�t�ra�uF>���� {��%��e�!}hP�����[���~cv�ݯ�낪w�q3�ї9�	���� �𧇱T�b�?����f�&��C������=.ȑ-�o�-���>�Pgea� ����vL������O������Yh'���Ek�Ǉ��w̗$���j�A�K���aQK?�W{�6�sc����D�(9$�wBQ:�S�ۉ^�ڳ�M<�@�q����9'�������ʣ!���	�Dz�@�����}��$㔩l۴�9� h��u�r��1�p�Dy�b�&��m������iQQ=:��)A���S��v>P]=������kS���]5*����C��Jv��������)}���_f$��eJ�nѺ�D4����9E��NXV\�9|=�r���Ԯ�4=�z�����XEN����.0Z=���=�k�����:)!�c�1b�h��&��1I������4)��6�&o�Ѯ�K�~���Ս�֐k�~uP���%�}���X�
��'��v��Q#�W&�7m�v�-�[���/�Bh�>8T�v���&��A`H�͋�^�J~唎�%��CV�o0�x懟�5���0�ĄM�'RVðD�sN�2���Ýjr�	U`��,�b�T5^p�I�rE�lyuyR�4�DR�o�R5�_��X�uDMA��{ax7((������@�,p��iٲ��Q;S�č�`�ţn7��p��<�i�inԜo�Ȇ�|�a9�79����S���,5���T�C1���`ZoS���I�+�N
(�M�)Ʌ�9V�w�U&C�f^��u��ch��n+��8a[攝�̊�+�t$.���;�#� �[���	|X�L/�R�]2���^����1�0ٱ
�p��঳J��&�).��ܝ�yz���{ ��"��o�����v�&ݮz�s��۸��d�T F"2�|�P��nV�٣w�����Z��:e�d�J3B>�k��ź	�H�7/�Uj�+�������b"�R�v����'5�k  h�J�{-��3
Y��_@��k��7��ւ��x7Q���sG�PK@==O��j�[�`�+r��A����4�[�r��
��\j���jm&.��hEĀT6Qb0͆��N~�=���e,%_�-��x⹏%}�$,|�ن��*���C���+*��G{�QS-�'�\2jB�9�y]���zDJkN�v���ў�˦���d}��fg�<�3���u�@;�qПPKQA����TM�b�]P��<�>��9�$��hh�!'�n�l�(j�f�z�ƭ��fV
��mA��ӡ�S��BPh��R&b�
�-�����U�u�70@���6)��P���^A.���yQ�L�}-�q�p8mZ4B���`�e�#�~��L�j�#V|'���wPL�4�C�~�����,Yl�:l˰Z߻���� ��dT/�U	X+�+�:�	]��$g��W4�5H`Yv�:��j��ԋY*�ah�+�:g��S)Ms��8~U�	's�(İC�s�e/PE��� L��SdU�
���KVw�~�? ŏol66\_u/�) yhe�t��n�m< �T�E�p[i�����lU	,N|�<�	���ͻ	���P����5�l]$��wO<ď����p��٧բ�ՙ��b��ˠT	��i�����#����t'iwz�l萓��|D@��Fs�lCv{]H-*>�_�#7eT�&z&џ��{D;��Wyf�K�B�[5�
W�u�K�t����|��!�']쨁A/*Ӳ���[�1�
��f"�O]��K�h� ���
Q�LGȻD$�o2�L�9��t��-F\K�"7�/��?���T+Ř"@ܬw�� �i�?����p��</:��l��+q������Z�.A�hS�#�g{	H�u�<���������ս ^L۞����POVn��֛28�ڑ�����-���>!���+��M�����4C�_Ot���	w�c�a<K'4ߝ���^�%�U9�Ñ���u,����t�6�K�&ݫ�cs�Xl!1X��q���X)I4�L��Y,���r�%~H/j[�&�t��#9����n�T3��5e�j>R$��Oi�C1�9�a,����Db�O�㞨�yNk(0\b=������ێ*����:�;1��0��S�U?�_vE\��`l���1�8��I���E�w-��sW`�Ҍyl ��4���=�i�J =�۞T碒 �Խ�E�Z�=�Fm�����e�$����m��R�6��|� �!N���yzi	^�I�K1�P�O�R��0�l��{<8&Y�o�g�\�ީfD�����FPx�+C��y���.���N�&�/�}K��l�pWXp�ghk���ay�y_2K=�S�>�,+�JB/�<���~��5{5�[]>��5�G%��Ju�h��E�2y� �iŤ13`�ƣuC��g,ے��V�=bYd�/?�˶�z=,
�-�h�a�J��ú�T�nyX8��|`ϵ����:��*Ux2�.��r�e�M������\Ԛ�aqB���ɵ�P��6U��#�������:�Pbc�Xh��J>�).嚵�����U�	��G��i��NY�{��|�*>M���A'���}�5�°dϷ���⨩�Z��n���]E�oO��>>x�gS�.��g��3v%+j�%��'C�&^�aL�x[#���Q�qK�m��<q�>�i����l��)�)�Ki���(�s0?�����G�/�b�c�ew�"��χ�1�����=#�;������9��>e�������{�o����2�&���E[,�_��S����<����➪�L�_�Y��Nn���,��q���J��u%��[�9Ձ�Ds@���7T�4���R�W�Xu�u9�c,[:���@��C�j7B���o���p������%������/�f��AњƔ�K�'��� �?m]Q���秭=�+5���{Ȏ�����TƂ���u`���ǲ�
˼��䷞X9��N�	vN$��H�f��6L���}��U�d�c'��u~C��@��m4-)���aҙp�y�z%Ҏ��eHZ2�<]�����=Ac9-;n%/܁���c���>��|��ၑq�D܋73�� Wʀo��M�n�0evgܡh��-� �;x_�f�8bV��/�������D����De�m"��r��_Kz�!3�kU�x���Cuס��V��QU�MНDQ��K4��l^��]�|ozW���`��F#�;Փ� (fE+�SeCΜ0�ބ��,H�s�6�4*mquvy�ZS���r���P� ]�$�dt-����o�����g>�75�> ��)�|�����_7������d�`��v+��)�|�j����U��!���OC��E0�����Hj!�!�r���Ї$64�7�e"#`0�(Sm��'���@-�%���la�[����qC�� )�W��Oy�}k�˺wHɵ @?�@X��<DTk�ł%b-� ��
��r��i�1�a��5�O��7sǋ��,�z�$A(Ȥ�U�1ב[]���o/���:6᠍��%��������M�{x�LqЇ�\~�u=��,�a��?T�L����O���:)!%�h�s8���W��ۖJ&8��X�\z��x�/��[����>[S�-��4�&���&�\@o��_X�o��s���пe�)i/ŜǍ��l�w;-�y�����-�_n�us=����I#*�#��ߚ��9���;I�bWi�8n�讦�,���A��a�y��j��l[=��/-��BF�[2�����7�sfii��_�}&ڮ�8��zj���+UG�Q8�A䕼���_ɳJ��x����?Z��Vl���� F���w��CT9����=a��ўz���62����Z'o���d�vj�)w)m�Qg������3��=�����Ҭ�ә�N{	�:��&0��'"�Z�L����GԣO�l)+�ĵH�D%��$���,`��ԒXC&w�4(%G���`�a��^*4S��A� �3@��^��fm@��-s��ޞ�r	2\YR����k��Ш0�)mGݴ�C"j�;��GYdvW���vT!��n�?��9/�	��]ъ'�Sy�݃Iۇ©�g�Sѩ�q��������ZG�e.ٟdD{���p`����-�!X�-sb���x�_3Q�b�ľ�@�d�>=p>��[E����l�L��d���Ȇ�4�[J�/�d��(U��`��5G�S�|S��*aGjҠ?+d�qa=�ʆ���M�`o()�7���~/z�%.�F]߃��F2�����Zd��%5��c9U��m�� 3n���|P)fN&�$|O~�/�������!�60|����� Ok��fT�i�9�R��'�g=�х6䪷}~ί,  |�;<���fVַX{y��������Fvړ�6C��-��Z�ch,�Z:&W�{ǭB��<�Wc�t��P!7Ҳi[WĂ�������y��t �4C{h�ŏ ��egx �U#�Y���!��������z,?˓y����̱QY���N0�W?P�z:ƢWۋ���O�p��Ʊ��+�0c*P�B�j�qЧ=$����p*�*n��{!Q��Ba�oݥ�6X����Ǜ̵H$V1�[9s=OI�18��3�r*1�ĒL�z�Î鿿���`J�R$)ZVѫ��z��ͅ/��lk��L�"��N�qk~r�ժ�&��/}H,)B$ǻ)_f\�s?=ٺ�Up�^d�xvox��S�[�(��ըP� :.��.�=����5��<b�;Ȓ�x����e���oa�AY�;)�ܑ�(�ap�TLKy�cZ�yu�~�|ݗ#�B�M��r[."�h�7�Iq�Z�@Z�Յp��<��1�8]��{�E���N43�y���P��D��a�׌���3��w����X�2.*|t\!����r�!���@F��:�$��o ��r1�������>�ĬJz:�[��N�i��)t���N��P�o%VjOe�ח�(�kt�q�Z�̼~Sk:"] w�?]��s�0��_�ɩ��a�CLsR�U4��P1�J�S!h>��OyFlȒ'�>_�����ͽkb�xc��E�uѝ��]�߼q-6����JJH�'�y� ����
��JaR �ב5�:����ٶO�iA��َ��d1v���; ���֠@� Y��yM�^%�m�� "����o��뽦C��ĴQ�Ac��}��Z���r/��%ά~�e���hH�o陙�]�!:�˝ѭS�4ϧ8�C����7�a��p�̶�]��zM����k�	�>u�܂��$)u<\��xty�B�7;ju����B�L|��,Ra
�<]���#��;Bh��(��+8+�)�4/��!�v�$?u,����̆l9y��F�_�� (������?���Y�,��붍���V-
ib��2��r�T��l?�D����G�.B``U'��W�d�Az���ρ'� ��G���պJlcA�^T4θ+���v$�|��;w���tmTѩ�)�'T���x����{�工�m��j���;p)�C���Q��9Hh��f��ٯ9}_t��WK[Avk ��~���W.�'#�#¸��ǉ��`��?��l��놆[0�{B����Kk�
6�ƹ}YU�P�L�fV�ٛ�ݣ��#K*����̣4����wW��`"���(5�*��{]�}y�̷i�F�8P�Ĵ;�����ED�_�i���a���*���j�5��?��[�O���{Y`?���c}�2��NF=�V��x(��
��<�Ba���R�)��žn�M�4�ne/Vp���wr�a�i�2���OY���I�s�Ԕ@7������ 	�88���p���PM�V^��L�D��e-�YE����
�Ք�ۅ�>S$`��Pj�5K$9�;��� �i��V�Y�}��m`Z��X�J�;���ʨ�K��6�ֶ�sr�+�ZC���$v|���ã��r���V.�9!ev���6��l�|�>���J�f~�a�)�W�T	����j�I�@;J����`	��EĆ�~�%��S 2�+5����}�?0����
�r �#/��r���o���8�v0���=i�Jc7����糓$ƪ�c[�؄��{�_��ziW�r���a)^��~D= �8��t4�eǏ�(9��	Pٖ��n�*��~!(8��MW$�.<'t�i�9���BI�ٮi�F��KU�3��!��ۈk���q���鶍����ܟ�����۩�+�0���PG~c�㟺�:}d{�g-�:R)�1h�3+�ͳ�8�J��&c�F�D��	��T+G
qT����@�g��kvc��c� ��Mߋ(	#Rzn��mw�u�O��y1�4��4��- 6�;ٻ-�59�	�vy�ϚF���E���	��[��Kr«��uM�n�C�;��\`8X���o2�v3-��M��&čf\,���ke�'�kqF�A[q�N%�=쵉�C!�ل,Tw�i����<5�(��6{�#�Ĳ���hL�pm���A�cu)Н��!�3QG=<c�s3��-��,��5�k �I��Pp<nQ���	�s��p�*�D���d�YT2OS�'���*^HJ�؄DT;,�����T��T��`t�m�eЮe�mkeJ)�=��*uqD�����\�|ԇ;��]u�]�_U2�p���rP�yOԑ��9�$K� ��TJ���.8;�tP��C�K%n�)d����v���h�sLLǼ-�4�R&1�G2�&/:�L��L����Y,&lXl5n��\��T��+��TR����ā�|��x�xȟP�Iw�k��D��%F������9ʶy���0)�ͩ�e��I�� ş��K���@�o����;S!/��9��gNݿ"';����!E�y�1/BdɧP��\͗�K����M@�䓱��X��
~��k����Z��v���R�r�Ǯ�zTT!�h�����B�v�,K./�l�T}�+�e|��8/ov��]	���w��p�4�֯�y�p<Y�TK�_z��`Wɪ��Or���ΣGo
�N&�+�ox;ݐ��:����v����I+���;
��բzC�,�S�r��r�+.~�~�63@K�򲍽�6hY�>��}�$��}\���a��Z�"A��Fë@�(Y˞
J�~��t.n!�k^��������5�l��r/�����HP��sT\� ��U�������M̟G%q�jW���]��tOUYĕH^�Wq4�X.�g����T?L�5<Ҥ�nff��w!�����4�g9O-�=�Ņ�UѮ��ѥZoG$�(H" ��\�]\�R處��^����	,Q�}�2'Ʊ�>������ؖӻ��q:�=�L�����y��ӊ�m��w�s��ږ��T��r�c���#ֽG�xv�=�p�!Խ6��G�����S���b��
Tn �I�L4���������v�U�P;�'W���љ0+z���Y�����t�ܻal�5�L��dp��A7C�\�U`��㩏��
�K��:���{S��,��売�a�2(�	�6��j�ӷ�A�l��6�����tkI0����`���}�HR�c��&�����I��D�gJZ�Q
�Ȋ��S5�n.�Xu���hH	�7�H�%"�HI+���!�Ӿ��u�*&��M�n~vFHf6��k)�3��4*�Ŷ�V��BI�"�0��T�$� �L�V<9a[�Q�&��B1[H(<�z9�Sa�neV� �2ϸ��/it�J�M��Ȼ���^X�r�: ȍc1�V�,�����ڸ�#$V$���q7=d����;�ޓ�k ���YshL&HڻiA񴁙O��d��{�������c��R��ҟB�b���,���{q�#�Bn��oJe�l@�jT��{ı*�>�i��E�V(�V���x�)p$�S��c�ʄ�~�_�c���%c�z	�-O�u�EO����b0fĠ!��ނ?d�ZJ�<K�y/'֊�+`c�̝�I �^

��?9�O��V�T�"�<���Сh��`kW� ݁���t�"�>�̇�S$���TJ��%�*Z��(���Òk: � G�92O�X�bn")܁.�PPpo�����k�� �����
̆y�8���WE��P�`��&N��W(��ֹ��õ��or��D2����E�TL��~������-XS��uOz�����\q{�p_0�&�i(-Q���6����P����<ȅ�~����a��nUç�e�p:�D��M��p��H��B7Fj����^�J�"�%۪�
���B�C��f����:���h�?�(�(+����`Ϩn��E�Dw�Pz�W�	w8gq��4��FC��6A<k�3h�wZ�W�-֔ p�x,�@��Ͻ���\�b���ɿ�,�;�������T����>�>![t~$4��M��M
������1�:E�q��E�b�<RX.�W�0"`���G#b�������-�[�EõeFzפ�f�Xq}��p�y�Ѽ=8�����P�fd�u�胘o��O�_����J! }��L��
24ǂ tQ��a�9�5����N����ځ-��\hly�@[r����#��3��	�v� ��9���y�GO�|s���3"ڲ�ۈ�'�C�o�����٫'��(cp�y��(��L�;{�y�P_Q����9���i�u{��"������	���4�6�pyܹc� (�4̪Pu��g�
�V�<8�	��oހ3��ü�����rm�����v
�0@K����~o�M��ꔟ>�=�(!�����^���i�M8_�L�
:�-$;ዸ�"رUl��o���QF�d�&�UpG���9�ܴyP%F�]b�֔��#�V�OHs7�j�� ��'.W�v��jX=h����Y�p��r8���1 �豄���B護
N�A"й��/h<�@f���i�b �����6Eɖ&ܻK�3��Vf��_�qt]1�'	β��+�my�����Z鳥<F|lla�|E*�@���kQ/�����N>uؘqU"���)R�ni�������T�[c��_��ڨ�HA�����'���Cȳ��~#ڻw�Zꮧm���l���ª%B
!Ik)�9�࿞�N�Jo�W�h�8֩j��+C�DڸB�rx�hw���g��^H&X��g.��7�+n��N��.鞀�Ah~*_������a1�nZ���F�#\Z��~�h��?6���!P�v�H�h=��$�h�jK�b�����tyN��U�$��&�4F_h$�JE�v�;V8�� �Y��;��;���T:UQ�E	�R�����|K���>�!ۇbӺ�J�iP�o��Ɣv��Q�`ĥ�O�#ҕ��g�?��@s+�2����zl��M��90H��h�+�^�s����L�l�~	H2�7ptn��BGgh�C�KjD���R�ۛ#�{�&�d㿀n+�s��B(,�������H��%-�JB��7�Yq�Z����%I)�Ҋ;��͝WE�\��>��E^�,��OL6���<�fzg���wLuȨ�#u�Z)�:Ѭ��.m�ʁ��w}��c���L񉔝@�O�8��J�%P!J�SP9)�w���i�!��)�%b���#Fv~��B�D�����$Ebl�sM�Gⴓ�
������I��	�ſ�z��ˋWF�t��0,�B뽄���U��#�΁/S�174��|��2�.�(j��x�w�� �?j�=��*���P/}�A�w���#I:��(���Y�)z�-I�*�mD%���I#Ŕm�>�4|,lό�qJ2��(޾�x Il����QLD���2���j�UВ�'��<t=��4�O`^�b�w���T|�k����%O9~a���i�(pUc�Qv�x5P;���8v��I���96�Z���kPW9ْ	��0��e���-+�u�ܨz����LB��ʁ�T/mGL`��8ηۖ=ی����Ϙ�	{;��?�"�н�G��)}���C�i9)�`��Q͠�T�VT�0�&���ze!E��f�#�~��6�"gE6;|�����$E3�u����0�U�s��iah+T=�o��n�Y]:h���~�`��!��~jy,�3�!�T?!�Z���Yz%��Y	���&r�����K}��Q�pdg��H%d�:1��D�Q�W��D�L��u�$�@Q��7�!���=s2R��b��[KԎ���}�-�)��>�#8���� ��8��&TLy�ƥ�\�����
��J��d��IN�V�>�OK���D�
�1�R�å�B��o��5
�@ܷe3��)��nX�Q�+�MV���r <�T�7I��BְC�<�9��C#�R���2���	��i�;�4:��~�s7o����~�!_��O���'��bøӨ��Q�l2�(:摎�ye~�O��͕�vPj��82ʯĳ�ç7�N��z#��݈1y�*$SK���>��:�l���P�*���T��X�_J�B��+S���Ո���a�m�~���_��B9iD3�n(�G^v�;���J�����d����>�#&J .[�I @��c|��'4�-�d���{��Ptw���Aim�`�!��ʀ���P�Dc]�Ҵ�ݖ�3M��ۉ̈́+��|1��"r�!��_���:J��|�:1����ѹ�,%���a$�Aw���)gk^�\m�:�\3�'����V�ep0�2��a�o�����Cz��!#�v"���&����0
���2iy��X�NݯB���a��V.�B�OC�`����
/Lb����ϻ����B3�E� �o���<�	"N��f|�,$��O�N��,�u�T�Gj�в�=5���NYN3��%cP����6��A��&g�~@�H[�1 
-qϪ���geia�z���K�����Ec�8ɪ�ɒ�b�Z����b�~S r��������q��݅R��z� �/I��Wi�-	}Aڍu��ş���Va{T؟��3]�:b�+���L;�uCO���.[�'n{��=W�+��M����1IB9hѩ1w�euB���:�*kB�j�(��~�����M���yjT�����/�11U�tN*O�	seW��k�
�����\���pή����ll�[L��[��K��]����݌xMё��3KU"]�(8�.��t�T';�<+�="�%#���F��%��~h�21�لS����g�"f�L$q��5�'�0\� ЏzS&ُ�.�ҽOZ_9�ʢ�����Z� ֟4�+ǃ��*�!&,���c�H㬳�W�y�hz� '�ں�z�2�����I؈;�}!�N�'u�^'Qo֎�NH�C���'��Û���#EzZ�B�F�'��#O^y�*�n��M�����5�'�|���t�2 &qF�,��G��|r�+hƚ%�=���>��h�X���u��:]U�,���3��[��K�pӯ9�� �)�{��Vn�0~Q��+c��"Hvh^)<�q����p����HR]�8@,V<��\\�*�=�~�a�Zl㙄>���E:r���%ֵ(F~ǃǖ���X/g*��O�r(*�Y;p��W�����(�|(����;�N�)�ar6ݝ�C<��e�ͪI�}��l&k���J��w@Z������}�#M��%����:ݔ�r;���	�
�[������N�y�?ޝq�H�m2tw�fa8�Z�8E�(�@����RCO��k	�	�+ ������ ^$��k%hEQ�����$f�o�A�&��*F;[�[�2�:��p�Z*BP�D.���hzA�y��GW�Kσg%�u��������M8���ed�%$�N��ԅ�F>zTq�y��oX,�~�+�>�f΍>��s��T��(T|�8u�8Ϥ�
���D|���V+�!>z�ӵgFK)^����4����O�0�y�ݻ��vk�Gl�*�mdm%5��Bf����|�P�D����g���+B+�)�Dɩ�� 1m9��*�"�&]!�Q���lB%\�'UM"�aUH����0��J�&s�U3����,�
�߼v\h��p���~+�T8�o,�NԒ�bM<�]�4a��V|ɸܺ�
G�:�[
:���$a���P���~vNX�V�|�s���gF�&�����,2{�E��/��bp'�&�;*ė���W�{�)e��D�o���A�4*�L*vc>ܟ}�`B���p���W^�������b�Օ�yC�vD);�/@��7�rl~X�Z��K wҬt���Z~��C�0��9?�ש�H�kz���H~����n���rK�<���f�f֖���M�"�]��A�vC�E�D�5��#�	QX�;n�%������(ȿ��/�4w+�!�������{�8b����ZM�eI8�RȌ��[@e��XLG'FD�u��9u3���9R���Kr|����;�Y�a�9k���a��_�fB��_T�b��bF�\Tp�����A8v�$T-A��k!�?��?b;M�1g�����e�� �}r"�6�qJ����"��us���䞣!OC��qhi����~�\��n*jS4^��\�+B��I :+NӔQ���;ؔ�E�
����`�BHZZ��t��(��N�34S��+�k���%�c/8���PK�,���$�mp�M�����n�ةe�#@��æ�|H��Mۋ<����l(t�S	�gǓ�B��j��
�%�II^��D;���M�_S�#�v��#f��-��%>|��f�7�}��Y�Z���n)�+��j�,�A׷@��>�i���h0Z�\�D����R]kW�z��U+�Wd�g��%M��8\T˭� ���⾡7�υ�x��rQLb2�T=�l�y�:P�,�3�J�����o@
��B�Sb�H��t�Bri��LRk|\5�� ��n���kr!�ᱺs��(;���6�!n7w�_�]as�͚�١�f��dެ��'��(0�����j��C_^�6���E}����p$���ăl"�i(��1���^VQ!�
(I,˂�},G+����c�Urt��!�2�����C��l���v(0|���~�h����ė��p�w0p����V7��)DM���ܜ��M��x�+��˦��V��<{`��e��;+�r7�I������Yfu�vn��0���U�6 ��se�8��)�8^�괉�-���o��
c~�W��T"\6��������C���d��P����YM��gNڋLß�c�Ct�����5G;oF4�'Q�ֶ(����ĭ�������.$x '�?���!�V^�������>�#���BDq�|h���+��2��k�׹�����F|v�������K}��t� �QjBT5 �y-���𖞩�o�6Rڼa��5RC�&mȰvz�P �B��bz��<�Q�o��}�D�)�����n�"{��1t�b�o�#C��0l��]C7sFxJ�f�y+J=������b>�DA�*���5�p�>".��h�p�������Ҥ��3�iY�H�5>��cW��9;7ҥ�4H`#C�sW�kU����;��QӚ���!�H�4}V�[��|�ZY�%�Xa�Ccz1��1�q�����奩�Jq}���G���a�yz>��������v�JR�Ƅ\FSD.;F����%����]�E"�܃j]�&?�[3�	�,$�����=�����H�¶�k]M��!B��S��~�|�2��we�;CE����giqoLA���L�ՙ�0�����U���ܹn�<�RĬ	;��B9E�������0�Cp�0I���σ�y�^C7�y�`~��z�;\C�����t��������A�IS��
������@��4�-�_Y6ץnHHp�όW�m�fBRT��vU�ߛ/~�b���c̈́�VG�e�iy��m˄*��}�6P������3f�Y��ܤ�(�x汿=�J
{�9��HCJ�X�����"�sg�,&&��)Hݴ.��(.���O-���j2	M���Ʋ�s>8w�[�����>z��~o�e��s6wޜ�&�?�jʪn\��\}�'��<�������2z�ꦁ�.''�r�iƢX���Ů��
��ԡ�t�-1W��A�d���H�X�U��c��TF[ƾ�<�=c��ׁ�"�r�������������C"�nP�:���e�%����:��`�2�z�\C�Ik+�8>G'n��&�qË�롺.ܼ�#6�G�0}Q8T�$�~;ϙ�!��"��|"	���H{N����$yD�ދ�	t6�f�	��������:� .Ԅ�`B��j���� :������!V����ӗ��g����'@w^ȑ����:C��\IY�R����� ����Su���<�B�<~�gP�r�P`涞Ç^3׻`��H��9����S4@����__�U�Y�Ġlv��5`�r�6h����\G�d e�}����%5gj{��'�o��}s��(���3"w��`�f?H���ɈƤ��ǚqSP��sn&�����y�ף�AN�S�������@����\�� `{p�&�8�ne������<�F6�p��6��ڷ�,�
�^�wI�����n��9�zFJۻq%)�-��k�i��"T,������	�w��[�)�R���ŠX�(s#<-E������%�Ư�8���h!e<e,�����]{s�Ю��=E:;���5Vs��z~�M��1�1'���k�'.�8+9�Y������+��e�j�[�=c�w ����U��zT\�1��_z�{!�[Ia�=������Q�)�#D8k��9�m��i�d?X{{o0���wy��6x�v�@V��J;�.��I��4��a6̚�:(F�P`��t��>�%��I��g��+�*ó��q��@�
xW+�=d~�B) N��%��e�hR ��������*k����6���p�����NNx9�`�X2��To�m��y��@��Z���$O.d�k��)�U)xߑ(}��}��|��ʋ�'�*�[��q1֤Pɡ��8|T�P��9ռ�����w��om?�:F�t�3��鴼������PAZ�u��E�9��zDP�T���Q�h3||��N���5���Z-�]������oc����(N|��h�@��o^1��}(��)X��xլl��c��ޔ�6'��5�D�z�R8Y�l/��%4��N}:��j�h,���@��@�>���3����K�J_H�P���F��/��-p�ǉ�mnY��U,ZDt{0o���61�*�ß0p�t�;0Qt�\O3w"Fw\\7=X~Lch��
=�y�����)��ص-�P��|����q/bh}}�Ho���N6���KI�x�71=n��Z˧˥c��M���o�.�GQ�3�� ���Y�Y�nNKr���ۄC~�P�:uT�͟t��c�y4b�5��9����؅x_�m���Q�����[C)��r� ��:n���ͤ�m~3���ǐ[�E����h�1��	�3���,Go
,$�m��ϥ9*�nhO��w�@C
P$�I�p Ԥn�yԱ>ů� �f�ߋ�͇I�˔�>�D#���0�yz2��Cr�}��4��(3��@��
��3"�G�C������qR�����gwM�<R⩤x�ک��pX���k
�ē<@�w�&�N�O��>r ��'B�!R.�`�3�{Iw���(��OV'�@���G�����h�u���Y�	Nz�c-��qo(}s�g�}`��G`UJ`L�"uF|�D�l����p=�U�_���Q_S�a���m�w^�,��h�k��	ȒU�̳�z)0�:�����^��˚d�v"�h����	X���ś��z�fs��Os4�M3��З��{�E;C�c@�ug���,l��i�]����o.F"6T��A+��Ӏ��ݔ5�˫K���݄4F-�=���Ce �0�Вu&�*�
n+��[�h���q0�Q �w- ��X��~���a�Z2о�)u��M�95��^l�]l�xa��ϐy����s~/#e�'8|N��^[\N��bc�W�πB؎����r�V���̤i� :�&M��e��C!�t��H�^L9�<�ï��7�U��<Qu�a1kFR<��T��u�0֙'�E� Z�lH��󁐱Cܟ�m3k��*L�Ѣ�O'�t�M���Ԉ��>�>j]��q�Y5y�{�X����d������&0!�  Q���t9B|���q���RH}��5Q���&b�l$�1�[�do��ݍi�=������rj&�mٿf^x�;͋p�=0����P�;В����ɨo�fn�����.Z|:Fؚ�t�;c%rNQ���?��A���W�޾�az�{�^�68 u�@���rp������2���>��f�ޅ��@��7��#��@�o�,�������c��bhڬW�J�S�W8��D�v�\�X��X*@lw� ᒝ�Pܪ!���V��|�ۀ��X��0p�,��e1�kʝ}ɂ����(e�(z2�d;��X�=K�+4��*�T&˾�
�1J�AJ#$�F�u t}�!�!
����LaPEK]��[�Dv��H
j�M�b��i��,�b{a�t�Ը
?��.�J.��G���Lw$�/c��^�h�RB8i�b߸B�ʀ��iÕR�'�NյY�����=ΎW��z����<��g5F�e�cg�d�d�8���n��:��ۥ�b�2��������*=
SD!���N@4���E�<�h��o�p��R�HQ�ZH9�S�z��Ze��;���(��Dl~��]�z����%'�ώ���"�/��'NQV��8���%4�pƉ�A�M���<�ˁIlP��%]+����ٚ��?���	>M��N��])a�!���2�Qy�����K��	x-��E��aA���(k��hKq�aYa��
_�x�ȈUCG�ǃ"�5�SSbe��1�����	���OL�i�;��H]�5/je���?k��i{x��Y�	g&$�G]DY��z%+Z���޵�5��W	6>4s�*���ħŪ �&f�ج�%��.�x��WQ�o�:�\�Ӫ�cqb�|���?$���3�HrP��$D�y�T�!����m��s�ϼìlc�vb��s`m�����`U@+�C���Љ��
������#�@5
����}����e�ܝ�>Y�'p%��0���c ���6ꞈ�%^��f6���1x��rʓT?c�^:�斔i�f.�Ld��)NG)n�{�j��g��
��"r�χ=����d�xn�&��ܖ?4�
���9Y���w�I�� X����w��ak�u��`��;C����4�,��f�#`!DA9L�B�d��ёM��R�Rh��"��A��iU|a@�'�D��&SI�@��EW��4v��<n^?9����A�w�ʴF���[٨Q����硵<Tѷ�� �S��h����R� �ov[���:� ޮ��9p�=A@��-��͐�)���~�HgK)�Uc<ɛ	N��w��ؙ��Y�4��xF:4�̑p��J�X�q�����E����e����1�`�k�o6����*�B�<�qL#�2��8	Nh"����:�S��T��h���uwo�X�&��X��
�nA�{cfJCk<�"{�p� Q��o9���a����1�HR�Ƚ�:5:�?��&����?JF���
����ů�d�R,l��쁺5�[띚(�a>+�RE���)��x���<}%�d��T�6���*�T&��H���5�/j�=�S��~��=@I5��>� W���|�p:枮;�u�ME �&�2}2"H�ܬ�!�v��p��`v�_X��N�T��zg�)�{	ka��*�߭a꒗�KR!ec�}�[�����S\_7L
ٮAɀougOd����lW����e-�(_ ��X^���9x��>��5A��$�U���Qj-L� J�%&݄�+�:CT��7�w-V"r�S�h�.S�ɛ�&٧�l�� �![eV�d�Q[j0��R��%�`�����[)�-W&����tF�J?���PI�L7{�J��-�7u����N��=�=܁R&d�Ԙ���Rgv���(J%4�6�����H�ʂ�$��bXI,*�B���H���������E|��|/,�r�����("��7� g��!!Ro)��D��U�8���R&:�t���9}H�G�Ӵ������8&�!�3Yo J�D��ts$���2�V�� ВL�
�V��1!=��
�5����I��sTn�C)�J�d)���׾�?�|���[�����v��Yf�.Z�l����J�Y�nk�j]IfHM#"�����7��)�8����[��m0��X��&��hL�;����s��p[g��ŏ@EK%i������jX��,��<������?e-�b�~9��v0fX7��Xe��؊��	�Ps��Ow)�g}�^�E���1�sR,8`�t��.?/W�EZr��]I�2�h�e�2R������Q��e�a���Ś�1��g!�~m���	7��fkw�ُ�'�j�h �ٱ���l9a�_E�-stJ@�Z�}Y��k���u�/�PN�-`��ZsrK��J\���\�<�JB-^��LN���rm���Di���ON�,Y�����<��#�h���;�V1tu��]5����"+��w.��q����
e�yl����4�_e� I:����[>���p��~`/_K�h֚e��O ���W*�^��d�a�5k�4^����N���SC���1�7ېc�aR�f]�ipHO�Ҷ�8�^��*��/�N:�L�����<6G!�?CV�ӀH]Z}��2#3���۴
�1�E@Y���m��[w����7�8�O�@��:������&F������c��	�1�i��{J}'m�|4Eߍ��q������F�X��e��5~Kcă8k#�L׌uaA�_P/�/�|s}(Ya#K��8IdJ���p�bOK`�%5�XW��	���C��4$���C�^\m�-?�T߾?5@�ۀ���}�(N�s!�U+���b��"��S�D�z�'xv���q@�t1�+���)�����(��4�D�V��d�p�4X�-�,���)M����fph�AU�\q4y՜®R]�Ǟ��K*�Z��(Z����/����eͧ�ܴ���/Y=�L4�෸A~��� ��Ӄ��Aqi���"��6lҙ<t@yO:�ac�=bȺn�r���C�k���
���IԂZӛt��ײ�0t��?���_2��nvy���$�=�3_�ڙPz��#�����I�Fߝ	�.m"����dC�	�F�+���P�(7r%�۬�r{����q��������m`9�P��!�_n��}�5J�h�|�"	�]�wlj�����ɤЪ	������|���"o�Ü)��+9���7�O��	=�\ 5�~�'TΊn�w?�`��P��$�] 3�{y+,}�.������0z$5���؂�[���}���9�n���IF<�2X�yq2��6�啑9���5 Z�i����D��z���q��^��!�y3je����$�2�		����pZ�1�V� �mâ]e^��S]q-'=`�����c�s�c㗧^#�4in{�8P��������#�|��7���cs��'�i�)��Wv�btL%� v@>�� �`,�t�f�e�(���\�R��q��g�k��\�fLl��8y�g����N�uq�̬��ű/G��ݏJ^zz�ݮ?�C���9��kE_����_�M���e�M)@��}F*'�ŭ藍ɭ>�_iY������9aC�;�F2�8�x�Hnr�����%
��a]�JG��Sľ�C�*i0�!����7y���{q0�]�o������P�n��B���mL��:���~m�؍ڼ;�Ü!��ӥQZ�w5����!mu>E�pւJS��DzL�U0�����ip���,���H�҅0�*�1&���Q�f2P�����sOx��� ��,����>t[=v�ݳ�.Ixk����([k�7:����N��R���3���[,���s����
���P)�C<.�QWcv�U
fۑ�Y�>�p~���U/����7��*�s !@��[���=_N$9�xMHN�0#Βu�5GW��b|&�#�:�@����=]��	�S�.y�{����8Ƒ�^��X���n��HYd�cVH��w*`e��r����e�O���+㡜���4>�0�>/<��H1YˢSH���7cvCNIȦѨ��?S<�Ý�Ώm��x[�NI[�u����u�cN4Z�y���ؼ�a&�매Qwk�����'�:j$���;�S"��"��++	��(B�K��Q��P��u«��|;S�
��4� g�����F/� w�~��W^S�[d�<�h�[S;��mG�����[<L}��:��9*�܈`Msku� ķ2�PNtG;#�C���<Ʒ�Z��@�1�GPs�Tƴb}�k����Y�B�:ش,̢G��LS!k�pU�JԹS�r!5b>V���i�d0þ6p��'0��P�����7ɽ�Б�T"�ң�$�~� h��&���9̵v5�uP:�Ǚ�\
�2.�_�l�*���I������n?!���EtzT|S4�T6߬���V%O� A��/�!�0:�O�d�{�HN������?ߒ-��n��ZUE�K``����]��2�-6f���.�׭2=�T0����E ��;%)�>�a���:��0�� �S�f� Px���x�hY9�����a�`}���4���t^����,�%���b�u�N�#ݣ�l��S�[�F���L�$�]2l_�a)J͟S��/�Y|J��K����n�N>>^���ez޳2S�ɒ�o;�Z�<����'���©����rH�,�Wx�L����B䝐����0�)�T�..�Z
pD�Y���93�b��N�ef^1�[(P7�t@��_VE؅���Z�\��o�h	��mx��9p����h�k��sl�>η�� mu|��|JM�2��o>ܞ�6�QW�jo?y��*H�VQj�҄ ղe��2��cM��y ����i�E�$m�H���9<���!��j;�/���|nc�s�������9�&���܂�F�J��P���eI���HY�鸯�j�"���+�d�W���4�J�ʡ=à��BǏ��� M��rм_�0{U�/3���/t{��5���V��]���@�1!�O��*�ˡ�R�q1
��U6��.v��f?)�v�2�t�p�D�n��}�j?��{
���_i��V7_��J�O�+���I��� (���]?��O�A`����1�G©կ~��wV�y3n~�E���k�P�W��^hY���ܴ���݆���`/���pCp�sZ�td��F�o0�\y�R<�m��k"�¹�=��e��ě��.�&�mŹj�Nk\�E�&K��ŵm6KC��4��6k�ꀖKkL�z:�8�3$�t����ඬ�%;�/i�Ay١<�]���H�c���y��(1h���-U�MQp	ƕCG�x�hv�.Ȅ����̡@鹉$ؑ "�RŢ)n1�U�ݿ�jϕ�J�D���e����1^�[D�+��� ����B��LK���b%��"$c���3)��Ym	��4�&��ךO8���|e��u'�H����ʝs�ӦBo³��+�T��9����K�:n<w���[��`ť#�J4_���uP��
:�\�^H�c'��^�r"��4��0��qM�+lKs0�;�Ҙ�b>�%�M?㐶�&+�5��Ý'8[��Fܟ!Y��5���䟎/���	V�A�?UvG�n��� }�z�nBY�G�0����gy��	,�����YΦWftǚ^N6�A��+�E�Wwd�~p��t���z�w��Yr���'whn Ɗ��B��B�� nT�(�f�}��k���Tv21"���a��O	j���`���2Q�i\a!ʻ���7w&���O��鷧;�Z�Z(_�q�g%c�>���}�rVǕ�7l걔S�d��#�:��B�Y��#�I��4s�9r�@�K�A^��7��GJ�_L��q>?6pyӧ�|Wa���t`_[:���>a���T�Id��g2�zƊ��T7d�5g��Lء��ҍ�4�}��BS���$Q���[�RG���}r$�F\]�1�©sUx�A���+�e���g�87
��M�n9���jRbS��F�+��N�J����������i��P�4�a���>GV"�ulP�c�%��Eķ��L:%��OWV[�3P� ����ޤ�s���ʔ.�e�[��F_\i�7`r������]Mc��J��>cX�Q�JD7��W�#d�;�0ESR��"�Q\F������� �g*�[���ـ�@eZ�>ޡ��"=[���)� Ԋ�f2�E?��?��Y9�x�S��Q�G��,��u�?�����W�C#O1�	�������^�A~��n�v�/�dm����\��H�w�a����Ћ�bB#GIA�ꃣ��m�����ᚙ����F·k��\te��c<"�]IŊ�<�:u�=٧zOlb��9�F��DD�I�S����ACȌ�g�!`I�Kih۴�LRE�c+�ng'�J��c��i�X}��������|蒎e��^�ڦ>nJ&�}�ݠw��1fU�9�Q&���E�V�'�C���1��w'�B��St��6H��`*�B�}�^��A�|Cj�pPd�9�1�,�8�Nbg�m��Ƿk������Ī�\��_�R�ʿAD�����`��~ �:W!��	�A�7���q�Z=M���ak3Q#y�S⹒��g�A�0oŚ�M3���𷑖�|+M�9u{��B����R���SKh�U��H^�[3�	��c��G�7���Vi�?C��1��;�*�lz�����-��rq\��\z/g���U?���@�s��>Im ?�6JHND!�����q�qﾞ�SZ�����[W�jF�>vޗ:�R�$C-N�݃ʑmi��Hv|v���J����?�s��aA�R�!]hs='�	N��$I�B�Nv�O���{����C̸%ҙ��j�2gK�9�s�jm�f���ѳ��9�f>%#�~*u~�5^���e�#��������
_\�Hu��VRPys�׉	1E�!7��,�s�z''�}g����LĔ��j��1 A���7<��g�a/틅������'�ߩ+�w��$@�^��;}�2:���[�A0^�N����
�'�nU�z��\M��L��]ǃ[��7t�w;hdY��Dv�dJ�O��%���P�4��V���ޭN�(b�
��[�'��B[k����%��|&e�|q�w#�V��&��F�����O��F ���:�'���uz��1�KM�BLpk������8�6>+f~D�/�'�[ޮv4K�N�s|�c4��Jz�KeԆמ���!����.���[̯sW0|$uY�'��'�l=�i_��r��i��n�7��^	1█Sl��Vz�Ǫc�N��u�%��������-V+@�՞��E���Z��u�"&4l+��t��t�)�z�Y��� v��>O�5e�4$�3�M����톷�¾o���OB�3 ���?M��6�*y�5��\Q�襶�HټQ�b�4���d���%��1�x��Lz�>���x�Ŝ�4k�3eVuX,(��U`�:���KB�����8Km&�U��ȴ�OӇ����	�X$�s��'�b���h��n�޽�.���P1���H� ��}�R�i�"TP ��X��Q�a�ފ�y}�U�ͽ8���La�� L��������!��	M�zh�->*��0U!�	�E��R���օ�1X1O��R>�Է��;��f�-�~��^djK���<G�5�����ܡ�����>:;��H�Օ���5�;�TZRy�>�dS~�"-xw��ӭ�ٻ���[��iq.{�?ٗ�b����q�0Z���J�9ڬ��T����JO��@j[$���֏��ğYT�s,�-sL���s�B��Zn����fU}�H�,'�Ӧ�,�% Ӂ�R�����	o��"��� '����?�Ĩ�ա���		T��#�15�{���$�MtӉ�(%��;z��E"�k����|f>�8�3e����
��R�e� �`��)ϕ��)�y�ܷrw�S��|q�a���j��<9	h�?�������Z��U�.8ޢ
��������k�� �:�$%ˇC6ԝ�e��c~&���V,����J���\�]&�[��O�7�C7��Pe�"�s{j�84�oa1J����>��_ygy�ܐ	�u�k���SL,�#��bZ߱%�7�\L�q�4�Z�h��-,D�����UdF�X_���4�B�Z`Ol�(��ő8.<�"<�)��YE��%����jyc�����"�p�+0��Ge�P��p!�U-�ʥ��WΥ�TR��F'sRF��1I�́�����͠ӗ�.N0|��N¹���Zby�ه&~p7%���0��fD�ޞK�e�~/��p/'�O�-�����OY�E�5j��hz�� ����u��{EH�>�Å��B֟1��"I��lEE��(��:+��x���=Y'��W��8���BgE��
H����˧F�d`o�DD��O��� ?��M�^�f_?�3D8HU�V��r;f��H�y^�p,�5�bA5p��\�F��t=֖>ĭ��S���<�^V�#���k���1K�!ч���i.��-r�y!��([z�9��߁�� ����#Js�q'f�W��ةO�߀��]��5�������=_A��V���{��/� ׉o�Dd��4�c�ƹyo���]��aw�a���4�A�H�� �	z�H~�P{Gs�H,ѥUK��KT����׹�0@�XaQ��w�����A*�kL��]��w\1�/��RF�ߘb�j�2�%�72�4Z����y_a��%��H,i��9yl�N�*�'OB������������#�s�3����h&��P)P��a��|�m��6���D	W�_�b�[e���� ��U+�b\�`�+pF��I���J���\B�{:d��%n�4z�����)s���_t�G�z���U=uEun�%�)�*f�r��"
]�����`A��zw�כ� ���u�#�mb�F�*;N�l��ޚ���l�l��ְ�:g)�.�\�C�H��}��*[�"kf��7����ם� k%oƐ�������D�����9�����@�&ie�����a�S
�g����������O�X[~� �4|�|��	2]�8�䜸8'�B)�N蠮�)(70�eU �Z����v����d��Qn�^�a@R`J� �����F��$��'Z�g�V�!��,�����A��K��ݤ&�Ef[�{9�^�v.���aЙ���e�@b�Va�{K��m��<roڣ�u^E4TӮ��#��P��Շ6��ϻ���0�/����7x����2�x��W'�5\�o#����39h�(���^�|Wإ��O��"��2�n�%���P3�/��r��Y�����d����ҷ��J�EH��h�ИZ֚�2B`Ѧ�t�cO���8�3�ӲͰ�H5e�?��..�0�+R���mdH�2��).2V�������pA�յ����F*���Y-�������BBl��ߑ�������=�\����f��U�7$�ñ�ÿAT���E(�6���5�{�o�������g�*G�����<��Qn�Oʧ(͇4jy�?������%�J�s�"k����B�)C��*�c}f�d��}O������� ���(/���0R&��b7FH��ry�����t�n�P�,��D�V�gtx����L�r�h�!��p&����ܧ���I�-�?��1z���ղ�W�#��]@�f9'����g�RHLղ9���Ӽ��6 Jѐ�S�����,�jH�>id���D�Q��a���cv�r�f���yY{gY����~����td����97��<gFh������ٰ�!�l����5��h�3E��jsT��M�f8~Q\ń���U�5�<7�;�Z��Æ���ǳ ���2qG�S�Mo�G��]|*-z�e���d�m1Sܗ��<��?�7�<m����|���mi�b�JX�.xJV2�q*S����ľ�)֞��D��f�T�Z��9���0��gǐF����̍����lI�͵]6"`���OU��P��2v��ͣ652�42��YE$V aC�2Qa�He�xl����?��'W�ˍl�Bx��?DP�#��$�������]���t��)�.-�	Kש%�1�
�軺��1	��>���g���+�%� �B�+�r椁�N`̍�W%�����qfS���OΘѕ� �}���I����9aUr0ni�Q)ߟ�2�[E|{��o�M��z�^������/��b�/� l&^#+9]\�g�ՠ�ˁ�T�gWK�R�P�?�tMϚv�34�1����Rޭ�2��t�����f��y}&�X��"5�~�ko��Jg�Nݮ�)���6�-{���_����CD�/O�sw$c��{�RCDw�,l)=Z�ң�P�sb�L�]-����l����/_F���ad"�Fb��\�k��ہ�(����$l���"��Q�d���m���LgS�a[mÁ��x�k*h��|�obA�A`_��`g�𝼇�)�p����R/�L����7L��%AH�!��kB�f��A�\B��M+�^n��^[���\�o�Ѷ6R:�oF]g�
���Q�����Aa����(*r�`gKE`SQ���6�� Bu�8U�*Xj�����aL�� =���"U݋ioh��ɵ;76i
&�O�z{�ol�d�Qk��f��Ȼ��2�Fxȓ���M++l�_��_��'��Y���M,K����H �~A}�H������?sO膱Y�E������M�8)���VNi��]�G��������$�-r�HK�Z6Կ�C�?���K�^������w�-��W8�tVď�)���L	R�M�p#��UPv�nV��3O�Qh���O��aZ<y��g�$�`։��S݈j:��P|x�0��7ī-R�?�<#��$�N�{���7���ov;��P��wǕ�+�m��ٖ\ �w'X�7F�l���ߟC�|ǳ����������ۍ�}lc�u�����2��y���Q���
z֛0i�j���Gv�9�kMj�R��k��#q'"QGʛ�5+c���,
��U��Ԇ0��0�YC0�̅�CV�>ܶ���?Vf]��]��O��_u� {>܅6�y���j�03�p�"���[E� ��l�<䧽ϧ���_ �ԓ���r�U���7p��V��,����+��n��;ﾤ�+��-*^�;��5y>���XMV����qZ0%��n��qw��c�Ox�6�K�"*��9#3K���<����Ї�Xfz:e�Q��}5N���P%jL�?wGA�7
b�$��cCe;�������p�^�|t��P�7-�W���O v�v7���z�u"�2r�U)���9 ���G�{PF��$��b:��P6܎���M~(1�D�属�Z�}�%U* �6`/�@Gs4I�UPS�g��n�'oJ�K<J��` �� �0R4*���ǎ'�,ch�>H��XHe���W����S��ER�ἚY�إ���h�C��a0�w�g�p+w��#M{�N�ޅ]�i������x���F�8��MG���#4$*�Os���	Z����$���@�(v�Y��K����L;��Qo��-�a[�hIÔ����(KjO����P�ܞ1Zl�})����C�92�\ڜD�Hhb����;���1�mEsߡ`;N}�.h�_��g׆cd�l�0��ǎ?�π�l�B���nt*[�E_1�
yjo<b�3�x�tX:Eү_Bo���
���kq/��^�|�1(���J�GlB�w�*�ǭ�.�ęyj�*���J(80u���bR��;"��vM7� �{�T+ka"��;ު��3Dre��*� ���0���K�%�������{L��g� dv����Q��[���&�ʱ� �����2d$����\�5˟��Vᶥ=_�%^��_�gD�3��C3;�Q��D}A.1����	�>Y�MTy���%�ˤǌ~]�]�#����xo�!�z'a0�/�1"=�T�SE�f�64�h��~ Џ��o��3c�2�a�B�ui�X!*�(��]��4�����iShW��4�:_Z2���1�ɴN�oNΞ��N���2�gX'�X�J�?c�|k�^�D��|�"48oZ�j?��dt�8��w�tU6�����*l�ܡ�Zt�!c�F���b5q���؋x��T���;v�9�vcy����U�(P�C1r��������Sj��/�&֝#�./n�Ղ*���"�8G������Yt�/���"w���9�Ǖs��᧼^���Ԝ皵�(B a<A������D��� �щO�E�q�� ;��@�x��T՟� l��g���/��C�ȟ�A*��߲� �U�v�4�]v%��2An�9jv�ڐB�#��J�Ǎ��Nw�O�"����_�,遄�m��"k�_cCHԺ�9�����t�MyLT��",g�p?f� '�nEu�ݾC�{��J#�ŝ*���?�)>'�'�Q��	��ܼ+�Ut�0�r:�3n��|)��U��8A=)j^� �]m���jG�����5���d�+�u���IWV:gA�=[��W�X�����6���S�z �^P>��P��625��T_�S�P]�M�h_2qQ�C�TD^b,��p�yfF�ɼ�s����o��+uA>�ʉkc
��b�夭� ���ew��d e�5�nj��׽R��^���<bEh���m��wօ@��Ҩ�g�T�קQC7
�֏��Qөi�x�9�@|ꪑ�#����M��pI4eoYU�����c)�����מ�W/2����+5]���
�2�α2�4};e_4��%Û3����%f�_Ȯt
��px�,�<W@��H'B��I	,�0&����j������ju|�"L�#CKEխ�X��ڏ��e��6��!�do�
�ہ��*��>����^=.�ʁ1�@��2r�ۿ�wŰ�.�IK2�ѕ���7RwrX.F�g�|.Y�YHͤ
,Q�{\0I9.:�G�X�}(_ ��q���Jm��W�!��[��`�'���],���5�3�߷��S���Ti1�L�G��5IwU��0��8����߀
N1 �n`d�ˬ"�rEJ^�	�x�t_vW�zL���O�4��P���|���On�y(~��)���Cq���>O�f������������PS��8�j!Y�I��q�/O���LRI������\�_:����8#y�s@���4�p�7E*s���4n������y�cs�<��Wl�e /[�t�'9}P��5��R�BY��N�T���)lT�=�k���Qo�.�m��;�L?r�z�U�iB� ���*�~JU%Gpׁ�Z�3�ƺ�x*Z�r��߼o��Ǩ�G�颒M���n��e�(�ޡ�ƾ�Q� 03OA#:O�
s��j�ѣq��+�Ե6�ѵ�_�i$mQP���/�`j�� U�'�j�k���m:)�b@�L�2i����O�E�>������q���.k�F�!ȓ����������>w��u�$D����[�.��pm����vg�o��9��Bþ�n��B�E�B��&,�U�"�VA����������+����^/�5l@1��-n�`�?
��=��c�3�W�}��q�cCZ�D*�u���(	,�/�o�d��Uy35�hȘ�5��1�������i"�N,��<k䆹�?���Xd�Nr�PػQ)�=�Q&�^t�i���mcb��5O��gŪ�Z�:<�}��G�SD"�͘�J� Gx�vgOd��΀ۡ�6"��V^��V�P�k�V�*��
:�!�o�Wa�s���!{g�U�j-�8鶟/��g$�Ή<�������A�t9��d�3�n2�j�����h��g��d�������<�����޷2��n��aa�oc�a��w|�잸�	�����"WR�
��@��ޫR�Nz���_<'&nO�&,�F`̬���K��(P����z��J���;(�[󊄇��b��T�A��筿�L!{& ��s�:�l�� /&�#/�$)��T�q24K�7޷s�	����d
�w��p+a&6���bߏ_3�\(E7��Gd��A�&^��F�����I�n�W�xlu �q. �,�Ã1�L���bJ�/�+�ۺej��|�T�z�,��l���r�19�2��b���s ��9�c���L����M���oX�7ar���-"��_��WP�F�n-^����g����7�|�tME8� <�5����$���q���D��G�$��Dt����>Z4-�����C��h�����^�(v3��tl.�u�^̴<�.Ӏy`(�z!$��p�2shQ�j)�Ma.�P'��d(I� 3��r�n�(O\�^�T.s*�����w��������f-�N9;t��,�8�h��-�ճ��U�V�|�yqȥ7�1�JMl��$�����Ə.s_]}1�IP��W;��$��-�Q��`ߡV�����i� 4�T��ta�k�9��0>H�/�EP�R�d�>������uUCM�`�%�a,2=y�z����}����h�.Bm_M�]#!"�O����� 75���n�wR/��~6�}�PS\{:W'�w�-�I��0+���M+�������S��<N�����,�-2|�ܰ�.1sZ���a�}1$
�R�7�zM�E��O㭴�9��!Xѻ'�J�j�zb-�~�����Ү�<��,e��Z��{;��X��q����Eȯ4uf�^`�����\�ۗ���"'��@s��1���?�p��R��X_bǎ~��e��/)A�������C]9��W ȷ�9��^�+�l���E$��_����Y�ʇ�L�K��^6�=d7Z{RoV����g���Pr�u�`a�X�y,�=�a���/���L=r4n�M�I0��S�U�S.�@�?��(Ye��¾k�?��Σ�^�����i;���fC�Y�w(,�Zw"�lc��'�.�$�%9�u���Z�Jj� ��Pޤ��JO\d5��7l�f�HN��H�u����N+��4��LmuN��{ү��t{i�́��p�w.�]��Z�A�M^`�MWf��H7_"|aŻ[�b�IXu iϱ-�#2�H,#ċT��8���[�)1�o�5uJ�X�R�EԦ~����<�(!t��t �n+t�ˆ����q
�h&ޝNm���5�o�ۆ�;ԭ}��yؙ�Ə�hy�u�m�^��3�� X�!�]�����-��g��\�q���o&�����4|��� /|t���DE���S�D{�Y�\f�FO��#�#J���
t���
��h�^������#��]���gkʘ�a��U��;D@E�t˵U��AN{.+�>mz��=놡m�|�AC��9�zLЧ2P�Y3�	|3�0�K"�(oB|&�jiܺ�z-�ZN�6�U��ՙ��Y�{���WR��;�>;���}>�vl����|��1{�۸D����K���U�m��N>զJ��W�}]�3�@g�ԧ\��-�a�M0�#��ݮ� +��7SŬ�_\I�q3�q�^��V�o�i��b#�/Ë�T& hU�M�~��GO/���XT�r惖cT~A�HQ�ű��RQD6�V(��T�s	5��-#�g �O�p���4?��)�����^������F0���7�`[�8В�idlE�򫱸+uR�]�/l�z"��)�N���c�'��k�\���5ڠ��wd�:I*�r�AJ�fCkI�M�W��ԪO�w�q�K�%q�� �OYK��i=+1�+�"��agS�wP[b�z�����t�栊�Iu�97~��x;fj��`Jn��qb4k��WRD��5Sfl��x���AL��s	�+.4�?�����C,&�[!sk���^�?_���N(/��dH��ƛ`����mErk���!(�w�e@.��%��>�E�u��:����e�ͼj��Q��Ο�\�m��r^@�F4My#�������x,�D0��M��e.@@����I�
����_r���k
t ��F��kG�o��8�	�E�^�iT�\01�?8�e���Cy՟`�I�A���T�2�/���oF���C������o�����l��4��럜8B�t#)���iD����p��7	����=%1��4N'��ǀDe2��C�7�����s�j_|O��/ܗ�g�1�J�*��BʽIb(�38i��S�4�lu�
�+����h���K���r�F���n͡[f#,%B7��P����&\��ˀi}On�K���!p�[[og,} ��̇�����ar�'�0j1LdN�H��r�3f$5/�� ������ڎ%��H�s���������8%�p�ݍV�@��3k�N���w�����TgN�U��-�#�m[9����j��Rɧ����M�*i��H�A\���4Z8M�)]��������~�O�����S|��;�?�D�ﰇ��}�F�.�Z�:*��������t�/���vP윉�WT"/�s�0����53�G(
�&����D{-�YƔfE��΀8���'ug!��~���pua�ʩ����,�{�.��\&��N�R��K9VK(���N��D��bA 5�� @��hC$��Pg�Ua���Z
K�Y�"��7b���3�D�_:��֠�I7sn�'�}KM<�,Ј�'��]#����2�	��!��%<��%�E�
�U4�yܪE�r�*���2в�f�i�)sI��P��\u�;�<�F>Xܮ�Y�~���ш��z��X�I�6�N#jQ�}�>tyisQ>/����`+��ZY�����Ǆ��q6�� �#*�NN:(��ٰ>���(C�G�7;��VE�ر���}N���d��e�5��1?��pk�,)y��JX�|@W���];g{�{��@Xu��T�݂��h��5�S|�~�!��΂>���Zw�Ěh�g�ǻ}>��AU���t����O�쇻)������G/�6{�޲ʺO�]��k��/�?XD�``�V�9���e��>)�\�l�3=�4��X�
bw��0���m��{�`vz�iZ���[SϞY-7��g����>CxV;���I-�����G������m��Q{��k#m"wc�f���z�c��4ML��qLf[�e�����7��;.0$C�)ʿuS�j�<�������>sG|�@Tb1�ͽ�k�r\lIZ��Kp�R���V��'�k���<�$�>�g�!���$�d�N���1��Y_~8v$�HYe��h�	�6�X�r�<�P����B��uRr��66�ܮgK�2`y$��փL��,��(Ҡ��fV?$�����%v�J���3̾yj�������|�֕��f�P�ʒV�aU�l��ÿ�����(J����ηY�A��>��1�'�K&l�̪�N0:�C��,�a��+@��4�8<� �,�F ���y�5 6���T�*@:A�����4�W��(�3�?��k�8���)��xj�՞�֡�R�e@�m��7&V�[o,�
B`��QB�0)ڭ�#?�4�a5��n�D�q��V��^9�!V�����G�/������Z-,��R�ǰ��ɫ`Mǧ��r�lM�y�K���x�r��m�q�AM�#�AOF
ʦ�-�WL��@Tք�,���p���%���y
�R"�lp�e�bt�����bb��e k�e���aZ�b�8 ax�������mWHޯ���U������(��D�B)�A�� ?,�x�+91�hoc��;���QU�I��#����9�j5�Nyn�"������)4Q`�EӘ����9�_\(���	���u����y��,�u�����"X�9FهV�_�j$��!s��T�M�zҚ������!,w�y�X���9�@�:\�J9h9�Q��%�P1�\
��{s{?։�X_:�~J��PЧԙG3ӥWpv�4��5ͦc4ӭ֝[�9%�� �>�t��!1�y�bw�+-Ƌ�x�������2��d���64����,����q�Z�-�X�В�༅�V~QÈ�u/x�J&C��}�ө��VN<��l<^����*���N�����1X0y�,*�A�n�I����
w�x�"����0Z:g�ס�n���	BoWm�<�1{��twJk�["`��"&�jB�cM0�p�\e�rƪ�l"0�Ư@��2�"�
�p:�� ��4��D7�:�駻$O� ��I/{>8K��
x��<3f��">��^˧%�����ħ=�<����],�����m�9{JU0�1�zs��>�ޔ#]�Ӿ�e�4���t0v2�S�3~���t��7%����BK����DJ'D]
�K��(�>�h��܉��������Xn 5�ӹg�,m� <u	$�Qbƴb�s�U�W��^�	z����j�{�ITt��V�"�N~�K&S%ح��:�p#�﵈uY
h�O�ͯ�{e�o� ��k����!-�<J�.���Q�BW��K�~��3�^ NQ(,-���8�����(+�-t��,�rk��5�fJ����ڋ����>���x��z�[��E�MV��O�{a�W���e�X�&,�yl�:D������=���볬E�SQY��Ts5���N���~/ƚ�C.����ix;��KO�xy�禲���0�QF�aQ��;��2N.�O"�2������V�j�k����laO���|��H)c��-Q��[ccM�4�c+��q,0��6��_Y�I�g�b�:6"8�(Xb-�m����]t�Y9 �܆>�0��;�*�iv�=�%Ij�s�^t�:5���3�x^l�~�L�>a�Cq��e�,�uď�cȖ�y�ŕ��u�1���:���^�|�d�3�FLݤv�| ����7XC�q�'��?nݸ�֒>,LAYR���~wI��@�M��y]ulr x��*T.�ͷGx]�1 �3������[Hc�v�J�Ҵ�܈ĉ��:�D�� �D����}�pJ��sT�Ʈ�� ^$�r���`zbĚ�Ѹ`��V:����M�ξ�=�ܤ�5똵��L����2���+����]�O����O
0!�� ��������f.>z3�)	�Q1츧r	tw���N9���Jµ�9Gn���lw��5��G��T��)%�Ri��M���u3�8�iG��2�S^�nv	#�H�Y9��6l#Ǣ"���V�,a�C>"�I:�����62$j'���:X���pA�k�*�`�t,!�
/���53@C�S�]�i�a��x�����VRQ@͌��,��R#�R�$u�s�u�Mp8$�a�%	�����U�W��E�7�b�۪1aJ��.�0J���'�1�bMۍ	x �!v&-%_~\UU��b��f,6D�ÍH���QCN��/KU������l3L�.5p=5��1D�;�I����9Q�5(��8�"���=�'	��X�����j�y�|��6�g�F������ ����:Q��t��S�D��?J�81�"��Ԇ�I�B�gŮ�f��r�;Ru`�_M�3�X��x ��,�>�h&D9�x�#�v?��ߣ	�Xh��ta׋p���1B��{{����Ǭ�<�ٲ�?��a�쎔���Aꓲzb<����Vo�m�����I������ok�N�RS|$��Pm�������[ϰ�x�ܜL��͖�5J��U��	�z��!lH(y�b�U�='|�4R;K#�fcP���"�VY��5_�����zp�`uֆ?l,e�>��/���D_�[�K՗,Zw�c�ف�vT���!�~�|L��s��:E�U����i�sm1D�A����G�_�e���9�jJ��5��9o�4�d�S�ޞ���o�{$GM��w14���mFU��%���|�'�л��c����E��a!�=ղ���v렠����V�b��_���2�ᛱ=���!nV�"���c�)!yt�$�����2��4���1/�L���3'?���L�V�ɾr�˶��6�0M8Qj"a��,�]>`.M�"�y��H�
����t<�� \�t�i�$��>y��d�!W��Ҷ�řZaV3��q�(�Z��4��)H�v�!��P�䫗�gz�r���r��{����Z�C�Pu������m2�&��@l_�H�f��H�,7Z��:�%@�(bT�|��6l^*���A6��
�UEZ�V�2���TTw|2JNX��.�H9$kW�	jχ����,nF�e�e��l������c�֕�m���UYh���)�xD���Dn4f=�c��ړ���b��b�U�kQ"��k�>��@�Ԝ�]��������W ��I+e�r"��4��<-H��=R�C֊@쑙�X����7cZ��ce��IU��(k�)�o�iZ)$�1M�[����6�^v �U��z�xnC�h ������@8�!�� ztFZ�^ɮ�+x8��ڲ��E�)���j�)�9QK��؉�y �q�j�:~� �̐Gİ����9/�6Vg��*��"�~~�g슟�y��4��Q�U��x���(�ǳ���Ҥ5ߩ$��i!=�,�[Cv.Kd\���S�0�r���f"��f/,\
m�M��p��m�� �zR��M�Y�z�����+�$�X9?ʵ�4ǨñjjMq轈��Hky*k�g�Q1�G�Vh��.X�����p�X�"tP��l	PN��E��h��r\����<��\����;#��d ��9��D/�*
�}��e��(A6ۡ�ַ+M���p�B0�Gb��gV�Y�aB�z��^S�sT��)�{�/�W�GC��u�����aՄ�Ne!Ĭ��M��:F�K_h�6p��ښ�@���z����&��fh 3P��5��-O���/}��Rl8��Y� �f>��Y�ک01���}�w�j���+%Ҵ�'/lSsO���V�sxO�Q��J_�������Z�t�;��p=�0�c(�	5�>Vi5��T�Рf���2�M5�D.�2�΍	��_%�j~o9?BhA��h��`��A�Nѡz��mj���U=Y����l�W�#��0w������#q韘-C�,i;�^���5�e��4S���y���!.���-�:�-�x��f8�eFu��<��	m��B�6<�O����:�c�W�'�>�w�>�*�g��8
-��e��,�,{���>��!*h�9 �E&�	��wv[�L��G���~�,��>�����_�p5vS8�����폑Z�C�n��	I-YG��b��I��Y�, �O��k��؄��E��S!Bf�E�?��rp�试�#`�s�R�<��x��#��_�(ԔHN��*Z�pX؋��'ՙi�NY��Nu�5�
�"��4���˥�-ҿl�$�-+,�~җ�V�Dв%q3���Ut��R�*���8�nP{��������I�O�q�Y?r/�Ϯ�@�آ��}f@M�d�s�o��qB���5�I�@�eb����.L[���#JW�۸����3���viP�q��Ze�������ڧ_)�gŚ�l�M��0ޝl�i`�,Yߠ�ԗ;�~�d�l�5�7_Y,��Nj�V�l#�0�1ON�����Vlu��I��'�P1��E�8�W(��E�����Y뮀}�\X� �ië�T^�Q�9D�ZK��d����H��b5�ۏ嫬P�b�y��JQ��b�h�.��2~Α2�9�pmXQ��K?����"�ܶf�>�_�n\	�����Q�!�Ō��t�Q�����#�3�6����4�m�m����2��f3 �L�P�/��f�l�2
E �$�(aQ���u"� ��V�V��"�dտ��F�&?#��1w�a�쟗R��LXz��ֽ�9?QGf��,5����=�o�N9�Z�"w��neE�̗�@:'a5(�۶�@�֯|��A0�d1"�3NR�z�0��8 �u좫�A�� �k�z��Q溋�.�IF�x�
�k�)q�xI%��#�`IL�?Q^�;y��,(����������w�u��e����ǚ&��-("��\��w/�mߠ��޷�g2�m�v�����S�;4�69c�߽��MvbL��?U^�����I���/W�t.wl�
�PM:��������ҏ��,�0����� �]Ax�E�i$��W�H%���匰g>��y;�I�)r�?!��};��w��$j��1ӦF:�>E��kI�U�O��I�l9#��Lb�_{��W|2~��q�r|�J�A"�u"�A��k�lMI>��E}]>�aE�����!�<��@�2�%�Sz��H)�1�혢�~e�~���@��=��ؒ�6���BqZ_��,�lM�Pd�x�D�q}�%��`�)g�Pu�3�*';�8)��s���*�!tQl�jD� �S�����6�gk,L꥚�^.Uv��J�� ���Ёt�/S^�QG�(���I���)��j��=TM�{to�y:�Z�B7r�Zt0�վ�8��T%
�!�o�j���v	�tW9$��p'en���2��şԟ�0y��O%�J�-�o���@��]0��)�5�(���k�:j�� �}�R��=�'���خŇ��;�1Ȅ�A�`_������!*x�Sδ5��B�o	���T��8���x_��1<�c��h}���u�1ZR�K!������V��h��Q��ދf��R��3����K��)���eH$2V\�`�Y}n���S��q�n�b�%��xA�ne�f������o�8"�h�{�����͟9�oD@�e�/S��0E`{�rZ2
H6%*�:2�<�9�8����?���9��3�ⶥ�0�g�Z�@��|��xb�x �l�f\Q[]��N�3�[;=*��)�G�Ud{?������`�6�ٹ�ֵ=�7�-r/TM�hL~Dy8�T(Ps�fy�-�e�Лg+��o{�
OV�;D ԉx��(�C���m�co��ͩo�-�Q#kc�͹���<Y���aׁ�-f�.��WH[,U�<�n��Huy�b~e����	�+{�@���j�\���LJ��w哟Ӿ
�����D�etz-�F�H/]��x>z�ܤ�sV�)Q�Ü;�����DL�^%�4w͙S�Q[�dߎ� =�J� ��#�i#�t�P:E���hb�Y�e y��6��O̳����0���ݴ*:9#}<R����xE����gc��}�ȳ�E
�������f����1"��{��KbTxA�?������彜���ʂz\���O��֋��"�����_Ig~~#i�g[g Z�ˍ�௾FU�n�ma���@���P�Q| rǮT�Ao�)��-�!Ҿ����&����J�]ZV�^�&U!@˝$���ï���l����y�N��T6����u�8Y�k3��o�h�&��hJ��d>$���.(�(XJ��&�+yL��׏�6���TP/]��f�S����1��T�>.)�>u@ۥ8f`�
E�����y�}�ᔮo���y��b��
�}��A�+bY!� },�h`��fÊ��fypb��@w�wVu�2���gL�(壵 \�e�)>�n�%Ɏ2u���Ȕ�8�7=�t�?��o�6�(� #�ӁFa��$E��]�����5ʞ_  O���	��4��VI�uY��EJ�Q?�Õ�5����t���N<��B}t���� WC�<��}^ii��ʗ1��YU@�	7v6�Jta�5��6�:Zj�ä(�.N6�`s�k�j�
��������1�=� MVP��D�s�񗉭p
r�U��f��Dl���g�[t@�2�Y����n��V���_:�b�������إ�@D�i7�� �����D�W(%2����hN�P��n���tC�E*���6m`�f�4}G��r�_\,'?��L.��xYr0�fB6�#�(f3ك�Z>?J���N-SG�iT/9�s�b��d��M D[���'$�M&�bor�l5jA����	���]G��4�~3�R����7��53+�e3k5��Q�g��gϝ89Rw��k7i�~b@$$�����l�J��_Q[l_���ğ/�v��y�������Oy"�̌%UI��<���}wz5���p��q�D�Иv��/@%���s�{���4�j�?�Ts�����*(9�~?-A����g��_� K��rv����U�c��QH���8j���M!O��=���!QDDҚ\Q��4e��S	#�at�R�`>���[����g��j��r�˱�Vȃ�{q����칋<���D�J���?]y{����D�q���9�GC&{�31L�v����N�c�%1Ci�t��zԧ���ߠ��t-�r�� �3��W�����7�NO l�ި=�n�2u,s�b�~��|�^U��m�!\1j�+7��>ER��{g��5�����[1Ѝa�8$��rJ����5!շ_�ڇ���j�j<��pg_�2K�;�Qxpl?�)�����Wz�l��@�;�^�Z�uf��)iL�գ�{G�%���s��,���6@�)�u�̏�s����$LY?;q�n�~�"h���7�5��wa���U'���Yş�n�/zϦ�gC��ҽ����s�����;���#����Hg��CѪ�WcU�G�����p�a�!�׫��@�����j(�[QR�[�
a��� �P�u`�������x"�]��u|%�Bs�Z�����U�����7jL�K�!1�ּ�ל}^b{ƍhc�սĖ�0��/����U�	�[�o�\�$�&&M��{��l��i��@���[��M)FNK��=n]�	��8CgI?�j۲�W0T���wgɂY��y�*I�c���z���{����I�y�F�*���`�I���j� Cn�A˃v6��\�����fW��a��@��02�}�{���Q�:v��Z��ģ�X<�bG���u�v���"�.��U��K�N�[|���n�덜�uM�u���S�l�Z���;y���}�'���by#�ґ���G<ϕ�+P<r����p� �����0|]t�#C�ε���!B�y���O}j���:�k-�a�֍�	%�p��-��)���γ3%dk�8$�uK.
��f8��0�@�9��2���k���ys5z���amp�S���t���fg�O9:��sDV�����Ó\�[����N�`}����	�&�(F�[K� �(�%�ɒ&q�k��ĳ��-���5Xc*_�f�I��Is8�I<��gE!񜱞�XhƵ���F�U��� �v��jYl���+xPK�6,�\�)C�)���x>�����߇�i����VhKp�͋!$b�撖5i�F&j v���n�6Wn �b��oH��Q��$ �B�$�X�mu0P�����x%�wE-U[�O׹�����S/�!9��&Z�^��D�)�0��:�u��_�{m�짟3S��j+N!ǚ�R4*P`f�kO+�lwS�-��*���X����dxp���E���~���k�Q�1�)I���0�,�a�t�Rvaঽ+2yB���%x�3
���!�9�S:��BF�(U�:�2�v�œ�m,�^�]%���)YQ�ӧ��S�ܶ��1�.�쉮h�a>��o��
�Ci��B�^z���񒣭�Ӟ�p	�=s^l���9	�.P�IF��J?�a�1�?��Mim���S�-�[hׂPV��|)3:�M���V2���Ӻ"�-h��ִ�v��{��K��/X���1آh�F�G�Xoj�Z5ڲ �d�%�f']�1�RJ
MD�u�4�ņ���W4�U������p��յ,�)t8 �CO�b��6�=9�d6IщC	��_�l�	�Ż�G|bF1m�"�4}�[ s7������39�|�䶳R+�{�;+�H�Hs1����S#�k�`/���YvE~�H��ܗ�ա���KG^B��46Y&�<iT˛����M���Y/3��0�$}ʲ	�D��Y���N*��J�%�+��r �i�)��<KbZ��q�Iҩ�R/g�lW�C�8I������ƅ[�����ٮ����n�Z0]�򻂡�*����~�z�1Z�x���wM3N�����lEkdn8��qȣ_�'�w���M*��@B*�;�r�A7[C�
k5�fL"��s�;S4��8�����l'|;U�@��#*p��j:�ʦ�� G��^�ŏ��(1�Mf��үgT�u8��h"�cp���5�E�:$uY�q^%�b.S�H��ۼ�� ��2/g��Qv��ܶ!�?hU���0=����,�M�l!�������~$�K�%/ϣ��@G9՟��2��k��){pѫ(0�N%�R�L�>��/�9NǑ��i�l�w���`u�krZe���R	��T�ꅣx[j�1QJ.s��[�7��ï��V^�=ETJ ����B�7��h0[1��i���<=�Ru<�Yr���M��.	ot��������Q����zx���kb=�9��$I�y��y ��f(G��N��?R��]�Ds���j���#���J�ٶ��M�_��,<�ݖ�C/�KY��E��RțՊ�P�.�\��hHI\�ºs�b^Q>�̭B�N��ر0ƉCZ!�E�G�	�>���8���D����~!�U�e�䜄RVr��ơH�\4�`8U��g��+��Lu@�7�reby�w���R_4lB���jD����R���?�-�)諸�\	^b�q7�j�9Ir�*i".Ȭ�J�����c��P��_� ��;=��IBq�,0��8�L��kI�Fx�<>/oN��߶�j�����W���YX܃J�	�j'�-3���2w���ߘV�������Pś�l�j
�U�0K�]�q������r�pݒqS��x�V5� �H?��6FROӕ�����C���K�c�[�1d���~HO�"j���6~b��!�D7�]{��XX2�W/Tg��:���GO�F�'^�iL���7Pe�"A�e��Jb�4��n/�e� ���T����fCc�|ؽz�݁�`�ص�4ٿm���m0�����V*��t-z��"K1�Oc�Ǝ�XŐ7��3�=`r��G�.�Ğ!��bI4���ՙn�W���)�N��� Pb��̲��v��B����T�&1dP��_��M؋�J$�7О�x+p��0.Q!÷A-�
������1��oK��T;�G���_c��#)�`��Z��&���H����0!�_� ��g�D�l����ֿFþ zL��H/Td��;�"�?\r���麟Zk���Kwӿ��D��L�?t4!F���"7���C����)�@VqDݻ���Ȳ;1*b0w(U�[����,(ťB0#~�)¡�#|o�1�y0����[�Q�n�{2+j�r�y~���{Ҙ�d��)�Z&���>��IsH�m��]oW�AG�� ���!���&��c\n���:�n�����
{8j�?}��g��*"���@��ra�랞Z-=�b]CP�U�-%�@�mB��RTl.��nY�ގ�=��:ܽA}������{sw̦�~k�T��ƍ2�k��z�^�w�UD�"`�o����]�1M�'��P0�M�9�P�!P�a9gͅ>���բCÈ+xv�Z��4��uAQ�L��] o]s��&�%�>Ы����7�jA��Zq��*���x�ٛ��u�Ć�%k����d�JXs,"�J�T�E�u�g1���{�yخ�@��O��锁�)�����p�o��(��H�k�����b���I�"�)��z�3�)h\Q�
�t��(n�c9&��0a����lb�#Nի� �ڦ�kh���h���6���	_��#�A=0��;`#d�ɟ�ai��+����20���o��ɓ�^�=��Bp��U��3c�����х�����ؾ4�l��6�����9������]����-��Q��4%]���L̰�
ڹfso6{�Nt8q�7�:CL�h�iM��>ɔ���ur�����J�n/���#bx��;�_яl���v�9����"!�u��e��#�E^c�"a}�>U���T)�@cV��#\
��Y*��n�5��
Ê��&!�D�`:%�C��:�����8<����9�xx�,�¯q�Æ���Xm�vO6&�����3��hS=<�W�?,޴a8Ioq8�cC�+���\0�[�>��)\�B�
�# �$W'�5�M,*$֧�8�Ӟ�9T�X��B%]��,�� �y�hg��^���Y��ՖH)�}�G4{~�>z,B��g2eD�7���y�C�+r�
���)��4��Ѡl�$��Z���g��P�eݽU���>Q>������J�)M�\;9x����h�����Ԙ��j�����K2�[�]ͤ�M���\�������'��VK2h��b��Ee�g��-��=N���Vy65�/��� *��&�Q>�mɔ2���D�9��m�D:�N
�7+CK�o��c��&����ʢO@�͵|j��Q�[ .��	��SY�n��K��4�J�n]@���z�\�l!�CM�$�1���^6@׍��B+����B5�4���)�T~F��8��a4���됣_!���� Q��f��T+��Կ�.�-t�lƗ�	��c��M�ed���"�q��G��҆j[�S���{����,����3���S��{]#�V� l�b�Ͳ���r)!��U�`S.���.2�d���E���.�2h�a����,#t��Tj��U]#��o{R2Y2a���b��ʱ������'��5������o{�����sQQ%��.'e�g�a�ST�:|�����dzQ�l`�	�� ��(�'jw�o�T��~_Y<q���^��^bS�k��_���.ҝi�)��fVT ����<ؠ���^A��Wd)�X���;��_�A���h����?�Y[yn�9>E���R?��ٽ"�`i�O݁ŕ�)�|�+~�A/���0���> �����T�F�q�D�*c���nk�s4�w]��5�( C��V~td���eY�%�9q�0�n2��C6�D��!��K:D���A q����%l6�x�j'I-H��~"C��2�u�+R&�Qb�Y�u�ǆU�ꭇ&���(�W�<3�~�����Gm>\�v�2 ��,훭+\P�zy�E��>���.F�������\�H~3[}�c�<��5[fڎ��!��Aq�$�uq.y��<%դ�Ov�9`���������|(4bg��~J�:@�l�p:�vk� �X���'���w#CkJyX��L��3�J�[c̫���n�+����>5�;��V�L�H̦�䡅ר�W+�����KF5E�b�ּ�3�<�g��y�`�K�s�6J��:���fR:/����6|�jDw�+���^1�hz�'��ѐ�iOBƴ�noT=��	Ƹ!����,�0��Ib>yAz��\�&�dWR&�	�Ő-\s̪����v�U���X�NND���u���<vP/�����.�.�����g9��j��k�^��*|KyKC�$ȅ�t]��yT��Z1�ݩ٨�(�ĉ��n��F��0D+�Ɔ���x�ڴZ` �K�AG292Q���](��q^��ˁU�45���1-���[�x�s�oS��AV/��� 2�;���6�(���xnp2鱢wm�o(��$����X�wS�3�I����+��3`X�%�[[9a��Dv8��`�/ޚ��1�Kl-�-#(�P�uj�-�."�?��ô�X��9��B�7��"��f��
	<:�Î���5��r$��F�ہd��3�3zؠ!�jeꜬ3���\��c��Ϛ//��I�ꒂV�'2	����:���Ů]J��d�_��;�{F��k.rb���$�	>�>�٩Ziǫ���wT#��J�i�)�nr$tKE}i�U����UbjN�C�t���2b4��e r���jQ����X��[��`��2�ڎ�d�0��{c�k`l�:J=�iû�.��m8��.n5<K�yɞ�4h���ϝ2�' o��Q�?R�HO�ɽ���5=3(��ޛsG����|ᵴ9� ��[G��z�s�5�k����?Z�ΙMM��zTv3d�M%prp�a�Zx�GPQX5J����G8�ڦ�L�QVXs��=�ۣc��<�F^9zf��Y�D=i�Ҹ����;5�cj�GR�0#xd�1�r\�H�ue��&�-����Xw�T�$I���l�[��8v9\G�+D"�&τ�@��}��Q�"�;��~�f
�?-�G�9���ʝl螩T��+��N��Ӊ�8��jƂ)�b.�d���[�*A�����9:����ή_LIB/Z*p�pz��|�*�k��t�ik�+G�q39�6�@�ᩒv���ϣy��!�6h�=�W���ˀ��f�$�t��Qd�6[��wh�* :����Gs�HE"Y� �2?_qh7G
�O�?+�I�?S �̠Y:@t�	��n�"Y����Tm0�)x�>}8Z;�ơQ謷��08!��."��ۺ�>�8!�bլc��8�l�D��=�>�x���TUp ���C�I�~oQ��0Q�YG�|����HA�
c�ɉ`:d �P������;�����U�<}e2�zn1n��N��}�zO
qų3ݩ��s��|5���)e+-;'������#�>�ؐ�{="�b�,���I���3�s��<�>T�3�"(a �
��j��e?��yt�6��k�¾D�A��a��TN@���`��ƒ:�(a)�8:u��+�d���qry��EA�h�ǞU:W/d�E�W7��X��rɁ:�Q������KTxk@�!�1����-7 ���ۜ��uc������%�a��P��@|}���U٧�}��O�T��N��=a�a����/�@h_��e���R뽗�w(l��57�5�ܯ �R��Q���ݥvq�m��_j�U@sɗ���zB|TOd�>�/ԩ����F�!s�/��.��W-�k�$n�A^#�;��1Ug�Ǘ�'39W�A+�Zj���o�}+`2�Ԩb����{�i<��s��+�N�����<����и*{"'B�`Zū�
8�%���Kbޠ�[D���O�W�x�C!��6[|!�Ũ�l{��Op�ٗB��զm 쓶��������e�/����2F�?�iAj�L}Z���LM�	��N����5�7��V!y��+��QL{����ץ����������M�(��$�3X�dN����ڈ·�">�B,���$�$%����$�a#S:ӁVuO^ܗD����ӗHs|��yw��1��O�����8��[$��j6A�S������@B��u=o���&eY�)�%V*Ê袖�$�I�LrN&��_�{Nz�;�tb}��+�8A� �ݮ����vm�
�ǯ� C�!�0x�r��Y5^Q��$�眧#"��.��L�%����ڦ��b�!�G5;o�w�BE兖,�lA)�)�A�E~�P����\�w��@�y����J�B#���L�e'!&�Z�ׂ��f�4O:E�L��u�M�?�c��71PJ�5YD��eYl[oR����(�3�w�y5��p�����q
?09�L�GU|f� �׸:���g�$T�۵d7��W�t�~�s69e.57��̦�["?u���~�X&Bϰ��J�F��6$�����[mB�����N�9��Ğx@�0w�����h�D{I�J!��ڌ�I���R&7�^�=ŊVf�M���z���:�J�#�#:цw��~!96)�<���瑻Zsz���_`�it(s�b�=���+1��牷�e�*��R:0�r�8 ��f��RE1������кō1@g.q<��p�ߢ}w'�SB:�]��M�i�ϾZ�w�H5�.�$$����
Q(���-��
r���1�V�6g�a�v>f�P��I%#0���V�Rc�a㦱�;Sba�`n	U����A�5|&�v�����%]M��]��9����_�֥���%6���/v�#��b`]s�r���[�Ug�!�穵�"�Crv���=���4���k+���(�5	���Q�M�ؐK��4���4 �!�Te�dX��'��}FY�#�t�{��2�����E+b�8�L�i=h٧'.�mf���������X����öby�ri�AEwr�oV����s���F}���@<n�����l���>�6İ�oO�ouȈ��Z�;��\���䛌>�����h�+B􀞢���zH*��h���"{-Hӝ��w?7�[I�[E���V� �a�� �W�0'�[KgI�VLi��I�t��	V��z�CI�ǧf�dF�/��/�/$����-��Fn��'��gmZ��$�\��7�t��B^�@����	S4;:"���x�a+U*镭}=?�grAXP�Qt.�-?�H����O�Q���i�N��j�`�*��s�g���PL��H��ӆ�A�3ޗ�GKq��T����e�s��Xd��?������)�H��5,)I�;�<�ٳ�
`4�y��a�,|�g��1�Q��nv�?��n~w�iJ��3'HV����95o7"������'@G"X2u��DSƙX?ބ��%�B�렗�Ѳ��L�N@�ڑ	��lO�
��GҎM���?�d�D��t���A�Z���G���L'%x��K=ef�=�R�6$���8�������Њ�0z�!�����+%����{)�m�_��A%�p����qR�(���~�+�r-Fk�] �O��2���������w��;O�m ���A�Ķo$�0��2�Tn�L�I�=�5�ވ r�?
S��#���B�BέIp��Id܌/�ؿ��~��3G`�;Cn��JDL��༨O
`r�c�.a�8�
�~�*�9�2K<�8��72��Nt��7�+�����{%0ԝ�9�%	X7c����������D^���[�{BS�|D�
��|̮��R4S.^�����giT>j�󾏺�o�����*��'͵:��؟H�CEՙ�p�\��
�.taM"@���6����;��N�82�q��'��@�U�PK�by���ܷؑ��y�$��L}�'�<�8�Ӡ��P�l�Nt�aK��xp*���K6�6ֱ�18��8�C4)ȑ�[T<qr'G����yS �3Nx&y�Vc�Ƙ>���Y��P�7���&���	wރ��lz�+K�+c
Q|ϻ��a�!�ŇVdJC�+��10WPqm,��BP0`��ɟ^�'\��e�p,ܙ�g��G��|��<K�$�$^�?"����� _'fGL�_ZR���8�E�т9�I���V��i瀓�N!�˄ݫ!i�+ژxH6�d���S�t)S�[A����s���iO	��.�,
�{��4��y�H���~�O7H�Nv!�v�]Q�'p֊_�ȭ�mʒ�'�i/I�LE��utY���f(����1؂0����e��2u���K	G2�g��x�|�R�����s�HUw��V�=h��&����];A�
�� �7�ɜ�|$l�W�	�� �P�g�-�I�gSǲ��^�ꃜw�1f��[uG0��Y��G��ں0f�,^T�d��QE
��qw��&��n%���v�B��k�2-�[*E�@ݕ1�|��L</�����F��$a�����&���>p����r�ʪ7�+��m9�<<�{�b���0�3�4��QT����Z6������}���$�q@��*��QM�c����}��z�7�A�L1��}�$���E��,�9���r�����S�B��Crh�Q�2J�Vzn��mv��<�fe8כ'�>ۂ��CU���-78�9�2&Ƅ���ݵו��L1��N��*m��i��W���ֲ�)N��vv��}>�����o�ܑ�K�*v=3E}N�&�_j.�HLz�as%�S���^,}Zz̰):k������Xl��派��z&�o�wce6bڽ��f�P��Om���R�d�}�I��h���Cģ5��q����L���j!�8J�7{�ʅ�2��O3M9�<��M�^B�
k�%ꝝ��g�[�e`��x�-
�g���oĵ�!����n|ci���O�%@����+�~���۬�I�8wE�y��a�D�h*�%9Y�����i���*g큪�b�ZA�xz�f����j��7	Y��S4�D�q���B��!!�K�j�q=�_�!=�zh �~>���'E�M��z��ց�<f�x�ڿ�G~j���\U�@�:}"� > �T�����9ؗ�N���g��Odd�+�Z�䯤��"4˵ՎR�Ƞ��L������A�9'�3?70�(KN����`����4���ߜ�J���B�܍�u��\�6 u�B��o��:\B���1R6�@�ћ��7]�M�;��S�Ϟ��(4��9�O:n��v���B� ����,N��K(h�:D�#ÖI��W���t��[��,�d����`(�ȴ+w�\Z� �z����G
��=(M8��+����;��I1HS�I	�$`Gb�e���i�5�l���%ړ���ڕ�JL�y� ��% �-�]�r�ׁ��~+���{B���dh��Z��_`�[��ĚB*�K"�	���r>�\X� ���k)�Gl� �/���Ҧe`��=
�<o���{rt=�����[h��(Z'9 `]�����c���o���X�����wp�����{������<�����X*��֙��f���ņ3&Z�p�/5�Q�Q�)|��IЗx�g�4B��A���P����V���pFZF�*P���ܕ���;�QeȲ�
�5�Q���)���^2ew�މ��7D����`��"�x(�N�ԽG�g� ����h�)�d�������c?��PsU�G�[x�?��6U-���ڔ{��)��(��G`D5:���P�AO�ww�2��	����>��"ͱ��Cg�P��NXZP���ÊLZ@�(�7B��0�,�.3��oQ״	���jj�H�ֱJ?�O�E�Ra{/#8�%.�<�v�s]n\���ǋ��ד�^G��]G����q�Ѻ,Ot*k�����B���b��4�<D�D��t��w��bX��n<��o(<� ���ќ�\���f��bJ�H��힕�L��{�n�_���J�E]n�C��/$��ԡ�)@Ԭk� !�ށ[8���O �=�zu�]}�tꚩ��t��� 4�����g  �f����~#�P*�=2MM�b.��=��<��c�H�P�
��D���%�����	h����O˼<a�ƿ��n�� ,W�v�t�Kw��T#���#�	��[�ք��������-O�>����:�<	J��������n��������
�Kj��jObo)� ��R��h�i����dL3��`E���@p�s��]e
�o�^'�����ș�yB�F�$�bt�Jy�����k[�-6Ḝ-�u���	��/��R�Q��?]�-��g��mVS�f�M�ww�^�U�N��ŏ��������>W�z��<�|���il�ᰶt*��6�C���i��vm]��^��E{|���{�fB��ݵ�U�F�:����\�.u�f<Xd�ҽ"]�5T���/n.�����<Cp���J�����x��;�~�s�J�$i�p-��ȕ/���B�"h��?S� �[I��[=�<0-�v(�BGRd�=%#�T��a�_O��>�kKv�}'E��ʩ�L��w��6��@�ƽj��~.�@�bQ��f��շ�����5�odA���|�օ��]T� �!��F�>n	J��k�`{��teD>�%Q�B[�b��{
�v�pPs�-�<����ftp��L�:�Qō�Ctc�3UZ���5����O?,��5�Ծfr��>6�w�2�� n׫��R ]'��O��U�Z��{���Qh����2�c��}���KN�s�+�H�>��F������d�o*z�]8N�ׁ�x��n��$�W8K
8A-ި����8�d|Wd!��G�f����kLh%V��ϴ���\���ܳIz��4�O�ӀL��Y�̐4�J
V�~9�ox���ʜY�:e����;�ǻ�,P�}8D�(O��(\�	�ł8ג1�4k��,o�߰i�~J���iR�(]�2��ʮ�O�L�jb��0Oص�s �IV/�6�}ʈ���0�����s�dl�I?<��b��{��<&�oX�j)pʜWƇi�����U8j*����]`�Ln���D�6a�����:�}�@~4���3�xX'^��&�V��xf:�L=�7_�  n��O{ŀz@AB��{ɏڱ�G�V��wj]o���Gk�-x�ox�1	�h�6����$8����z�r4�ϼc��a���DQ@�*����� ��;nb�+�J�����y~���:"���9�_#��O��p�b,= 	Pw�v�w�~�wx�d��;#�!���S���@�^�.�������w�eφ�d��+��Q��"0���$��ST7�,�>m �rHY!Ø&� ӔLbL��#1��{��,����ܼ��.$��2^Xh��u�2�P7}?2Į��{$.�	(��N�GW>s��'�ԓ�ě�`Ep=&d�L�܈�I�Boo�	6�����F��Mw���F@�]{$�>��߸?����#���zJfOH���5u��&o`q�1�����+�Eg�(���aϰ$�@���#�g_F9�{_>F�/P�Z�$�MV��9�[j�wL�Y�n8to݄L�
�F�8�m��X���H�@ ��P�O�i�O�/KF����d�E��� ��b.^�Oǐ�:��kW��,��]IZF��Pc_.����w@
��8��K�ck)�|KY�����S��w�=��d�]���ꥍq/x F3\=��Qn�s��ь{ސ`�Ƿ�Tu]�)�@�$���<�5Ʒ(���6Z�D_Yp�ZA���u�I=
 -FPc[4&>�M�uK.Ȕg�"���VP>��:�sᴫq�J�G�X�'�Ɏ���Wg	׉�9'��uq`�v�_58��ڄ�|��&��[�(�#��z���.��6��#2#����`A`�ܢ\$b�9/����	��F��~��G�z�AQ���a�F�awR!sO��qJ�l$�6͖`&�s��J�2��oқcz��84���j�;߹鸥o��M2�.]��B�J?�O��F[���(�ӣm*Є8�A��� 6�g��J���+L���}��7:�s��+�r�N���/��˿B���ܦ�A5ñ�����Y�>�1P��Fv�0�Jx<-	�o�`�j�mY"x�����>�yk�����]!��g�i����E����Hx�:�M�a��k`��ԝ�{�V�p�����u��I��y7�{;�5������0��$ӵi&��k	� �����c �	T�"��K����h���Ή �9F7^��l����a$t1���4]���4�#oDp�Gm��� �Y;�s<�����d�zD\ F$t���/� "��B7�-v��sd���j��B���z�V��P�+U��a�GK�Oe)7��0��5	2��6p�֬)��v˰3�;;������.������9��[x%":� 3�V ?��U��E���_��P�!���A|kP
R�G%0�e$�\z$icf]д�Z5��#\b|�}��%"R8F�|�r��o�����l7I<���D �v����Q��)����`��?���|�Z�z�G�AL�/�ݖ4�A��Ό�5&tG��r��tΈ��"�Y�w?dMG�$��{����+���X�����Q�_���s�+��)g],Ա�/�?�ыE����5��>���l}kē��	.�&��6�ކ��a;�#k�,���ê:���m�%Jn^���`!�*� ���xD����i����A��8:�"��i�E�C��q���U{c�7�p���?�� )��C�#���� u�o��Ȉ�\�My\�%��EJ�������J��V;�/��A��~� �+�:,�6t/u�$
�''>*���9.�MT��|
���-�%�ʿ�rvi%#��m9��Re!�S�pφq�Qa���e�{o�OM7C�~\��B��-=�|r<�i�攼���c�$Wx�׋�����AzR��ظ��X:��R:@ן�#��J[ɀZ���	�D�	<�j\�!,���n~�ag҆�?F������H��(Μ.�O�v����ɳ�G�2�������ؒ|�rӬZT�� �R߇]���;�Cq˅��Pw"�|�o3�|��7�3�h��M�]=IT2_v���@HT0^��u���l��X���Q�n4�@����9ea�/��oN ��(��cc�E@�u���>cQ�U���4~q��u��� ���-7��C��O�w�Ү�He�q����Lz���[�����3.��tP�����ڃ����vء�eSE�<G�+7�2��䬍��ռ���7ַ��^Ϥ���zId��s�n���`*WM\�_�1���d���$�Fv���X%�%�$b_U]��m�Ek�	���Q6�q{���ω�+������6gH�c�)S�R2�#���6��&�ii^VA>a�!]�w|A�|R����If�D/`��o:øF��腯f,�+���\^7�s��F�M2q�-/��G�Ib �,��������h@WK��K_ݚ��5���l**)Y�r�A���$�Ry4��k�r��|4�M�NfJ���S]'�'�d-l�}@��9u�+'�z�OM0�k>U�vJ㈊t���N����5��!���K�y%C��l�=-�Q�&�}шl���[u��X"�0d_$�3+H�cC?TP�*"��1����qN�`,�mP޼Z:���޵��D�ʔ��p�(��2�l��fi�SzN����7N��tr�>O�A|3�GӰ�,���0Ŷh��`��9�� i�%QH�*R~8ID���sI$i���tp��c�U`�>_Q��ь������t^�g@WJd�X]^�x�;7��٨u���O���&��rG�X���p��|#3$�������R3�w	k���	8�6�����;zE��fe�F�$���0YU�䪒�����	!+�<��3[4o.I:�:���p�v�P����N�Zv���U�ɡ]���� ��[����ﶚ�g�v�em b9k�C��t\E��1HyUl�+�_b���4 0[$�vן���:O�xS���>�{�����'h���k�e�5WLh�s5q�NY-E]i1���@�I��>5�E͘]����m��!�=ʖ��5�G��P��i��1ji-='.G1�G��EnGb�FQՄ�e�G� ���u�/(��1TH2����xh���#�M�c��_�^疣�d,�O���9 �G��=��r��������8bK�o�_������y�0:.%��`��=�u�6����{=;U��{�C,$�iU�0u�\b�3d%q�-
�_2�0��!u���Î�lw��in���%��֛��౳���
.���T$��F p� ��F|�S�OB��/z?"���u2WlL}��G)����9��=��Ao���7���Q�3��ݔ��ғ��(E�ˈ�#�����Z"}�^D�z����ɪ�t'��;&�������s 1D8I�0*!Yp��p��x�FJ�K�Z�f뱉H�p8W"�gѫ����+�>s���o����������KTO�w�W ugW�9�+���[]�k���Ӌ4���o[�P�WV�zU&��R1N}:����xfXYL��s��?j�2�/!1D��2�n	�q�Ȟ]�+1�vȣEđ���n&<3��1YW��Tn̇�3���bK^����Q�m@{63/���5�l����Mԋ&�1C��W~8$?��K�aXC�-ѐs텩_�es�3��=�����B�z�%[l��q4�?��T�4�H�}��஧b��aF�j���w�X�*>�%o-=�~�X:ոW� �}�j��גs=z��!����e�lF1��'�9P����� ̷-֦77�	JD�}7�x�N-���f1���*LO���� *	�@T��ٿvךn6wW�r�8�����o�M�Q�-:�9>	e_�Vf�&fi��� 3��AI�j�@VDk�;XEiV��$s77�ۜ����"{��e}�<rr$�7I�T��O`�R�b��`����v� FzULD�
OW�0�ђ���]����'���l��{ �d�!d�YO�N	�H����}�Ä�=�)^���ǚ��b^7�s���XPJ��5����cگ�;���=[� G�)�Q�':8�{t���{�d��LنD�G|�Y]�o�"n+�O�
�"P�^�z\b��X���Mt��c�BdW$�E(<y�fqG[g��y/��f�5\׋�fwPL'K>|�!s=R��\1$���~<߰[ �m>C+��i��)Y�!�I<�}0͂���}t��R�0b��$R��+EF��k����?�'n9�m�@���)�n��F��	l�>����@W���+�lx]���~,z�l��!*�2�ט?���qD~G/֕�nUX����wi�̛��y�j���lh_`I��J6]C���N,�����,�%ݗ�p�mu�ƫ�;��9��D⦀�P�KIgsj����+ض.1�Ы8*-��?�3
�lPevmm���Ҡ5�'4��⡬��y��m��fFf�G�i"m�~�z�Q�b� #��"�Tz�Mp�|nq|�H�OaV�Ӊ������>�ltآ�@OL������Kp�B�%`8ISxG�%N0��o�w^��1�`�T{�r��\g\� �����PB�^��b�Ԥ2��fk*k��,��_�M�T��n��8F��3-��(�+�ф������ᨘ�8@�/S\�XH���� 4BVK9�gO����]�]�FF��g5�*1�$ ]6��;X���8��Ey�����`P���^����H��.Jv��q�JM�2���!r�&�ܺ��Vˑ�V���0+
Z��Pt�U�WT�Dp�y�#��x9љ��S�o��Y0���.�G�Z��ǧ�ȖR�W��p6{]��: E���/3���dM�չ��8�.��DW�%�H�h�p�,�L�\�K;����Gqg�g��B<n�����&�/���\�oGj�)���`�gΜ�'���'�A��fjft�	w��c����L�o�%��ʔ���Wg���������L�a^�,���Q�|���mH3�ąl�@���fg��##>��Wy�PzK8T���$�@J41�Ձ�D'�5?�sp��6���*��aƴ߷rjV��Y/z����nh(JI+Ƒ��/1�@��F�q	�N�o�.��X ��S9T�'�Ƙ�D�X�;};8;� }e�>~}a {K�Z�Ɯo��u���� ຳi1��(�~=��W��lF�i����v�+�e^]���Q:.T�P���I����cc���� ��fͥ�e�|�2���Pѻ7�\8h�S�ū���$����v������Ģu���x�|�?�ק��o`= 絆Ej�|�k��b���-cyF��E��7�Rp�#ٴ2dX�P�|�x��v�����]�>�n\����<`��U�Zf�}���.7��|z$o�I_�z�CE89�>~rmC��;���#��c~_r��|f�dIC<5����kd�B@pǣu��js�A��!�i�/�gHuf��9�����j��.S��i�.S�������?��wF���yϓ���=ME��b��e|��s�V��N�t����^.�\�����G�7�2���'�V��P;�K�(U�t���eF�^�!b8=��4)��Ɨ��*J1�u���$�"�+�i��&t]z��@嘐���E�p�����s������F~�R�������+�	�� j�q$���K�G
�)�(�i����.u�Ý��Q �Λ��Ǝ����T�=�Pݑ%���|����3V#L����H n	�6��C���~��c�M&wo��������fK?zό���
5?O��f?�W��#|������bB��ڳB����A���gS^�!e�W~�s�9��X%��r����W+@g!)�oD����yO�B�[�d\4;6W����,���������Z�S�=/ ���\	���+����^��Oh8F��_��r�e��:���?� D!�+�o����'3�1��)0?�6�jV�&ɰ�<J�y���>�<v �g��c��&*�Lw�+-ī�7J��B<�4�苚�,3,'�Vj�t�� :� �>����s��2 ��+��>KPӊ,�Y���3���/���چ:�Vo�K��r_g�J�fX�������"YKE��BJ�[�D��FQSW��&DM��U�R/:�7~$��g�1�'*�ҷ~�2t�BoB������|�M ����o�Tb��H�|��h' A���G����4���<N�1h�{[m�
�2��,�/�<�����,7wq+$"����7�^��R�
���,ށGϸ�La��g�Iܣ�ф�I?����w�+�J����k��F/�	�ܛ�k��z�P����E5~i��2z�@��I��?��^s��sV<#����xO��+|��ċ�^�E�`	;?�Anڨ�H,j�Z�������`a������o�� 靈���k�/ڀ� fz�6�}4I��
Ϧ��#������k_7}�ȣ�ܖ꨿��H2�3�d�Z���1?���[�t�Qҽ��F��4�q֑\�)k����Z��c�I�f'M�\ѿ���+;��*˳]Q�z,:�	�F=b�Vӑ���Q�����d[�Et�#0�m��&m��S'�n��9�q0��"�Bo��013����A���|���5
;;G�ќ�v�V�BM�Is/7鉞
Pt}"�go�|��1)�9�e��5@&���W�rdP���#!�2�:����5w���C�if,$;L:t��&��qH��z�t5���:t�xb�$A���u׷!�U�~1(_��� �2�K��4�!�h��X�ʊ��L�װj����I�Ge����0�$C�Sh�4��|d�8U���(�
�����wβ��y7W�վ���f�Y��I�����oL+
���ƻs��w���?���r��/��L胠u��IiKve����*��R����R1��2���޾�6�;
Y-H"�a�ɢ�(˸��[/í�b�s�X�R���Id箫��M��4q4r�%��Q nF��Y�8�YWc|�6�
�%C�-)�'��(�9L���s�a��������)-x�0�3?,�����V\W�Cm�p�E
@��?ƭ���^�?�R�E���B��\��r+�����ݫ��׎��X+�]��m�KF%@Z��E4г�
w(���֊��*p�pb��Ee�(>Q��f_��9�0����~��/�������s�.�>�J����\v� m*�RO�V 汭�aaȺ_0E�?/Jl�5o���~����Ռ<�-�޾um��৙�}��b��K��s
�6�~k{��B�X,��t(��`:��n���90�vڒϧќ���d����NFt̏�Z5V`������p�*���`�0V�]�`hXǏ$�̑助d�i:7��w	��N�؎b�����6v� �~���/h����@�)�"i\2T��I��hϴ'"�����#.ܚꥶ������kN��d*k'f8q���N�gv�޵�r i � DL����,XD/�"�'v����y��I+�F�IG�r���V���3�B�$�J1x90gYE0��N�3��������}�H0U�`��3�CH���*/u�"�e����ßj�K��C4�b��H�pe�(�C$^T�P��<��~׭��[w�΃T��[�#���e��Oӡ��5
W���3��@�\]l'�\P�56�B�q3�>�#��ضG=f�[@�e@H�Q!鲮(�� �
�����l/W�7�،�l�}r�����L��vJ3B���5@��t����L hYL�z���HK<Y�yN=&����2��T1W�d��[#yBs�Z-u})07��(+�3�~׾FІd��qoy�����C�Q<��Лg�:o����EiV���}�$
��23;����C�#�4��9;�K��F;B��Җpzw�ԏ�`�Q��ʋ�m��=%xñP©( ��-��񷭃X����<G��'���رd��r����_Z���jNw/#����k�7Y��;�d��M�;��ci�V����\�; ����QF��r �7R&nc�*^�j��)N����I�7�Z��d���oC�i^5�Ҭb�7t���-��%48k@��M���?�v;�j���W�IXŷ*�P(�>�.�m��A���>����/R���Ce�q�X�+;:mӂ�eg��(�̉�w�F�;��OL��ν���)�L������<jJ�|Ou���E���J;'�Ĥ�RÕM ���9�.��VRj��B��Ó8 �s|��^E��N@_m��[�y!$�;M����F��`��2���d�(�[��9�0������X�*�%�����x$�B@lc9���W��o g�ѧ�r�c-se�&'���n`�B�ɔ"�a_	��7l��5�*�BL �~��d^c�����(C�-^A��k�"���<dv���O�����ⱃ�̎{C@c��E���ޣ��_50l"X�������B�2�+ރ(���-�#����!�b%H���/���6�8�\���i��U;���I�|�ĭ5�h<�TB��'u���M�(�n��B�Tx	����{�v�P��@�4�9�����䩌�c̒�؝��Tt��d9E�D=hC��7�}Q��]�c�|�7��� �T�Q*_�^_���7gF�'�:�:�ƈc?Jn�F̟�b�f%��	��#����~���>I�Q6Gh?�JS6_��N<b��_^���	��u(Q%#��]>l3�=p^|y��"��߬\�r���A�5	.'�Ӱ��'>���!�6����R���<$�Y]h UxTM�*�!��� ��Q-��2T�\����hC}���y�a*ɓ�R�	��!�X�XS�\�ʥкE��Җ�����1�Phik�Y��(�sb�Wi�G��:����DV?z�@2۪M��z�S8e¥�M�)s�.�����oAp��x���L�&�S�Ǣ%ΒtN�@��b�ם����{�^"w����5��� ��߫��������t���H��T���G�=��N:y򲨷���&��O���iB�����_�IE�e���]�����#}l�%�9���ź"�Y�Q��T��*i�5'��ڝ�5T�l�IYd^^����b�י<�Ec��ӥ�m�q��.��f�#*S�8�m����������Y�Ň�դ��5�h�U~����JK��08TLݷb�H}�łRζړl�D�	füh]����=�\�ec	�FJ���v�ͨU�#�O�I�R�׹}ؔؠ�9�O��uéP�F0��r,�.6JY�������S}C}1�b#���1�s�X�~n0�k�ˉ��5)��
��Jv�E���(ž�{T{\�L/ v�0�����y�:v��b̜��bG�WA�>�<��0�s!A6g	�'���_n��4�\2�ܦ��������0�dʟ���1 �̮��6����^d7IR�4��sǠ$�����"�4a��(��+I��"�l�R������w7��
��i���q;z�pIÅ�J�����׾V^���X��X�Vx$7Bo�?���7d��CG:�	 s�({�J��P_��j8��ni����H�𸯛���o}fY<��8Q���M�frN��f�
�]~�].�H0F���eȏ
 ��3���5�ӿ�ToS(�E���n�L�e2yG�����-~���\@C,�R�{�7i�aV�]���	S�[������sdFX8��xN~����1�X)�L�cN씵�!�G�pQ�m���Re�͠4�(������J�;&�7��3Yv˨����w^�2��=���a�h'��s������֭���$ǒō�� � St)���E�,�BsK;k�r�q�P�0��5X�$쥁'��@��<��o��bwNƊה�Sc�,Ϣ��MO3W�̲LW��TV�i�\.�4�3}u*�q��k8`���}��޴�2G�j0_����k �])��Pױ���;U�:���#��c{�@q��E�>�U� lfhY�N�^�!C�3Fa�0(�`�
E����;;"�״<=��tj���:�ٵ��=�&~$�?���Ǒ���Т̈́B�kG�;�6 i��ڮ��SUQ�
� �3R|�����E�饌��)��!��	'a���)�]�.���"3�?��²K.����3�h�փ����͵��3߮Y�?�xDD���,e�a�4p���B9��Hl^`��4��#�֠�K4�d|�`��脰H�Q�m��Of���q��"�+�>���#�z-n]'�s=��C�����8��sR6c��m7Ȭ�yY���}s��Iś�������΁��&DOp-�܅��*�)#��ᇐ��&߮ul�5a�	��FP��"\w���;��e/�2b�ۋ�-����}��Xױ�E���� ��.ʓ��:}}:tH���!� ���d�����Nj���wW�L���L�v�
�3�@�?��� ^����c.K�K���	dԒ��ż6����c5fa�ʸ'�\��Pb��w�����c�'��)�� �#�	xG�@f���>°?��]/l���� �
�J�Hʐ$��|�h�]P��]�b�yUPJnn�9�+�����X���{��*x�vA7�w�9vB��5��Cp$���0�cB�9�!u�F��y�z���-X&����� m��19o��6{-E0��c�z(7���pRK;�s&��Yu��GT�3�Z��F��B��w�}�ٍ�-ryv�2�����LX_�@��y������985ق�~g�{�9�T���{kP%���G���kR\��߂��5�%���;���t�k����E�� ��G�-�]�˄�1#&!���;��i���=D�F�c��&�� 6� ܸ͘�gڟn�b&i@��a��O��ߜmYEr'+M�KLB]49/�\WL��	��V}PJ�~ч�s'k����b��!%��+��P��"�X�m)5?�t�[�?N|XD���!;�b�<���ْ��2�b� =�hH���C�:`[g�mng�0ݢ>6��uJ��/O8ur�����8�25��23	��R��PDX��;RV`�w�����Z��b�.�������	n���D�ϱ�ȹu��ky#�Qe�? ,�,����u܄0�Bf[���KvŇ�0z�W;�|@���a�	��d�����P8��vTQ�~HU�6.oS�gj�Nyj�6���D��=�5��l��
j�G>�s��J%�)�b&t���*�v��<jVZ��Y���>UC^wO��o��O���k��+]ޗ6��Yr�.�A��{k�������� �;Lǜ����SS��0K���K�#���4��!�#���Z�M~�دQ��N��܄���dB�<U�?�Y�xeL��$P���%�)a
��:�����O���|�)�O�WZ��b˙�T1Es�r/y"��\���������ޙs��rx3M�m6��7�pV�=�A66/�G����H�2��""ڍ\A��֎O�/^�P���
!�5��ח��W.P$�⸀ݣv.[]0���f�;�	� ���� ��$��ΰ5��""���˨��yDȼ��m��8����fe�R:}��&��h�c���绋?Td"�Ж�4�v�~�Eu*1��ܣګ��Ӱ{dĵ����u���C�}=��x/lb����
���@V��.�2�� >�����t��b�q5�?�i�G3γ���Vs~̞���_�
\��쎁��w�0���]��p2�%��r�kzWT.���&��zs�gCL�ᖡ���!e��4n�gIs�G���[Y��'�w��[�Q����ݱ!�SA��,*[�r��t�4CL}[��S4*����;��{��"bY*1�I��i�/���:�Pq(�r�B�w�B�.��q����2{�f��3<��F�
d��~�f�/����V$W�0Av��'Db�I3>�*�6��&� ������}��SB��7`��+<�ܿ�W\��f��~�^�.�vU��(g�� ƿ�j��*����u`��ߋ��z���s���B�D
�@|��P\�)Lן^��:��!
���0���8}}���
`�~��\+o�$�V�PwqKz���� �,kk�B�7ޥ�����1ei�:<��/6C�"��(}�F�Ҟka�rֹޚXgmIj��p*	�tu�x�1	B�UG={���`�\K��f��3��9fq��Օ����^Xz>��:Z��?fu�A�ϗĻA���)��԰��!�*�G` �PiȜ�9����8�Br4-&�p�`Jra:�_�a^�Ǟ&���3Bͪ�3&��n���	��7�:�~U�Ҹw��6�������	�f�E��xS.�yi���^�	����Dx��O���4��n����r1z������e/Xs�3�t�\��8�,�fZ�v=�F�x�HQ�E%�;\s���Ӵ詉	�����0MD.PWDKM�
�:����0bK��g���;�ʵ��s��8zn5 Wudu�������FO�1ԍ,����+w�y ꨥsW�l)k�)4�q
�OH�=]��-?N�%G����p�(�DŻV�x�E��H�_�ٰ�}&s_4QHc�ݟ�Y��k\d� ��~�ܓ�o؝�Z��r_��&|+8%�*>̶,5)�k�����ӃƷ�f��k2m���~�[�yw��lmo�Lp�hUJ�t{?СG��g�Sng"�b������ʗ�.c@���m-�UyV����(C�6Ef;��7�Z]:5⵫ѥ�TH@�bg08�rQ�+Rq���Y�%�Zs�N/�xq��T��Z�ޔ�9�(̗���#sV���So.z��´���ݺY��A�"}kI��h��g$�����<�(�F�/��W�Q�������݅
��xE�p�|���d��N��L��;��g.D����d��GFxr�CLz���>�%������?�x�+�_�qP-���m�/�o���C<������:��(���\�rس�:�.S���I�P{��(y�t�Qޙ�t_�j*���/�r�:t�$!�7��	�n?�<����S�g�3�
��kE�_�dUK����d�c�Ĺ��}?*Q����d&� �6W�����n��qk��(,8���sC%�0����� t����&��7��L�8yE�J�Pe�uKs��w��+��_�8<��NiB��ū��[�mi�oNaǧp3���zo�W��W^p�J��14�1�e�T�}���d_X=��|-J�k�5ݡ����ӯ���i~�В���U���3��V�<sV�S %���b�]���D���#�� u� �E�V�%vi	�]Ɏ�#Q���!O;�ŧ1{���k9���J����`�u���tb9o��/zN�n&�6_vgYI�0���i��ܪ?5��ܝ��;�HmR�Ռx��0a�F����Ճ|h�׃yC�������]d�7l^�b��hR �&t��z��Ք��H��K�, 17�\�ƺὭ�Lm��+=�����yX*��
��("I��>3T:<��\�O���M��^���Q���5��lm�;X��Q��n3)6'�H��cVLkzx�u^I0C�X��+���A�l�t�)RO�䗑���Y�O�4ߘ.�@�>8��GTL��<�K�yK���9�oH�O?)��Nk�dM��S�>�u˷���Tt�i�6"���nҠ���x�콘��bcy���7��Ĥ����g��׽!U���� e�p�Uy� q��<�ap[%B� ��6��a*��H�2z0�O��/�St�����OiEEY+%�����jf�M7��v���������~ط�N���7@LDm@����	`D��_D�nӉX�,Mf'�#�q[�u0DR���]�P��<���:f�v���+���3C].W�̨�8b����M�׸3�)�q0Er����Z��٫��0ԓ��� V *11|�zD�wmPn˸�D��ƗpU�3��f �Gn�� �?�',^��pX�t��p�U�&,, ���%��м�� ���3�Q�/S7Lwݣ�h���@Rk|W�k�.~����֘��޺��دB'��(:(�؎� {�@���s� n���Q�;�ں҃ ��N�40a<#�W8��OeF�fQ�q�{�dsr<r�BȢ��r��eB��Dw�؎y��?����u�����248`��R;[�m	��d&�1a��A����b g��c	S��jr�'�8:�HK�֐_�m�/Y�a%���"I]?fhS)��`���S�9���=eN�[��yΆj%�%5N���R���c��S�� *�`��1_����V�3�=JVI	#���8h �BO�;0{r.u�3���=,��o ��!tD��x��P���,���q2ٷV�s2�������Űɭ�mX�y��&��Kk (xP��?ж3�+�q�)�G,�J�"? ΄$�]�9�l4�-Ԇ/�� �y�m0����p�/���9�W�j:^,�@��c�P���m�_��Ҹ�]U�L!q2]"�O�ڪ����y�Q���7i�n=�%�śz_����Z�W�P�����sЯ�b���S'���2�Sy㲧N�@� Σ�$��=ݨ_��[L�	�L(�-عkmJ�C��.E�C����p���AC0�V��l�)��G�ED�B>�^o��w^{�*���#�g)�Դ/kP�'��N��#7����$�b��O�2��w�*G�*�ptk���<����z[�WF
����<h�c<��ׅH/@��i:�~~\��M�ga�8`��_o��{=W[�Q�z��a��ޅX�R��J�Ʌ]BU��a��l#>U�D0I�[��K	���3{����(D�D�4���-q��%eu<a뀈!��;~�:�����8\�J<WtS`;;���Z�2$���U��}/�;��MVr"����8�\���S��vt��J�0m��T~�/�_�I5�w�Ҥ�en5��ob��qK\ப��V�*B���ܽT���D����� �찉og�G�A�!�%��v�ao�f1��xn%E���}`*�}4075R�҂&�����dܣ��ʻ�HW���fJq������ڑpMjOЮ��Ot��Tyܽ��Ht:gE><l�����= �9`	[X\)��\�UˡP3B�2���tD4k�|4w�W�ۡ=���M���tσ _^}ög�f�S�_㉬<�A�r�X�Liw�*�3V��X�H~W$L�Ս&GT�Nr�yD�X�P��P�(����^�E��ļ�dnK�{ێ1$-����W�D���;�d))�x�.< ߦ.)�a��FP��c��|�?ֵ������Y�!�!R,���"�|J <h4��Ü����)A�0C�╜V.���VQO�e1��I�5H5RU:Ə䷊2��Y"�g57�|�����|�-�U���)��%$��F}oX݀�1���WaO��T�R���*��wW�}wt�8�Ö��k���5���~s#���^r�$\�U���->��aK���=_n'���/��kd�4f\�!H�q�p�̥J�\[� lr�@���/���0U�����cMa[Ĳ�.�	v�4n��C��H����W%�I_hÊ����[
�+��$�v�i�!U3��fb�Ln��] �qZ@=m(ܹ�/Ĳ �t#s9�|O�5�+@�M>`l-s�ktB(p�.1T��:�&ٟК��)1�f٢�ט���O���ظ�y �D�)C`�_R�Đ�0��e/�k��|�~Ɣ2"D�s��Mi<`����A��g��������է�t�c�7Z$e���{��Z�B﹛����[f�T�xƉs}�Œ�(�s�/�c���J��p��@�q������a�s��\�u����� �W�sQA�-��c��^�����j�I�����Y2C�q�E)���~��u�L~f,X0��	8�wݴ�FD;�8��d)�L���O~Y��B�����O��|��xt�x�G�j{�H9���G4�aMrI�Nv�kTޅ�kEk��9��@DNY>���˧ j� �:'��jf��J.U^����<��z�f9S�F�N���}�|e3/ڽK��P��7"Z6�sL)��n�����N�R��:����K��'��r޶E����饏�f_3�~E�[��nt�q?n�q�-��P�P�z{��k��GO9:�7H=��!�1���uyp���5}�F���+�VNx{��v
�Y���`ޠ?�#�$@�К�'��&���K�4+�!�P`/�.��YnG{X�e��e���Ymv�G��v�q���.Y�|�Sg|���$_�����VU� jքN5��o���;o���jv7�����Y�Dg��kQ�Y���r+6�ۡ09zJe����5�iڜ�6ɯӔh8��椣���S\Fr#����O���" �좮�r%��Qd�I��c��\=�ϖ,�o��C��R�w4�G֒"[��p�3Q� voF��̔��2���{��oӉwa��S���D��`�Vx�ب�x��."b����µ茋o\�w���pw��7��*�������4Z>	��۞]�D?��"�z���U����"���/����Jcl	��	�S���s��#}2D
"�o_d��)�P!�?-��I7X
U�O(�p�?>r>k��Z�iC����!��� JCͤZhY�����T����1�>�����D�55����N�q�gW�"��i�r�� ?8��ۀ����Q�xM����|?��SF��Ε[�v
e��-9Vᇤt�ژ�8r5`v��~wp���%���Ig�w]}��P&�M����b��#�`k�!��aF����_Q���-%�U#@��9<�~1�>�cN�����alC�*��0��/����F}(K(�)�e���Y�XP�Vt��
�q:m�58�M8��"l�x��R����.�j �y�&_6��&���ȱ�!����7���tӈ��;�����W��tr�i�G(y�Z��d�+q֔��oO�rZ�����51�^��������ZS�����qJ�̇�C�W�[��w ��y�	�J���c��t�/TB�|H��nM]y�N��$�p�?���P�ws�����l~�ص�ؠ�6GGk-\$��n��hGn�'����;z��R���.D���-�!�B-\�H�h=q�}/�қHZ�,3G}Y�uh��;�.>{��0D��������~�$4y�S6+���_;[T!���v��`�A����c:�i�aj�{��5(q�i��*`Y�L�U.��@��l�����H�Ƿ�q��:�罼<C�$-��V��]�>�Q�j�»� L>���m^�3�����T.tK��U;��@���{�Y}��g��}���o*���]7��t�٫!w;'�(~H�@�e&�;�ƫjA*�>{��$�%f�p�1K:O��Q�Y�&���̋��-H�5g���<V�� $%�8xuǾ	%�`�e�t��gI9��A8>�^3�^r��x,��*<Y�����hᛐGNC�m��pkv���Kz�U��I�a=o��W��9�s�2
y���Ոt���z�h&��3����jg	,#s��d$SBML�:�PHOH���mfS�x�t%{	=�QP��$aF���]O�e�v3/�K(����e2﷞/���v��B�(��j>�˴u\��XO��6A�("ᏚJ�Rp$��ީ�1�d=lp"�S}� 
�&���,��֙�>]T�cW��.���m���Pt�pJ��%��f;ȼ�yG��d�ّ�\a �D�f'CTq�ӳQ�o"�yiWE�O��'^�h����#����mjV�ca�[��:���
��R��2kc'�KZF� ��
�@|3W&^�H �meW_��9O���H�0���T���n�1Ш�(�heۏ�S�4�/�-@b�u	KY/I%[�����3�CB���+Se��.�˽C}�#J�s5Ųް�����b�X�5Kn�(��B��>k�.��ꕢEj�#��rA�ur�dtT�����](�Ҋ�h��k+���*N�e��#uxbo܈�xku��AU���F�qO @,~�2z����02 O�r�H��!o8c~6Jb�vAe��x��AEu�m��eR������&��e�c��#ݒ7���֐�Vj���}1�"��K���V��[���0,������	�]߷D���fg������3��~s�}w0=��B��T*S3}#C���ƫAB�;�P0l��o��{A-o�������_��C��G�X�ɇ�Ϋ�4Z��$�YF��.�vj�k,*:`w8\��R>Ru�W�Y��g�g�C���`E*C�#��=�7�k-��q>f���m���.�����jv���Z�[f�̞*vρ�x���[��u.�W���UG��YE�샏����8F�ӈ$��}���[�ҘK���!��z��*	_���k�K�VgM��*���B��(30��9�V������!��3�Q�mo��s�9	v�^�gj��D;ه_���0ctT�v;��?n���1s�A�0��l��pm�t���
.�od��ww:�[eg_�9��j+��I΢�;"߼��U�r�m�����K����L�~���RL\��WT�|�d<�".���_� �nr������:�y��e��R����t�:2���Cu��\�^�g+&*�����Լ����]�6)����u�a��zX�"�u�z��-�I��:����$�avF�P�nH��&Ӵ���V!n!'����3iW�~������[�A��R�41JuX��Z�����\O�seY�#r�o&��-����JC��S\��[X���������9�|��~יy8���fF������2�_��_��^
J_R�|�3�!+�ɢ��
 �������'��!�N!�!��H܆��������qt��A������S��߾�k���
li����8�r�+tZ�="r��3O������*�Z�eVþ��7\��_>I��5�3��z���jL��u.�EK�W�?�?Z Nv�K�0�H��y7'�~���:P�i;��}�C��n,r�f�Iq���/N�7��Z`�e��$���������Q��i����/V�3��i��G�}��ZYv0��zԣ�nQ����]$4|���i4�?�@/7��h,�2��
��i���'s���5��e���ag�D���X���zQ��>˜>����R�L��=��|(o�1���&Ɯ���)n��FS��g��`�W���w�7-/�E�]oߟ�pآr�����H��I�ԏ���#�2ᾋ;S3��HƱ�(��@���M�"D��S�)�l�F�g�z��a�L�I�Spч�������r�]���U�U�����}"���)K�V������1~�\�Я�ڽθV�����v��d2m�҅��d%�X90�Z��P
X|�˄uo@����5��:E�O� �n_#�AP�m����y��}t��v�q��Ҏ�]��|~�����ҳ�����]f�L���j�R���+w��d��z�?���=��*�pM�eLo���&N>�!Us9�o�Lb�������S��Q-U��#�3�r,_�kB�:bV�1�uG����&k��d�%��pq�ب/�

3-y5{l6�7�4�	�����	q��$�Rp�9-�;�F�ۏ[��#VŘ�4�w����x)��vvx�Yfa���g����*lT�6'���P���}O&Rk8
�1�����+ly���t�c����#4sj��ߊZ���'����o`DϜ�?�*[\��D�?��J�Јx�#�����y{{�Gڞ�.)k����Gdܢ�W���^t���i����0�}f~xr��Hꢬ�3�#
�r�u%�x�]�Z�c��P���~��8�O�M�G�b��77��,��T�	[|�S���q����?B`ɺ�P6�m����yM�x�m��I�(����(�aY�v�^��TB�vd$�(E���8�����C{�Ͱ�aX���ҩ�,��R�N/r�#
j:+_9�R ��Y����3<#h �vڟ%�9 �Z����Ayffw��:(\�����j�k�:&8��[�1��3|4��K��L۱��Tݰg��Î�O��Od�	ゴ��}3��9̛�n�/�1�ITz���O�=��C@�KxE!9���D
�������F�`|"j�W���Ep��dZ����<1���'τ��,���y�\B��]��]�L��gy��i`���*
-_F)��`\o��}�T{��	�B9z���g�-�y��O�DG�T }Q����|��[υ4��#w��yv�h|d��k�Y�c2$���{��	�>��w�{��-�{��)���y�p���|�a��c����D�H'���!�v��Y���I.NаT9�U��Q�u��Y(�Ł�fB{��3��x�8�P�~m�Yg?d�{�<8x�$�N ��<IL㚒'��[��2y�~��{D���+�{�ɞ�� Q���gĉwBZB�@�e�@&F��v�������`�VĨk-�;{Ҽ���CGK=0�-y�H��óq�Ϛ)5�C����H�1e�ހ�N�?�F!_�mw�;Yk�P��-�w��G�Y�޲X�=,������Y]�e�7�b6$�@ܽ���3�T�d%�jg�BW�4�7������Z�sl������8���'HQ�o��8��P˽9�%5�0!��%�����g��������+�{���ӛ��7�<�u�x��l�v��"^��QW����ܷen��HO�b�-��R݅�2(��<!Y@cV��҇����ș'o���004u�2^��xFt-I������e����*��5�b��>�-=ѓ����Ε�@��6�r�q=��D�R�����E���塃e��2�h�ޤ�Ai���i�B���a�Px���Z�lr��c�M�h�\�d)�)R ���H���5�L�%�>�H���_G�����z�l#�<��|��3�=)��F�^�;R��g�4x{�1i`z��c&�NZH��d �WK���,4$�~?W6L���>N�'km{$���m����xb��Z��yw㙬�A��-A-#�iflV�4��"^�=�~�V,Q!�:H�C��XGE��sg6�2�t��晠 ��l�V�ѡ{��helN��V�RpI�SN�Z�k��8�<^-��Wz���Y��O`�yP�`ʪ��2T�_��]�wEMڪe!���W)<9lӼ���GPF�``�]�'^g1��t���U�c%���$�3���i���4��%{�%�=�?�����nf�"�QN#͚�*���n�(�a-U׸�HC_>i=�� 2�5YX$�h?L��)�N�i���r0q��}��_������[�0H���h~I\�J�(���V�#��7t��A�!�a��ÚS\.Ch)�����}:��N�u4��,�ƈ��ʸI���wb��T� ��5���(����#��f��ū� \<s�~����s�Y�R�.���q ^e���!N�&[���¬�T&�P�OОU����j�Ӽ�J��y�!;����Δ~��7׶!p� �6�V�vE|t��=>� y�1�"����%`�f:�L	�u܆���iP!!�AOS	����)��g���ܺC�����u�x�M��R�T�mC�6���d�^}%�c\8��/��5z�-!&��(��/);z�g �X�wī�kb�]���x���K�� �\�0�:z��Aę�k��Յ�C[$wĹw�g��WH���V�[X��ˋA�7����eLP�b?�ÐKs��U;l_��K�}-U+նem_��oR@Vj'�(��>����@0��&��<�B6;C����shN�_F��!���AL��){���Mx#�ə��7 ]`V$�ޗOݵ����3��LK�3�~Ĉ{51�%]&|f&���c�R*��Y��v�ĳ����u���8Be�pu���L��`����&�L�k�~�!�6z�Z� Չ���.��Q���viX����=:�l�o�����@)��Wv��<:5�h��g]5m"����0h3�ʢǈPv�He].E`$p�Y*�V���;N���ѯx-���F�^�ă��*��kDD��aE�"�.`#���s���d(�R�� .�xó���?R>�]�{���%wE4�{{��5 K�x[1��O7��Z5���80�
��F�15��o[d$3�����g��K8_}�a��Z�����Yo�2刺*x+����O��*��R�A��"X�D�́�a�ED�2R�H�h��B��ɰ:	m>O�4^Z��K��\m�OQ��nnp�(�X[Z����H�a���q�}�"Q����7+��lݷ?r�0K����t��Ō-�� ��n0����t'8M�� nÇ=]K�;���A�BM~z��RwZ7�:��	�7�;�}�r��@����X�H�>H�mD��3�߶=U��B¼<��U�W =����<�)� 9�͒���{M��P߰Lij�FXQ��l;!�Vm�H%�L�Nn_�n�t�����)ȼ�f��OkT��ˑ%��Ot��'�Ĳ�)�����h�#ʩ��H�<���/?~�߶�&z&����PW��Н��Ju����Ab�/�-mp���v��%v�T�_L2� ��8�8���5�P�`�ٸ!���gu��?��S�i�=��Pw��G�M�?==�"��J�w�T͘l|�S_��HǊ��YR����ױK�1��v~��k�%mɺ��	��G�\H�n!��3_��=0�n�C�u�\�RFeR1HK��F��;&�.^�	l�H_\r��X�ܞ�1mz>V=����±��ŏ���'oQ�#XEѵ=o�(��DB��������O�m@qC��b��m{���'�:�:�#��]+B0N�E̷l�*j4������'Ҙ � K����Ɍ��%��_đ�U�v�|�� �>��;@�N.��yDG���}��K��͔7H2��{��6�ײTr��y��XV<��л��P����Ƃ�s~67e)���N8Y�:�ؘ��x�D�K��
����6�[>�Y�?FJ�E�EK��#����w�����* ���8�[E��*�[�>�l3Bf! ���yjQ}���Y
˃�N/s����I�`�������z�3i���;Qk�y\�����ߏ,ڳ��^h^i���*��a�@h��������R|�!@��k�����_��-���T���U����<��?�7zc	UL�{uu�v�V�z���W��%����M")��P���'�,=Yyk��:G^c��Bˬ�X�!�ߢ�BzV��n�0����W1��|;tX���׹��}׷���7�1��,���|
Nǣ�_+�ǹU�6$2�P+��G��C?�)1"�w7�'���)BI!��s��z�j@y�H����*Pz�VO3Zm�O`f��� ���-�z�E�3P3C)��@v+S��	l��<23E4�k���{�������~�xU��<�P�U\���+<%�c=��e�S�#�R��U���������W�I�?�� �qq�sʹv��0��yr��NV[����D3�o]H�:e��&"e�����m�ߎEUFшy������W�]&*����6�my�IlV@�C+�fS⡸�f�ņ��rK+]�\�ʭM��b�����}��Nr�=�[�_m��`@�40�y�#�psti?1�����6�*��ښ9Uv±K�O�*Ipt6K��{j�UG���8���p�3¤�ZM�{�84���j��,������'�BR_ø�J \2*|ʨIJ��
P!��|�<H)�!���mz�4���{TQ���1��Gl˝v��N�Dbn�ޓy��<�6".�t�Q��os1{��p�ň�BN��@$�!˺�����QjԘ�N����#��7D�n��h�KO�;�G���}��Juג��@0r�{�*���8��g�?zyB?���!�W��+��a.��@���)P��-�h����M]�CS��l��Y��jc����P�g�7ג>���w�r?'h-T�B�X=�i��T��7;����ae����� 8d�������S���dq|��=�r)��k��t�
��A��u��s���.�`"s��.<�lA����e���nę�P�����7ozh���u�?���"�2�ĥR͔97�Tn:=�=Բصף��-K��ē�A.[��Q���F���E��:�!z 1�!Z��G�*���c�������"�hB���C��� Ú��QSW(M����Y7�zx���U��N��6�!�נTJ�bLa5 @'A>�F����ٜm��=%@�b��:"{�7.��L�_�R�"ۓ������ku�X��[t�Zr){��W%X9Z�{�!h���Z�F�v!e1������c7����8�o@�+A�(K��I���s�c����;;�r����X���	�y�$���bɄtr�h���6X"�Z�w���!�\�⣦/$|L�n�:�#Z��TV4L��Z�'�����D6�V: ��rd]9���΢�:�Zzj����8b���Z�	��Ş)#LB_���Vae�82AՅ����e^Y�{���{**}n�Xt�ؾ��n�Y���|�p��i��Bڒ`i4?8`=�O���{ll�"�lb��(���)�~Lנ�.������6�zs����&��j��߲]���$��Q
�!��}I�j׋Z�7����+&Ҵ�ݒ�� �	�P�U{����c����Ur9�R�ٝ�����g��^f��Xh`(
P<K��}Wn� X%��;ܣ��p�.����B���rړPּ	g������s�^-"4؇�;@cz	c�)i#¡��v~����v	���tY�Dk��r\akQdT���� L�iK��m���K)����YA���_H]�(q��˖̘�⇪q=س�`��&�Z4�������SpȽ��r�۸~9\��V�/��r���ڊOy�/�52!�B[���3릛�@Aq�Id'cY�D':����:����F����c�-K�k�a>$'E�S�$<����C}�>����|���*�=����ޝ����М^a�ށ
;"�
�-��l�{V�TT�7� ǚ����s��0����6f�SJ�\��,�������2�*1�6`����yx������,N�`��$�d����۔AC={�܊�OL?[�������WZ^��;�Bdw	��׭`���pj�%rk��t^�p���q2àUt A�Y|����l�\|�!��7��4λ�ͭ�ۺ���i3�͖������G�7�%��|+(g.���]Цj_ٴ�����L	W�,UV�HV�"ɵ֨"����w�W�p�xAFcr�T�ڋ����e�]� Dr%�F�]vP*�	fg�s����1k��>^���ԧɲV��괱��I��H�8�^���!cN�6�?��^�j��	CED�z2��fE�|Ή-C\��ΎuQ%��;�v��u��ćL^����s������l�A��|��6*C�pե�웤0K�*��rv���z���$��('R<2~<2u��������t�c]�$��m}-�А�'�'LD8S���S�x�������zIÅ42�XT�I��s��UIz�i@��]qOy�t�X��U��}�~K���:1�zZ��0(�h#x|dj4ø0Y|۫��Vh��3�{)�IBQ�^��ܤ���
E��X���?j�䄫ˈ��/��}�G�mLBn���A���sd�b����Ki��zeA /WE�p]�O2��N:���p�J��agL��uym=S�}�뱀=-�-�e�{S�[�!Yv���m:P��L�P�$�8"G#�o/��/�`���4�k/���9����{Gs͜��O=�Fr�F����	�?����f�<t;���7���G��N����u�IpA�¼�Ӌ�`�&�]!؀�%�M�l��|9�;�:k� �$t2}i����~��L�Όg�(�����p*��)/
�г��	C�����|.��j���j &T���<�rK� &(���J5�?Lїnmӻ(��ڲ�sÌ7&�u�S��Gm}�J��g�`���F��܁� 7��6|�³����i�)	�@��ԋ�m��w������~�2.w��<��)��"�,�d��9lD�r�]�ua�Wc�Di<�5-����2��K�+�˯̪�h)j��=$F�~DĖ�5�_{��nFc��=h|	^n����օ�k]�(qN���~��R�x�{ˢ���!�z���\�	2sI}�gvlJ��AK�Mu�v�$��цϏ>���{9:�3eB�[��z���`�?��ϭIC�%���!բG�f���Z�A�L.��u{��{T�׺����Ay�d:;t�d�<�	���RF|d�MP��9E���@1ĳ_I��7w��%%�@���KӷA�A5�e���xLc���<�!�L���
j�R���z��� E�'���y��*����]%sr�F��D�ʋ$H�g-���av;`��v�}�%�%*O�Ȯ�*���E��\'4Jd�^R�����n��'�Q}�[G��&�!>pN]
��/Sܩ�������C�߄h�*ܵ���=.�~4v�ۯQ=��#ʚݙN��W��RnYƩ��p��Oc��x�V�0��8ٺ��,���� �a|�x^�S�HJ���� ��۹�tcy)�P�ա٢ .>�)��-%�41	�P�t��pO�i���V��6��Iq�Wc�*�Ȕڐ���UJaN�9	�,������?F�9�	KKXq3B{~��a����'JB�lS�X��%�M�W���6�H��h�A
�9��ȝoT;5�@�����VT����Q�b"���ʄ��x�E+҄�!˱��ޞ��$+S��[��^�?����l�;�6�U�9dD���s:�w�{�A�X��R���tVf�ʫK�h:tp&?���o��ࢬ(6H�����d�ܻb.��-�t�E�i�JV�����n���k���K�KφSܦ��_*� ��ZG{'����F�㽯o��z	qB�"�m�zu�~6���7ь m�~VŞ��I�mE�=��˚Miz���?����n���5��;DJ]U���2�����J�O8l�JA��Ag��&�"���`LX�/���+�\����A�݆䠥٠
E��@g�bqU�Z����q�h��vҀ�|���v}��O#�h�����C0�� ����Վ�Y_oaڛBzb��m�� �FΫ2�ݚҙ��_@���^#�Pk���B�㖧���n[?�D"��o��
����6��ߧ
Ǯ�)ӛ�i�j���B!��)Ch�֒]Ȭ]�	�z�5
яܯw{��ǙR�4����TT��؟e'=̾�D�����>%�N$��Y��	/�K�pwߎ&��i��d�R���Y�N']�U xk��2��ԝ݊H��&=j.g	k/�㴶U�T ��F�f}��x0 �թ&��zk�A�L���:�W�"G5�%-�m�my�IO�d�A���������Z���
j�%��� ��rh���ӌ�TH����=�ߪ���p;�*{���m�C�ɇ���n.�~�I�("��aԾ������L:��w*~_�/�	���\� ����Q��]�).��?�=�TJ�
��r��{�����[�!��U��e3�X���E�A�!���}H�x���o|���nv��z���=��e
C�!c��\��{њυ�|q7��H�,�&�ڞF{i3}6�%��Q����iJ]'$�'ME�������	;O��_�]w&[�	DmBMEQ{�(����'7��=�}�ߖ�<�ﶂ�5���h�����(���fW�؅�n[�QWz��`��תh�͘��.��V�9Mg�wTIqLb�Qv%4����@�7�t�$���ׂ��&���@��K��ޕ�1�9gl��pѡ�LF����1����S��r: 道˨J�iS�|��T?9؎�9���j`CĲ{/��W�S#@�(�\	�<\JpA��l�\Ţ���x��x�~��{�%����R�<��z"�R'H@Z�s�m1?
�]Q�k����*�ª.t��w��®�l!��lk�`��G�U1�v��ԼU8�i�y%u��ZO�GZ�"P���@�R�J]��M�tQ��?��!j�>EE�3��m�I��@�p&I�@�\$��^�FX�zZy�)�&7�nDs���Z>Cʼ�e\�U/�[�ȥn&��
+*�X����g��֌4p�R�{S)� �i�U����U�B�N 3WKc>��uj ��T[�����Í�������b���Yf�+V���(;yEPeV�r��3ГL�I�q���6�'뒸��F����Ci�L�׽?�ƻ%��������ANv��M���O�VzQ�-8y�72�*���qP>rb�`���Z�b���aߖ��.E�à�/��8�7�yO���drV�d��l� ��L#�9v:�`HH]������c���uSf��QHLITՇT�������g?��g�R�HO�������6��~@�&dbo��PS�:��K�p@��E�}���g+�	R�y]�7)�t�!.Gg���|Զ�[� ƥ1�
]�IV����Iz}������Y���[n��@O�Ӆ�	͋�+
�!5��L���ԂX?��p=�b?nʰ��>)�~W��*}2����J�:�9q��~l �8��������mr/��ƺήWG3,5���� ��>WH�k�}_��9$��)��)�oڟ��12߉ɛ�fu�����p�ɩ<�	����"b��xā��{�C�v���<�bx�b(W`�83�?3�aj�L��QՖZ� ?Z��*��$�W!�LR43��<_s��&j���lK� ���]{��%U$�:����8���ץ"oҗȇ�Ӏ��WY��P��y�;H�_�Yqu�ӇTxD�A �k;&,m�Z�B,F{��.� ����/H� c��Y�4f`"����<k�O-,�g�F��_��YKGǯr�Z���@]8l!8�st#~-b���4V�U��/����2�`P��R�!����i�(��o��(y��VI�1�zFy�Wi^7djtR�ʀ�ՠ���ѰŅJ�����8��n�b�PZ����K��7s��@��8���#��r(6eʘ�aA~�WLϹ3�}-I���_�;�eޮ3p�/�t�[�1ȱ^����V2���k+�n4��k����D�B/��&��U�~>f�~������Y�w{�PD�0���v��¨��7�(	y�Ӧ�V�0չ_F��:���*�%w���E�'@��Ki���F�u��&��,7IҦ��x�������Af��hE�����A*frx��oj�Ol0�����xŨ��:b�K��N{���~��A�1���u/K���EW�#UJ���J��*�a3-�U��fv1ir��V=��x�{�O	UD@��Dt��P���k�	��0d�S�u�6�w����/�p�=�+����j^-�~-�yRvL�����Q���Y�Ŗ���<}Z�@ޢ�g1�\*C�ՙ�[Ɛ?��:}��
L��Ҙ�O�U��҈K��9 �?�a�̆�،��S��w��{I�3>��&o8 FkJ`�#��� � ȫ��&d{�.	�����j�\���bc��W?_o�D��W�����2P���e��C�1�;Wp0҆9%+϶�R�_O�MI��U-#ЗL���#����Q�1%:M,v���tbɰm���3J5i'w^?�dL��3h��.*��m��B�ع�yP[�9#4�f ��;����u�9���d����|.��9ĕG�����vJ�V6N�p��ԙ�|l(�BV���YК�~����N�G.���nx�����X8��KM$7�FT��)�²�,I����m�4�"��Lz�cc���0���!�|3/�Dq��F��t2ڹl�D�ގ�iI����h�=w8��ȶg_�hL�3+�+���ȋ�p��ބS�+w�+8��Ox/lft0����1߃i�(��a��Z#���v���;�\���n'��p�Ї����7u�v!�($<�:��F:�=���ۜ�L��k�d�|����xU 9֧�Au6��|����˴u�#m�g�D��7b\9��k�ib���,�>p�����t��VEp����fG�V�ij�k���������}7�}��ğ�d;͓z��pQ�%\��� �E/XT�ѡT�A�v�!:k���}����qO��G\A�����F[�K�16or�*�fw�^/�d�����[� I)1�XXk� ��[�9�0��R�{f�ew����&ˡ�OI�1�_��X�]�?��rBvq�c3��'-�*��e?w�2��?:>Q r��qDN��L�߄�颋t�4��Z�+��ρ��y����%�Z�����;VV������Հ��~L/`wmV�	$��VꀸJ%�dI+۴���1���Ur�I,	2����[�`;eׯ�i�7s�ڡ�O�i�x_ �+N�4�·�
�{�u�����'4��L�H7{xw�W�/�*I��i�j��@ 3t�䗖AؑbO?�y���q�!x������~8.!LNUq%�э�ҥ���_˹�4좧�(�����y�;s��A]xsj�'�>�EQ�|������<1��XKTA6�A-�����o������d�P����2<��C�����N�3r�(���J�§}�/!���8��S�3�Z��_�����ړ�� PԊ�s>��;�03-�H!���t������"�8�X�=K�����Tzm�����f�	���٠���m�=�+Gя���`Cq�';ک���*&Yέ��= ��b���J#�j.
`0]~ly7�#�2>�7�
['~"c�8�y{ N7G�������/�O�\)������ʇ``釩pPb֩�br��4����@X@��*ltΈd[D`*�o��+��59�
������ӐY���l���qrIMf��k2V��SQ:""Q�%�B�Yn�E�h�0pT���Ғ��w4���� ��+t)�� ������yr%ūa�D�4�cQ��!�� iT�����L�=8���V�	�
 V��Lq=�O������LQi�x�A.(Dl�7�2L�y1� lq���6[��V����ʺQ�XCY�.@R����gx����([e-�1�,�" Rp)wO�Ҙ�X�o�,ͦ���]�~W�t�eoK��v�q9���\]{�i����!�(B*fHC�FT��ȕ�u�ڂ.�7]�[p��#�$���3�WX�j~\#�ֶp�8�i�Os�����:�࣮kf^s��<���^���(TD�0�Y���`͛�Հg�\2a���b�4q�T)+���iT�N�#� ~G/�ݠ�j��2���eʈGb���{�oL���~��d��HB��G�3�M~���7hz�������\e��5y�.����S'����\����?t@`Kk��}�)�"\�$0��w{��,J��g�����4�����}t_:GS��BI�������/���T,�W��K&'�/L����2F�a3׮HPh`��t������m��7Gv�6k���G�!��5��g�0��G���*S�$D�;�8��G6��E^���Ni� Gz_|�����<WR�߬[���q��qh��R:�4sK�U�$��'�K��X�0���)n�����u�穩�s�a��b�6sU��{*f�5�3��� u��;�*>m4���w��T.�.�V�D�Ȧ���bI~�Dz^,?p1������-����I�А���;C��Zqo����.���Mg�LO���M��?B���N�n烘	����A����v}ϋ9�JM�܂�S���	�	�U�Uw��BOW�O�QC�[I� g�s�(;�����}�l'�h�嫊f���z��-�������цH��G�s#5�UXb�ؐp�ZX������ l��%�u�F�f]�9f��)�BT�|s�-���nS���jy�-'���P�;�������q��39���95Y
� jp��TjC�L�{l8uyl7K}�cW�����%ܖ$�Δ�¤ф��^暇��5 �nW�����}�WC�nO���A��Hd�p"*���F���<�FAV��6����c���H���m��%N\��%l�=��;c�J�5��B�*�S���B�k?���p�H������7r����Zq��{�\2��I#2�u��`��:�?8�0�F�w�xw���p"�]�#ߐy�kd(H]u�b�;&$�L�Q���[g��iQI�[�ݤ��'��Iͨ�A����V�b�7�45l[��D�b�</3!Bv�9�H>m�~��Q ��t���I%���M~��j;���L��߾�qh�8���"���~T?��XQ��u	�H�p��	�D;�.3̡�C��P˹KqeI��54��
��fZ�����3��c��B�+��_�-ؕj���<,�ܺ�������=�m�`uA�g�xɥz���L �X��XHV<2�p6��jm!��<�E�ͤ	n�O��ၓƧ=�D���䯶�:R&���C�L�.���L�F�����9�Cƀ;���/��
��J{r1�<���l�v�D��d�p�54���C�V�m�E]�+Z�D�%It�V�2R��m�h�"ĿlU�u���0��T�b�Y_��2:y�&��t+�L=FS�Ɨ+�W�xY,{W�q[�͏O=��I��b��R�������.�o6R�	qӗ�c�g�l�<���6�o��4B_bE8L�rU%K���[��c�tC~9ю�r�聂�}ء��qٶŤE��H������H�b��h����I+Z7<���	+Y���J��Y%@& ��~5�_�3O����z�o{ý$��F��uEA�d
Dv_v���Xye2����.��6�U2�W������{�/�V���N<�<�On�pr�9��5�<����2p�Qu���4/d��}�n��A��eY�|����,��\�͂��ܛ(��ř�y؜���m�'>������>��^�ֹ/����ȕS��*��Y�3��e���M(�����戳Ց�T*Ϋ��}�Z���]�l�ȿTb~#��:�B:��ȁy�>|D&ݡ�ؽH�^��ʕ�͉�T:�q��M�_P��o׆��ɋ�S+��rh��y�?<E�̗�����r��m���iF��S,�����0�>��ȸ�u⺙��B��� >GK�T|Q<1�F�v&��ߩ�^y�z�\��iK���h�K����a8da57�8p�A���\ �$-�aH3�Őyb�Kޘo�	���p����rh�B�m��ap�ڱХ�;��K��}O��<����i�G�r�>�ެ�:$��p*B�T���ip�!3B��C�T�A�/�Iq�u�a*by���?Y���|f��'�`�b�X�5�`K����͓�ᰫ\ ��ۜ�7O���3�/��c���s�o��䓹^շ
�ب�ݽ��_s�.�b��d�>Y%���4
u}-�Ocq��X�Vl��.�-��b��Nu�Z'�R5X}�y^�W<�k���rr`�KSwVr_#��{���Q�a�ߟApqƋ��<��k$��9�,)��R�%jxe�g��r���l���#7�T�@�M���������=�U��lX�� ��TG��M��[r�q��s(��C����K��Jo�s�3k �����h�p�������+��d�-z56������:1�V}A}��zu�/�Qv�h
�;�h��Y'��E��ڊ.xLQ����崱BR_u�]�V�F�
ȢՑu��]�([����_n�R�)�i�k���x�'��Ñ��*��%�e~
�i�{�>��R��ly�n������+�G���{�%�}I"�y@����b�k�DA��o�ȯc6���r#Q���m5C+����8�gg#&˚�w`�Q�[^��>��[��C�0�U��4-��=%�ȔV����0c���
�[y���c��+�C��A�^��0��n��Mb�o�g�F��,\��7q��CO��V��c�o[_��z� ��A4�i�Q@	�oRD�ؾg�XX���kX��;�Fo�{��6Uƣ������0���u�J��K�����T��}%�t��*	�����]UW+�5�J|�����t�`�q<���Q�$ �v ���	���W@��>�VC?��!7��^-���Ǣf��;E�W�ԡW�7�mx:"~Vr(Y5�*m[�y�ď�u�����G��2O:��� ?�V�bc*Q��]҅`;$�=GU��*e�dK!p���)�t�p��~D�O�N��-8_{h�ә��
6���{ �eb�0� 	���ގ���w���o�T���W�6������]�$V��b�W����8���|����Bjw�k'QT���X
�?{�R�:°��$���]�?�vH�.�(���Dk�m]�+o +�<Aa{�n	h]3���[����,4=^"�/S�?�<N�����(�w�j��qm�����پB�x�ip���:�YZ2�������T��'���9�9l��t9Z8��VE�Əԝ��{�WW���-��ˇ_��t�����s�5\�hW��L��f�(�}���j��"��k���]��v��Ȇr�w�#�~q��c9��v�V	}QWVݓpu�q�*� ���%z6fԢ
�t(���A��Q(�Q$�|L�wɼD����
t�_]e��v9�,Q/i�T�)=�:�;���k�l�l�LCR�%�q?�ϾX�dp��CV�C"7��;�Q�� ���{鷜:[�}%����u!�3�ڎ=���<�d�48��=�栿���|烜�����q��B�(̤2K��s��<C�����ӧ�ϒ��,r��-���(`"��xK�O�3�F�}'�}5<(\զ����R>h<BP:�ˊ�f���4�"�,��9k�2uK�R�]ė"7��?(}C�H>��w��\��Јe����;<��@��j�<�S��Į�E�>�*lv2T�d��/��(D�	�
��U#�W�X>�!��U>�!��c���ʡ"Ũ��Шl�ٜ���g����\�U�<)�Gi�6Oq�#ZHl�r��u.Wt���17�
_>l7�%�(dٕv�8��l�a;4�	�����Q��G�s�pK����:��F�ʌ}���]m;���_�v$��[ɝ��Ӣu!Z����Fj�#���.D^��)�3M�A��ef��F�1��.X��m�B�&���.��ĳ;x��v	��X�����2����R��VI�Bd��#�i�$�C�~	F�wԭ��&|sB�r�\����F͖��f'���/�U,�Cw���6��Lܐ/bg"�}�9�P���N�Ȟ<�N{Y���%���=/3F�~���/P�8iv���'� �$7_%ֺ�?�N�G<+����h���Op��Ѻ�f�`��l�7�X����[��;Я"��uOCb��J� ��%��2 u���4W:T���-��j�!��C]IrE=E�/�`~��'�|���PX,2��PJ�}�"��W�o�o�H�X�P�!�۩������$w��#8�/��G�c]����18���(� oxܺR��G������mS{s�X~��l�/�0!�t�鈢�.����(�Hbo�����`�a��Ba��ژ�m�1�.�`�Q%'�a[I�?b���gA�Cv��H��$�LC'.<Ρ���������<
^�،�;�s}�>p`XFe@���6�����!�N�|�Z���T%S��E���
p�1���������G�p���ú7�	Q ��R�>�l��O�Ѐ�mV�&ْxnm��+�6��|d�x�c���ڥ
I���
w-��]��g�#�[f�tZ�2���6����~���ڧ�A;�����N)�Q^64a���8�y8q_$�n��J�Zl7�6ĭ��>�n3
ڷ6s�b���K"ܵ"W�����mTG���U��å��Ē����l��D/��Hv�'���8c?<�!��CTm{����l#��/OF:l^����G˿��&�wp�yT�e��� ����'�m~r
��6	���h��GE��n�g4��r|�v+�� q���h�My�|��s!�y�-#�&&%�q�r�"t��ո�F;ϴ�,��V��-��sWn|%���[�(Ȑ9�n��X!�B�R׸��Lt���g}��9���9!��j�‖�X~��'��}�lp�G�R��LT����t�7�g�W�{����!w��8
�Yl���U̪L5���M���W��Lv�~"��/�[/%�p8A�;����$�Ć.u�'�a�z�&��\B6*0�R�/�#XM��}�BG��H���>�&J���V`��+�x��:� 2�~��J �h��6(��L�t9��u-��S�!�-1�,�O,�
a��KE;^e� 
��y������|~>�7)L�7������T9��r?ᦟ�f1j�
aQ<n���u� Cg�.�{�K���W�٠AA6�O����]Qso�?/��������P	�Cw�	A^;�v�[z���f�C:�z{5e������ ivɎ:���Ph^9)	��N���+K���/��d�6���F�d�$��4K��!��&q��.s���|G��e�D bm�cy^��z�ܣ�_S�qK�����̡��rj����j2���F-|�si�i{������Ͳ��N�{��2����wԶ��0$��r�#��O�$�л*uH^��%���=�5�rɘ�hf�:�m:,��N�QzH�"s��vYP��S�E= 2���a�kD/��T����_�����غ���[x�݀�VX��ِ��T�7s� �o�^޲� �1ʕ-�ܨv�bq�b[U�-r����E��ѐ���G)-�[���Ǣ���T��Z��;�;,g�kk�,������(���5�qa�&����̸2j��+���qr	��ߖұpK���xΫ��r�����Gf��*.(?o�a�s��Ӑ�����%�Z��n^v�)�f-B�\'�*����T;�U|"���e���ѱ`J״�i���3�5 ��U{�4�f��v����u�ZL��Sex|z��_�����<�)v9�3�٥�=�	C�4���C��4�%(M��-��S��w/�Ā����|x�� 7�.�F=������=�yS?+̽�OIg���9h�U��S#:"����N���~PӚ9�Uf�*;�	���u�<�v��W/��)��|�zn`C�Z�jb��ꅛ�	����]^�F�+/)�}<���Y�Y^�Q�%Yc�\M�u�	>:���%`���b���L�=+�kr�'�qk.���uj#��^������H�Х1����Ci�7�bxH�C&��º�"je֝ ����z\Ǐ!�����?8����\�{�Hˢ�,���i��A밁fX���Hj��BDӡ�&8㰨�8�������l���:Ϳ�%��W�*�BL*0�I/��'�4D�t.*���p�����=�V�^w
���\yP�:��	�����TZ/<�@�&�k6ޜ	�~�,�Qͱ0���"���F�ɽg[w�`�ok��n�S�J��,%$�,�2&�-�̓�ii���鑀&�ֵ𤞄HG���ede����Z���.�S���H;��e�)YsA)֫��lt��P*���nX��wpK���a�:����-��ȸ�ؠ����)-!���Cyo2n�@��K�����K�%a�%�<��(�y�C9�7�b�L�7��=�w2q���Q]�pA��P�=�h�����왼��W��o,8O/Ρ��\M�a�f�cj��L����RLåΏ�F�n���Kt�E�
o�mT���kn�j XW
;E@�`��^I-�v�"���Ks�1�W�D��$,�Lq]�z�3 �m������u��-8�F\F&��[���7n��ً7�^�{Q*���.��ˡE�~I�g�9]M`�d�ez嶩�k�� 8���]���=97�T}>Y2ti������&�ԅ�m�R6�\�K�	t��r��f��:+�� �Վ#�V9��:�A��A�)�ņs@{Ɇ�4jR����\�V������l�F�n�fl�b�plkw�'\�Z�KFu��a�$�Chmm��l�H�N�}��t?�At��@YN�g "L��{-̥t.�rF-�(ˣ\�7c
��iyL�p�m��g � �a��$a�5q��H�P���Y��%���݁�7���e��:��yަޖ>�c��lx�����˹��Ff���ߴ������<N[x��M�,�6s�`E#� S)�	���[@j��0�Y�cT21�KIn�hXB Й���9��خ�b�8V�EQ�.��mxm� -�I9��3YZ�c�hq�K�o�]HB�����p�w
�f���m��f.� N���.�܀����;* ���\&�]HZ���'c�5ҿ���_�a�R.�����F:Z *;[E�'�I�5�I^��?��e�\�̆e	N�������q�)�����{9r_�jva��&���ȣ��Մx$ď��öfP8Is�=}1=D�ڦ���S��#��5['JAEC�n�k>��V�*��HO7 9���B�dp"�ƒ���� �������/G�^���g��a�N'p�`Qx���kv��:�"�q��4�C%���M����iµbLS�)�{T�ݙ}L�R�� ��˷�K�Yi8��0Î�ܳ�n+A���D���<e(4�bLm%' �S�<�ՌHy�	o��t��:���o3d���M	GCm�>]K|�۟�Hꅴ}���(����qT����q7c�+���Ԓ���q��'�˳��@t��sW�����8��J���鉀�	l�j��"��汤��[#3S�1h����E׵��H>Uq��\+h��o7R`.�Վ�;��t�a�Ð����g��;��=x�g�/���۶�����E����V�wТz���q�P�tE���Ԋ�9�����U��*�/Bj�N.���\R��9fq��>����W�[��i{|΃lx�?��计�F\k�Nm�2",�4`���? �8*1�c:G@,|�)�2�����X��\.�/�iBº����Gnh8ൾ�|���h����M?�9sA����:���}�՟0}��!��_��h&[�N�ק��ط"!T �ת��N��bR��sT~�T�Y���V;R��h]�Y.Ǖ>�!^�N�E:Qk�SD
�^�K�<J-�m+���%���E��d�K ur&t��w��l_�<�Ӯ��&�W� ¤��ZX����F��w���*�����_�C�M5����7Ț�'��,�D�C��[�$ğUJo{~�ܭ�iW*&�5�����U�u�i/���w�% ��:�9���'5��:)��d Wy�6?�z�)��﹇������B|)�П�-w�*� S�����_�i^­z�i�:FH��+Ub�J%�O���i���w�)���P mC>-4 kX���ߚ��<|Ƭ��s +7=%�+��O�0��V~���`<1l=��H���\+�ē�� ʗ34 ,��-a�p���΋��w�i{����أ9���e�	�]�%���3�g剻?�ۘ��ގ�2���P4�O�dE�R�Xc
� �n��_sQ��d�7n[|���rYP�j�ױ��c�٬ڿ��<����W���f����\�6r��3A��fZ�[��/��Ez��4���
>�-�T>�^��eԝ�S3���𔣡�YY�d�����HҸ��WE�^qw���Q�B�v9 �k�1��$u
�_�JbB&������j=LΚ*"�	�^R�P7׌� �%~p�b�����"���/��PB@�s��MPYU�C�� g&� ѳ�|�k%u��DS�]�\g��7����]hG�f��3�m��nM���t��\��<�	��Kz����*�Ra;�N:Y�7E�9���R^x��X���~��1��ԭ%�K�ں/�s༹
.��ƙ2?������C�l�YP����f�A|o��j/�cu����J�~�%��M�P�ܚ��e���A8l�>OƳLt��{��<G��t?p}�M']tLob"�p��8�O��S�k.x��}FK*�E*�p�B JUKBM>�xj�X -��M����;�����R������K�=(1H0�|Pp�^���b�a'q�
���bsC̺JG�Z,�J����A轗b ��?�D�z#����s�:�"�S5��7~qp��4��L ��1���ד��UT+�U�1 �wg&
.���P)Jբ�^X��AV[f'�5x᱿rS���6��H�6�/	ǍOۧ��GƜ{�*z�Ҟ��`��3�%�o\3q.8�de���U�i��f�I� �lN �
�hݣmmct ����l��P�%Of2_����\Τԣ�P�cik0$�+�e����n�6Hf}<��FR�m�?c������J������>x�p:��=�a�l%L��t)�WV,/"@72W�����ؽI������8�7�^f�?.�I����9"
����9/u��݃.��E����U�YO]k��M�%�p��?�1�S"�d�:���m��]yF��!pN��|�p�M ��Z���=9P���A��ȔVK�:�mQ�l4��3�B��L�0�����ݬ�<d�2����=�p+5�Om*֌��S ��B��h���{��iB�n3y��7^W6��Y�[`�Ob��C&�Se|m1_��Ҧ�~����W$�����!�Ǟ+'��=*���,��p"k���ȸ�OÇ��{0��?a��$UfH�Ӣ���+S��8��Hg�ˍK�j� @3'�=��\��{S�6:Mu���jv��x:�4c�M脨^�ܔkL�Oaw@�[���O�F.$J���}�C  �f-�_Zk���&���{[��]vF<r��ii��S �����d5�v5A�oy3ч�|}�SyщK/qa�Qo9����ι���٨*�Dapa�|�;C���EG��BX�� |L���c|�;�Ԛ�^���i��6��Mz���L7���Y&%6��`�VX���=�QgG�X�./�-ۆ��L�E�^<�A���� �5@����[ ��gn�u}_7u�GdͿ�^��(ʽ��5����R�G��ٺ��)�!�9/�s:~7Ot^�|F���0��K�90�^i���9^��uJ�u�`�q��� Ouɮ8cO��V�s�69aA"��u����ڂ�D�F�w����w����iП���̺[�Cd�6�QO�J_̖��r$�
���d����ؚ�a噲eZ��n�7�c��5���VV��(T����0��[��X�.�) ;Y;�vsu�pD�3O �>�y^�v���t��i9Y�-Ã�w�#��9���W��ccR�U�z��k�S� �U
�5��2�)IDf~�#R֕�KG�dIǇ��΍�P�i[�Y��L��=� 9d�A������C�ʝ�)Xe*�5TR��װ�+��ô��՝PʌS*���� |#��	�����r/��-�q8�)g}~��XV9�}��1���%0�z�EI��;D�]xR��)�D�yϘ�$���.�����`%��xO�!�(ʇk�S�E�堊j��lpb�%�h6�'9�͋NS�!�����҆��MLٺ
�0o�h����{��>��;�=~���ӊ�/�1Wgop�Mn��*1���t�A#FHyߗ�"��	�\<Z��4^q|Z:W������M<�?���f}9s'�ؕHL����L�	@`�+��)º:s���[�/=�������IO�˄�x�`�g�cHSFD{�)c�P��W?�<����Ld�Z9W\���N��)H�1�F�%�ᚩL�j=a�<%22V�
���C���؃d�1B~9+z�?���� D�|Y�,�bW�mX9d�Vp_O�
����r�̉hq���)�Dm�}��c�iX�7~8�1�P2꫑¨x���X����V�z�����",r��g��te4��P�w�o@Etf-��M�[�1�qќg{8������ţ,w����[�#���|��a:|	yF��v�`�F��|!�*#cI���]m11�K��^���0�;�,Ë�@�����m����b�[� ��Pq�f>��ӌ�|U��^�+�[#�N�i���4��x8V�l��(�c>W	5��o���l��h�U���CL%��I�#U?�.���V�ߝ�q�����v���������v=p~E�gi��gE��6��7h8������\�۽<��!/�t GU
�|3Gf�H���S�69����EU�	����e�(�Jo��?H9��}� k�.��
ܐM�HC��xq2Rhk��ZȽ�ec)���E�	�ہ�OK�Qx�[�Ÿ��}U�ݸs,�s.�|=L�f깷���H�)�^eJ}��� ����P=�5Rj���5H��1P���h���
3�$��,%�F�-G/{���Jz���8'�(�c�(V�c�JL+�`q!���J�V�s�Nj˃v�WOe6�5TZ���k8M.t��pP�߷�8�~([�b��`�LX����s��8>mT����"PLm��j�ї(:@�B�)��.����q�;�~|��z��M^�Hj��.Uc��(��;��Dɵ��@	��V�%��=��,$�*��=�o"l ��<f�Q9��sv���uZ�d�5���?|x��Vzj�g�à�%���U��Љ:i�� �T�����J~u�Ɂ>���
�8K����ϱ�ܳ�E$��AU!'+�`�H��5.Gf_����R�����fnUR�����u}ȨU7¤�z�b�{�� B�&DG���M'�d[
�'��\Fd�*Ń$?S%%rd����G�D�<�u��@��pq�E�oh�q.JZ�
:�3S�?�r�l�UZL�'\@�Xs+lLև�ڔ�9|�z^x���SZ*u�!�o�Ш�̻m��X���@��{��7��$J6cQd��f����\�@��X0Oł`�2ُ�0\z�М/Vat��z�-R0�#�ɘe��>@�E�Z��Ɉ�^N��Q��J����'�E� ���#��wu��o[��b�W��P���7�!�y-WHY`��?9���	��t;.�:g�9Z�u�(-Dr�#� �n�tհ�}�ι9�0�a0Y�?�il:ώ����f�B� ���!�:2]�_!Cq���g��Y��n�Ғ�uK�t��Ϡ�/6~u���BA������K^Ow৆���w6���e�%�V�:Iʐa��CE@�.�Yz��_uf�6n����1�>0>X&�
c�B���]���7��d��(:e�#g���ݛ/k˅&Zs�>�����'�`,�ک	D:����Lh�Ů��Y����
U���((/�g��9HL�8�i�ž��x�c��J=ӄ�\�o��z����L�[_�+�(ItO�"�s�h���/��&-�r��lA�?0�R���$����9l�W��"md{gf�Ё��������l#D���9�����bV�H��Q�c���7���ث�n����6C�ݻB�N_u�	��'�!M�n���2l���c�d|�r@\�ӫC�0_e�Q��]�"KI���گͰ�Uۃ?��fWM�Є�OB��e�����[�͸Q��S��{ܠ�a�4�1�pz�qut���:(8����&��ɬS ��.����9Z[�G�M��) �����7�w�(�b"	{�7�vI���4�f�������a)U����%	�G�g@�翀P�z�n^����8�m��Q�j�"+��S�3�N��z�$�}�!7��*��"��E��]}0j��w\e��O���<T߸C�S��y�.�yK��c���"9��䛯�m��qg����A�Y��ܰ#WS_�-܆1�F���y�YQ,.�Rօ��g��3�Pb� ��6��~v���JG GeWq6r�pY�H N��0\����k�G���i<o�q���Y8�4������x2�*Y|�9�P���hd|~h��>N�B�	����~�"r���s]��?�M%&sU1!9&Y{��?�Tg�'�䬎�~�HI,1��C�D�*���L�u9C���;�C%U��~�7/�%�sg��Np*�^���|f��D&��'��Rz?�� ��R5�-�X+Y3j�m��t��P��s��(��b���ɨ� PV����"^\4ҟ���!�=��M�u�*�m� ��J��˥Z�(oj��p�Q�b�K�4K���F�3P�L��5HIJ��
��3z����a@X4�fv�5@�i�Oa�v�V}B�}R�l�S�/�����u�,��r
�O.�'R��=�հ��:��A��/�++6��%��"����~�#x���I7ϸ�XX<�x.��������`*���Ɉ��}�{����]n�1>�>� ϱk���w�z$�I�'m�������YL�`���/�w;ёx&e��;�s�1w�g5w�B�[a�>�Ju�սtӋ�E?�ވ�b"8js`Ds�T�k��τr�g�ϒ�q�`U�}�w��^�nn����	+yD�)��i2~�u\D�@�A�,r�ȃr�ʐ*�X�L�P*���ktH�����h�WYB���d��B�,
η��ࣗ�'��δ@T
a�H껝{���Cy��B@�=&,��_|G�	&��C^V.�.}�G�,d?=_=��el�l�-������M����@m�?(MK�d���DN\rD��@�T?=7��#�Y�:mq�� 7aw+g��ނ�����5?�����1�(�fc\����=p`�P�(����ōz/?_DKE��^Dş4I��'��	�ϥ��F��tyF��(�� 4�q���^���w���
���U�m�C�h��m�}a���2J[��e��4�Q ��9�Xn��= L�J�H^a6���P��oo��K��bo$��=�L�����Ԫ�	f��,���I�����~PJ7�"rӷ����Ÿ�����f�(�Ǡ��7����f?"%�S+�{�CP��U�T?��i�@`櫖��?X�(%���X7^��������#�A��g��z��y1�:j���L�$|T�;�0*��BhD��sB��dF��3�WUU�^�'��M���EA҇����b��1�Nv��mc0��Phx�M
!9FӼ�N�p��j'ɧRtUƏ~���Bٚ��F�Ȝ���;��)�����,��5��\J��'O}RFX�� �k��.��g�i��y���.�2�P��9u�Ɍ�+8� �&X?�]��͹���P�=�Vst5��|Yu���2P���,���!v� �S�h�5ȷ^��=A_��|���՘;�_4k�h�z����l&�:�?W����9�F��~ۭ�E	���@ZSJLy\�紃��5�][�5�!�g��4.���vT;�#�;4>@BD<���c	(��_�J���u�0:���׊ب�w&ǈ��a�K��jg�(y@�@�g˴�y����g+lȿ��=Q*�w�s}���N&�o;��Q���wl&D�yԪ����J
��J\Ώ��}��?D�����^�C�ʻ2���ȓyK.k�Ty�Y�M(x܁"�TK�[IQ�G�i�`���%�ĭV��B\%EV�=t�{N�6a��BУ�l��7�YZ��,󒓣d_M�	X��aodX��[;IK�~h���>�7DyY�g����L�U���)B^lqiPմ���tw�g��(G!�\S5���v���0�]�W�n�̐�?\�e�ݨ�Q�K�?O�i�k��_�%�=�;u�'�)O��$�+FG��1`iId����P�����_�_H��Z�'%�.,{�ڠn�
='�|�~1i-˒*K:s��a4Iq6�.Dq+ sm��A��˃x�U�V��V%&�b:����;1���\��Q��ΎĿ(R�7U.@�t6�ǡ?�J@e�R��� �^Ԧ,Ǫ-��gC�p���<��+���Di��qC�$Vb�^kD"i�.\���BZ�W�P9�g�Y}tp�0�ai��։��Gܻ7�{��RK,�Ы^F��,0��)�A�n��T�Q��������B���fD�=���W��ڨrE��W��N	�d�wd^���
^�؊Q͋F���c���S���n*���Ǜr� ���!�s��x��x�wSOj�i3'��4F�GKv�0�d��F���C[HbQ����P5��l�j\y ��SnG{������J�h�2����4���x���%����&� ¬sb�Qh� ~�R�#y(%D	�y�9��=<2`�2���3w��t$�[6�/:CĪEϱ!���}O���e�=�
K
��DnYYOJ_��R� nG(ڄ�b�S�N��e�͵�y���rO�>Q�c����|��d�Mֆ_<�T�Y�1=p�)`�V_z�ѵ�p�9ҙ%RB�-�Y�����8��v�ЁAW�_���JV�zUoۈG<[�=��Z{~�é�(�攅�ŏ~��X5�SÝ��z�d*����DDǒ`; =W�p���.5���o�jl%��G�N�r-�b�Ϳ9:rgY
u$�Y�2�.)>��]O-���'�13�TM+��h�z�)�y�!o| p3�������L#Q?�{$+��e�t���[p�vҮ�s�M��(` [	v��
�	Pbqڐ۔�g"�'�Zw��+��������NM�����!23�_H��@�F`�e+�<(Xq�MC�>*�������YųW���v���95�⃻qL,y���Ћ;����v@��AƊu6ڋ϶^�vì�Rl��x>������u�&'��~)�2��6�g�Qٰs���'�X,:�q8$�X�/���VK��U���D< ����8�8��t�mZX���p8"���@�+��ȅ�{�hV�$�kZ�d���N�e�ٻ�NNSEO���X	_Nn�im6����7`v)i�䖫ȆnE�g�νڹ�
�_~<O�#_�.�:7�--V��P��.d'�VMD_C��9�X�"Y��E���dh�͜�d�B�s�{ݛ���"� ���O@囓������E����W�� c�O�t5��� <��>Tɟ�0��O��'�C�_���vctk9���n�o�b�Xw���/c�J1�T�ݰ���s�:..:��-�	w1�=�����(�E�vag�N������;1Ev���c�٭�TE��?�X�8�.����u��2(�߄Q�Z�_�@H��F�t!�|_������g�ꪖ��m���u�P�D��ٜn�PaƏ��i��P�d98,�m�/Q�1hCf�d�@���F�����/�,��ͫ�/L�3H[P3l�G[OA����y*�}�1?��P���_��d7�=kU�^Ѩ1�&C�㾇/w 9� M���s
��{e)3{�U����JC=��k�E+�Fk���~��][�=���҃���jaA�z<�2���%���uN	_k�/�Ց��)��N��l�X/�ض�Ǐ�"㎺n�4^�3�a�lnB[ee��C]�NȦ�OFU;��$����q���|cunź$�f��MS`����Π�1%JtA�}&{�
*jL�� n�0Ț���|	����.>�6cl�<��B1��&��\'6q���H���G��@���۴ )��+G\����-x�-?Fv)=���HJ7O ~a:Iä���A�&b{U��7,s�U��3�%�&L#��f���\�Y�:ﶎ@�b�@�O�'Ç^��;k���=酈H;_w'Ъ�l��79�����m]�R�{���Z��v�ݢ��ﻹcS���ft�.�/��J�
W:N�M�I��Z�XD�� F���]�����w���QxS�LW��겤���R*$@�x��2TE�J-�X�A����T;���;��8^����#�0_��W�� ���4����	|i��eL"Ru$1$�%Ɲ�C9K�N��SP��l�{��_˹^�p~�LN\��/f��B~�8PNlGp��{?d�D�)E�$���� ���c��w���K8��x�cŘ�U�D�a�j�u�c-q]�8��Y�i4m��3� ��厲���~�ݷk���a�n�׬��_�2�+����]_gg�
'}�l��t��a��X�,{���)*s�P��H��(���D�-�!t�iD'�p����h��v�}8}>��?s�󺌅�p���}g*��8YM���A�wo��.�/ȆK���]H�,�yT�\1ahyƯ�	����ĳԧфC�*Y��{-���_&�jY�YE�Y,�Jv�èa�(�Y�R�ױ��Vg@��]
7�W�P�8<"'�75!�k�2+���ٶ§�Pi��N�"X	���;���z���\!g���RW����P�EӮ�.�d� S7�R�O�����C���KVC;ʢ2嚼����[��nj�F]��[����m��C��j�M!�#�'B|���0��M���]$���.�G6���F{)�(hN�oj �c�B7z��#���`�闺��n-���W:K@��s Uv�<!��#ߘ�Tg��~�}�d�W�A�a�^�6�fR�a��z�MJ4#��x[}t�W9��>����̱z�\��Tĝ�|!u���Կ��D�JY�����`�z�H�(bh�[Gp=��g+�����1+�p��s$�S!��P7�L�aUp�J9&�%,㑍����?�*��)S�م�Aϣ��_�,̅��3���b�U��`'Qr6�<����������i�kz��z�(�w�!���E)�W��]�?vlK�,�kO�.كd�؋Y1_�gz��ľ�Y�-2�E�eZ��b����F�Df�Ć��X�#�{�bD�������%�JG�w G0�9�^5|.00��FCE�b&��[7�������ܤ�ny߿�$���Q*������H���F�U��\c��]�%`áܟqɀ0�I��L{䍷��K���}�?�p��ϣ��A���N�*Y^��yr�r<��^z��ߛ�X�I����?7K1�6�k��O�T������'e�BN�7��^�����|�|�����i��|)��!p��Js#�e� �`E�a�� ���Z�\n���0g�߂I·6h�,q��"B�i�U��	S�I�N���g�����ݙ@�r����z
�2o�<@����P�˵7�)���0�q�G\d@��4&j��}��)�t��2�@���0IX�7W��Y���S�*���E�٪�5��$�E����(�!X+�|#aA�u5��Y�a8�=gW��^Y� ��L�B���WI��m.|�N��S��*�ېxL������\�(4`�
�Mw��s�g�r�'ѕf�"�*�\j�h�l����g��{�����6(�tՄ���"!EP{V�{�t��ԉ?dw�v&"������&�p�����4L�<��\z�� ���=&���6!�4͈Q�EW�gy������}c�!I$2x_=�G:��U?����a�I�k�M*���A�]�z�h �Q畏['3���FT�5-��UG4�;�����lXwD�
յ����4��{���.�3}��*����+xxl����H���he��)h��ٯ���zAe����@^��~�.�r�a�����*[	�?3c�?|�Y+M�ٷ}��xnn:3Y7`�w�V��AL�^tr��HD$C'���-{w�{ٟ�������7�%kưRU;́�"��<F�_��Eؠ�p�.�ŵT褺�I}��T&��=�B.�P���7<��U{W�,�H��^�l������e�Q��4'p�4���6���g�$��n1>��\��̞u��4�.%��+���n?�z�Ɋ�a�W1EO�TH����h-�I��5�s��ʽ����S]d>2��!�5��߬�Nc�	�a�_��4f�̉Rf5a��������k����-���"��tZ;+�J�JI��ֆY����T�U֦�4���xI,��@�����ƽ�F��{pA�O���RɞC�$��o�d�X��%�k�A����⣬R:4'�EvU����D*�4Z�.�v�7cj��1s�7�{��x17s����a������k6�?�ɀn�}�2��;(6�Ňnј���>����Y*& �]T��b���H�{��M�\^F�y��g�>D�(�K�`
*�B(��X�~0 ���.�g�0���U����"U���_��;FE�8{!��"�F��J �J6����V.q����F�t��v�� G5,��@��uܧ)5�]u���QR��m�}l��Tz�z�,��Ө�HGX��U�����r�R�բ 4 T&_�\nz>���ֻ�TI�@r����Y47�˳D�S:��\ū������w�.�#/���]�0�<�&qn������0>���?��9M�F�qsY���z�bO:�=G��-�����L�G�W!႗~��*�������.��?P/�_��A��J���e�<��tK�0%���G�� ���"_��k�)���8�3��Q("����N6?W���g��򮵩�۾g�Q��_\�(��w�U�[�,�Mnx�B��yޒ�H��*�]�Vh�	l�v:Ų���D�M����K�V�[�J�@h�����d$vj�&�[�S��8>A!#��ĩ�~qķ��F�7�>ޡ�&¬%
!!���Bb�B��#���fd�
�������u�i)�2��ޏ��:&;S�l\�z�����)�2GUũD�d��`:Zbp_qB����".���A���rf)�B
�k����?�����V0�u�n-����yF Y�ej��K%�䍸��`�-�����NݸWd16z[�PXwS��%��-%�\;@A��a�R��` ����-\�Z���-�˙�e��c�{�m�E �ug�׹��Rٷl w�K˦�O���K҄d�eE�<J��<��W:M����OM�/ޠ�
�X(��0���J���L�Ur��
G��5�_!��J��"1pk-���u�{��3�,���S�����^����p?�mY�jz,�.i+>$�&o]�C�w�c�3�� �2'�;�0��J��!ݨ�e�6m���d��8��l2u���S>H�萄>���J/5�W@N�4j}��V#F8P�I}��>����i�t��2�����+�b���dAebВgr�#�6=���>�AI��W��Oj�_�]���s�P=h2c��:uЪLH�p�-VMS��'��q�ص�Ǹ��x̞�b%\FX`���6�T����X)�h�p⼎�&(	�v(x��@�u�!��92�2�S�9�����:S�1��A�v�t�ϫ��H@�o�-Li�L��-����	�/�$o��MO�s��L�����h�[W�e��<$r��qW���<`�ro�(]�*�][)P˟�8��ƙ��ˠ3 C���0�Iӳ$��b[�A��z�6�edi���k���
������!�8ZR�b,\99��t���F��J����u��6fF���ٗ���5��r�HO���)��d$i�{�rqZF�K{Kh��D���1��#�*hR@]I�G�酞�b��b-(�;��x��>{��ͽ1u�.z�*Ĝz����e�[w_s�MP?$���3�p��F���Y�Ւ����mL@]�j�݀����������yP� 쁖��Q�kFZ�ӺE~Ǘ�)d#��p�F�/l�c��F�z[�����f~VF\ �2 �W�G�I7��_(�U��/Ch�i�ߒ~h�jXB�Ľs?��]aOrQ��l�,���ܮ���9|m��s��4,�H�C��l���-� :[�.���;����o 	�a s#-0]����Ad��M񆾂�:Jۆ~�ި�@�Sbt_Ъ�Ar!ϷY���*�
;�7�a��I�|�:�pq��K8�*F���ᢕ���T"^�2�~/�k�Md!a��^Jl�JX�櫶OV	q�#�̅���� 	��X��l>�_�b��S��`�2�]�^��U/^��4�M�:7���e�d���!�2K��_�+j5��66��<�;&�kP�����fsX�P�~�O���	�nl�\��k��&3Aa�ӂ=ˋ�"�yE�La�c�����u(��i�c�B4f����.v�@E��W��
�*�ǽ}i��6⠭��*.��;3fTA��"4m����!�)I6���|7l!�ke �圶Y�4W�2�x )W�y ��i�Z��TZ+u�0�Z��=}drn��l�p� ��m�ฟ�h���=ʮhd{���\}$���.����/\@�f���j޵�Y�D�Ը��6�Ն��5}qZf݃2�ڛ���q�xe������كPN�x�+�4:}�w�0�t�w�&���x~�+�@�k�WT�.9\�idN�w���ی[*�n�H�
��E-Yws�=�`v�l��.MS��>G����FS:�~P||�0:a�Kb�*b�.Lз�*pm_�73-�J=�e.��]��*q>͟/ ;L������Mx�^Z���p��x@�l}�Uo��ka�
�Y�5(�=�"����@��G�-��*4ȷ,
\W����,�H���x�_�4�[���:#4���s��:���N5���iɅKxT�qYz�F�e*G���Z��
��]�fCv�5d�9�c�?�-�0�qx)fOl@��%X��m�<�=��۶��v�7��~�F��AH��,����4�@�E~��@�#�,ϓ�:٢iMV��G��4h��]P�����~��HR&8�K,���~�k��/��Zc �RQ�!�d,ӝ�k��B���>�݃M4	D��}~���N���0��T��Hy��NWhw��_�e�y�����+���Kg��E���Sm��ה��>_�,Дvk<oU(T�7i�w�t�6Ap���{��4$��t�ap�,�plfK�t��r��nF9�:��=��27��c�x�������o��0��'������z�}w(g��x���.K�6�
��MWT	�1���-T�����s�]l��l�Zh=�NwGF�g������&a��"�bIf᱄nP�l�E]�h�5c��>4oy��`�&�^87�o�9�sO𠲑��®ʍ�L����_�� �-@�i��Sı@����D������k:zj�(tՑ���#��.Vؓ2��J��n�w��g�l�Jv���n��c��輲���h�~�D>�
��/�9lw��x.�i*�X�?Uð&���9[�GXD������,3Q��p��M��Q�=q����(�R5����94�"�S�	�*��	�|����T�PQYyJ���L	N��kt[���3I"K���9ؔ#�����۱�A)�o�J�.���M�пǊ�mǄ�׺��X�
�{<�!���8"���.����ܓ�9�A:�4^�mDx�i���3��-��!�$�q'�LXA�N���r ��Ĳ�B"�h��]��hG�c�4�a�	D&�}��H�i��T�̄@�v��z��D���M�ʘ*���a$�玽�uX�T�yY�f�(�l��;}%��b)��6�T�K?w'<'c$ U�/�h���(��ݧf|z�v%!}^�`؄�/�Ħ�������Ko*�*f�{y ��uJd��X�yG�[�V��[�������6�S�.큈&`�� ̣�C�)���}���I�g�2�|��� �{N�G��<*~���S/y�F����jB��?��H�٥����;���r��z���6���p�XO������Q/c�@�b�I#�6{[7�o���Lzٮ����W׵�"��{|G�'�!ษs-�����A�}��S�<äH���Z�nZ����.ʻބ��yI��ӹ�"��%�.{p��A�.~#�=�Wٽ5_8Y�.\�<	z�]����Z7�Sc���#XpK�����]%װ�7Cm{��4L��j9�4i����'_1=�T#�:�N���m�d�M������������^3w��pBn|���S�9�
���o�r~_,�?X�S��V�d[
�^ ԣx}�	L�K(Gԟ1����'<7k��tkǃQBTc=4z��/�w���_7Z��`����9���bPhGf]KnL��{�#��tW��U�˂5�$� �G��B�^T�����j��+ge���pF9yF���]�B-I��e���Z�<^%�9���D#�_:���[����})�=] rG&ʵ؊2V"��Y�L-�R�C���+Q�r��jX�>�˿.�<�һ%���xy!n�9����^�*��!.���}����Y*�I_����d�ӥ�%�{�%=�w�Kl:aѹן�����Ƴ1��݅��g-ov���,��d�*P����}݇�=V
ٯKMPvF��Y����J�,Hk7
WB�Ƨ���N@W������[������ w`�~NI��4��Ɋ�Na9	��n��OP����젤D]�G[���@��YEd=,�Mo������|���o�nKT�P^"i7m �$�F��ř3k�/���'�W͛� ��V�Oi.0��R��5�/��x�5\�xȓ!�!g�"WDf�����OY�q�j_3��h���}�:��8��~ⲃ�N�Җ0:�o����D�%%څ��$s+q��I��M�UN�o!��M4�pv�.���æ		����&��-$x/\��[ N�q�v��t�U����F�?��py�f� ]��d9��>�K�2����A�_(W������O��QⲊ+�3�(�_u>4m��Y��cQ�L�v=]�Q��Y�6F���@��U��)z�e�e뽈cr*�͗iV��4�ib瘄�C?Ɇ��b�7���u-8�I�N��}�Q�����6,��_m���+��3�usDZ��g�x�����T<G���y��~��_�"����^��#�����<_Q��
^ç��ͬHlMpiH�)6�'�F\O45%�5��P�#g�MU�h�ȩ�J�&��y�j�m҈���?r�#��2{��7~��;%l/��m�̩^��׮���g,��Y��
�m�v)�?q��΅dF<"�5�5�Yj����C@�'>�G-R�ν��rO,�<��v]J}㦊�9���X�j!�5�;ǻX�6v��Ve�Lx�Σ ���yR&#��Z;"��n��w~�W��k�U �*���C����s���_��|0QJ�}p�U�u��~��vҖ2����'��� ��;G�K�@�Z�"%���� ��E�s��
��\�P�^R?��geWu��1;�0�^	�j���REy��/+:Υc.�i���3�L'�mB�f���a�R���Fg�]��,��uZ�򡜳���nľ��ҁ���g���/r&�A��O(� ����#��!_XXo	#�A�����?NW���l�j)�hE��bT%�ʂ$.�w5i���]	oi��(^P��ͧ�Sau�����Wz�F� ��V<���T���AC��fa��N{��u��e�w{n�[�����u����ژ�)��W�-��P��Ӥ��H�..��A���P<*�u��ĬG!w,�?�-�)��=6%�n����'��J{��H%��s��j� '�0d��WnΨ��m��:0+N�*]En�#�f���<�dQZ�f���f8Pw�~�bM"x�k3�PR�X�;292���C��y��JU��r3��	�^��i�����Y��r玴���2;�@:D�#]��H���	�`Rʊ$���77!��#���rxW�*�����c�"<����os=#�ɶcCu&7�L��Gٵ�7,�=;� �A���
R��]���#�Kq-O�C�%�	�r�h���4��q;�P�/���E�fJ�P
~3�|[�q*�P�h	5��[m�[��n��f�"�2�]�&Z�k��O�s����1�ߜSb���26����ި����FݯZՓiq��0}� g���>$�a,,���l8J:lB9}h�
�D���(F��k�����5#�;�!Ʌ]�6��"7XcjN�����gx�.�dPI�I�"�`S��J�|��T�fR���K%�.�8�J�i��~]��{t�2���p� ��]��Ct_-co-(m�<�#�Et�
���}@%Ӟ�qq��-�Dק{x� ����Ğ��L �^'R5ܿy䵰���I�»�=@�it�s�'%���e��El�%�hnp&A,�c���պ-�h��Qs��+DǴ.3�`R���b�e�݄�3o�������^̃m�ѭ�[촔X��CZ�C��E�:���AO���!�Lf���$���.��lV��,(G�`��}%`=EU�E����f��wj"s��B,�?����뉔Y@�Nu�������y��� ���T�x5��No��"�a��-��Y��a�i���2r����c�>�PY�l5�w��O�NIaƤ�E{;�#>�v��b �8Y���@�C�E��%T���=��j35�my�25�Z����A�o�E��M�����nX��ǯ�	' a���&)���T�G���v�w{k�l��S�绚x����q�|-��-�V���h$��0[��\A&�9��������ޛ����-y�mw�����jȻl����v)�/���*ƘN�i��bJ5c��Ï��"7���3ȼMs�}(��
3cw�����^��Rv���^T���v.���-,��'���ժ��Q0p+�t�̫ܴUo��"�'����ŵ�l麋����w�a�x��6eB��͔>����~-���l��U�k�"�!l�ԭ�Yǹ�OD2��e��y����B.�*pR,��=��d���B��__5��O@�T�Q��H��_G��O��[�c~�z���K�Ka����%B b�t�0]�)�� ���pU�ptvq��������uxE�қ?.O���2�Mu���5���$躒+.�)�K=%l	d��@��@EU9ēA��'������9����k2,8PG��9�Si`&�d���k���o��&����c~�Ӂ�O-ôbۦ_N�EM��4S�\
��f�.��Y0nl;}��=P�m`n��4�E��G[D�������I3tj>p����Êt�⟔��� e�R
=�A�I��p=�VPP�[���2��#������/�?^:�,��#��5Y~���D*sf��p����^`��-�0��ה�%4K,�ˡ�c��MReV�5Zc煀>��L�˰��
���nQ%�Xkx_%��U�z�#Feadu\��L���'H��!��!���,ў�o�~�0���3:��:�i�#��j)[[\�'��U��q^ Ј�=���Z�G9d*;�z�s�Ľ�o{(��7�]d.#'����"h��r���E)(jw�bw���as�E�0�#�Q�&^����O��c��?Nf��L*�&�)�"��k1?��?-��j��2��$����U1���x���3p��P�BR��k��%��9�R��`�܍����
��%�QkXsS]�((�QvG��x&kG��C��h�O��3�.�[��ө��,t�$��y�YW�"��=��ނ֯3�՞YTjQ��}ϙJE�!p����|�w+����p)�͝բ����{���4Cb����v��蹟�i�%���D�ٷ�WE�}z���)���{)�QY�t
�c�)ۋ�OesD^b�p{w��%FlD6�����yh��e˓W�ВH��{�FIm����ۅ��c1T�S8�^���ꕤ���i��#@ѣ2�Ѻ�Os	Z{v���,��W}W�ɹh�٫���dC4��Tv+��+_�A\,Ĵu��h�� 8����mk�Ԃ���&�����Gq�ݐ�b����́;�*�m5'O���te���X��9�m����=z�]���e!�"��긌М'�S�1��0�y�
�
�� "4�G�C��U�����p���D��x�x���������PW���Cm�Q��{�CFtA-v����j�>J���FM��;��|Y�uK��a�}>���d,�7��������/%i�:"�"�vCrǍ�e�G*xU�r:�N�:+��S�1i٭?CBcb��(���l��>KX&��g=��Qz�T?w:�3�hS8������ �L<y77��.u��%)�~���>_�֛d����q��fι�*|���p@'=򆙏�o�х��evܿ�?-97}))����5�~N5��l��SFx�&|�{kۿާ�=Ŀu������S-RU�L��-D���m9�P����@T� pj�ި(���Gϔ�o="L)��Ҭ���p�)cF���λ��Ue=�Bw�����"�kJ�t@	i��rC1q�B"'�[�eg��¾�ڨ�#�)��0�%�������۷��J�F�a�v=s�LhH�/dx ~�3�p#��+�4�k�K��t��;�lg+�B��
ck�C����g���r�!�u,�5�O��^6.��`��k�-8�*?
�����ߑE�v"Y�֡��f5��؞wΗ��i����>�{��L&"���}*~�E" DN8�3� Q\�4� ɇ��f�F9T�D�������6�6���q�]�� �J�+�:�U�J*W�lK�腼�>�I%����h�ÓEuH'D+F�=t\��@T��������+<�1�d,W��T ��,~��va����tԧ���[��5<Z�x�H�k�8�t�8��.7��uN�NO�%�Ia��ְ�|s s�S��pf��Q"�z)	 ��#���Dw�>������U��LV�v�%�l8�A��5B�P?���N�� ���E���SĪ�ܯQ�i�z����g������p��
�������ƶ��z��0�Ej<*T��P�XD�����+�I(Ƒ2R_h�;X%� >���>0�Z�L��t$�]��V#: SV٩���p���/�Y�N�zC7'�'�Eo�q�Ư�����F���q��e�������#	=9�$���ZOO�o�E0��0·�L+k�ɂƛ�����m��� _{y.��#$>�Š_�^��=��f �1��!B�hZF&�[1��4�튟��f/�>�1�n`�`ϔa�5x���	r]�1�סX:� 2�#&&��˯'4Lr�[����-�b����ࡃ&Y��e�w;]U�,�'��}�M�G,�V�M?�k;��oõ�1��������'jz	o`�gv�����"#i�C�Ǵe�(��`�k���?Aw8��q���"$�4Ī���qő??���h���)o��G2;�ŏ�*ނ]���*,C}��hqG��J���-X#��ɣ��+̙S ʩF�]����>�,�������kP����#+f��yN���m��[@6�#_TB,��+�מl��"-��
���b>�6kt�6E��]�[
�+Ϊ��[ghA�������u0��`ȘE�
�M$�=�N7N����s	��#i� �ˎ��]o���o�{���+�YB�Rk-K:
���HP:���A��V���I"'�Z�\`���4�*��d���D�Hy�)�{wca��/!jU��A���W�t�v2+��ү%5e4�]�g$9	v`������|4V1��Dή�h�E�K��W�%�K��|L�!�Zw��T�]�x!?:���?P.��ÏL7&�9�����4�jǍܨ�@.5&��<3(ur�تO$�H�NisJ���׭5V
ܢ�G
��~s�Fee�-=����A0F���H�r���b̆��^�?�.�&�w󘧶kF��<�U1�e��. �x%��� zK����!:Gj9�^�4$m&��iߜ{|/��������a~��(��u��q�DD��ą���wq��{��l�9��g��I�(�þOwj�A�ٖ�~���tQ��qD�Rj'��&����ؐ8�6G$O1�
�Eġ&O�A��dә��:�xN�O���l��㸆*�H�E���G�w����@�(e�JXSB��&��ri-U���$FR �+��о�j����Q$ԻM_	�9Z�ųb���?>�&F�E��,5�ss��7']!��c}𚨥��hO�l֬Iz Lք(�4��*8_�[��cT���E���^�+/Ks9Fݏ���VXU7�<���?�'�j�|�I.I��ߎsu�k�mc1�f^�}��M�y!��j�ek����&7�W%Y��f4X-%�7{Q���+�����k�rۗT���Ӧ���gr$�f[��f���q�rL�ńg�m:`��îV��%a��������mn@��[�Rj�V�������L2�/�������G�P��nIH���y���0��3�sdOG�T~�څ�<F����Z`�z A5�k���~HM�W�!��i�*��ͮn��}+���a��v!6;Cj���y�^�|�!�GJ�^4�9�Nc����`
'��\~|yĩS����G)�f�D�:C9��z�[�h?��-���Ҕ�+��/;�D6�`/+�yB�՟su��%ϵt��h>�oS"��Q�`�1eX����Z���c���?�"���f��}\2��ީ�	-q���Y9�5�n���>o��2+�Z �w
�3_?�'7��	�E��H~�y�2"oX>�o.*+���ϟ������G��UN��D� #!+	��)����JHk�e}RӅtEp\�E���x&�b�t�_����(�D1��hogx�?����h����?Jϙ~8���V�m��������L�O���B��m��E��F�Y�s2_q�e�*5����t�]�����#z��F�qX�n�s�1�a�=T�a2�#G^d��Ƈ��� q�k��g�D��屻�a-tf�+ ��[�O��M���6p#Y�K��6��t�I5�Y�H��B�C���dh�8�F�,���@��Ѡ�H&�E�b6���N���`�-1rFV".�Հfva
��7�x.HR�q8�k̘Wz���J1�EP���c��"8� q�@��8�.�v��ʐ��P?��-�|�$��.��7x�Vb�k=�Y�ǉp@>�̝h����:?�Wt��t
_�B�m���j��u�{�W�96h<Y.U�*���6�.�)Z)z��|� /��a_�r7<����iTD�zSnQws-8���)����Uu]9_�P�g����-�$�;�����^���v���,���l�Xx|�i���J	��zK���OL�уS��3��-;�ᗖ��$A��� ����	y��w[[���P'��#�W���`�������z%�"�D��;�`:'x')����H�J�J���2�u	-N��h��y���mMS�x٫y�k+c[G�Δ�(����`z�v:�-��O\f9��;D�Z4v�C9d-G��o��\�bk�?�^���")�'���0�A��d�(љ2�}�x�߇.����b�-y����_���4�}p�C`�H_ƈԸ���/`1���NG��A��	��vl!��<�}�Zk{
�����an�)���w�>�w��	p�%�����'���Iv��$g����0���&|��i��&ޓYx�ue0��?q��Y[Ve#k f�iל�Z1 [)*GS��1�<�ˋ輷��ֵ�GMK� �Y�x,��ԣ�#@��{�5�QW�@z�F/�$�� >����"���Ą2M9�
P�&�&~�Dxq�͂�Y1巊��|S�}~H��Ez88 ��gTA_R����#a��2�Ѐ����%��������_�~�݃GC���$�ۙ�	|^S�?��2o����V�Q�Mh�?��G�FJa�7dN�P��4��J?l�U����N�G��+4ihV���l�u����'s䃤�2��JwBՀ.��o��+R��%�>�t�e���"
'&nâ�ӭ'�Nء�lKȤy,����G����V��LS<�#���xߚym���ppO(�c!�~!K�cO/c�Ŧ^R�c�flLo�|&]A���ų��VMpH,~3I+cHJ� N�O�M�	�*�vd���Pf+���?���(M�w)����gj^��(}�TWq�ʠ�pC��3��@�c9�f� �!a�!q�Yx����L�ou����5a�.hJKh<j��Nb�{L-���g>��ƛ1�9�u\-��������-Fڌ��d�t��2�qC���Jo)N7���xs]gI�������mTO���~�����E�>�s8L�։����gPa�+L�S�aY�S��'�����m�g��в[��w��˰��Z��Ms8���b��0�U�ڵl!�=iD�%jƱ=s|���Q�Fp��E�U_EM�Z��"��xC�y�D~��w�m� ɥw(dyf��i��ǮcO�M���P*g�ĺ`�K�v-)��Q�)[�;��wR�ԋ��wh*�v),���k�=�sY��5���_�y�~%��;h�m>��o�#�>"tR�~@0�b���0G���f��M�<m���T���,3���rt�ky�!*O�*D2�S��.�����]�i%۟�1�Kg��M����H�2+�I����k�D��	�#X�a[�I[=�3��+<�J�w������њ+�J`���Yk���,��|�pTt���蝴���rZ�ۦrn�'yA�T�c��J����~9S6�&��:6p*.��L�~qʦ����sF�H�E!.g9.���b� ��*k��|r�Ő$�J' �
��А�.�,��9����m^L�+d��N���cW�����^�Ґ�J���M��l�TR�tbY0"R�2�V+�>���<�e�I�BO�w��r�~����-�-Ko��e���7�(�)Y��Rs:ܲ�1�b��}�P�pP���h9ŇQs�{�-�(�h]��� 
0����Bs���UJ���®4Dr�=�8�\`��׆ Y:Y&2��8�ô�GOb�+]�`��?gn��q<��V�T�Z�챐}:��
˪�sGKt�QȪ�k�\W�hz=*���<?�[��z|��YͲ ��9P���}��ʬu��t�����Iv'��I:H��N|���8���D��4e;���(�F?=���k�z�,z���> eyt�񐆼i��$xG��Y��F9+�iBr�!�Y�3�/�Lk��P�K.ꝃ�tQ�>��s���`J����%"|����o��H.t�1*�3E��1ל�jQ�t���5HJ�2�/J��&L���Qy�Rޣ���g�e-Ȅm�봭@CAĩ¸��B�eΉ����$�/�o$��P^ⵌX�oSCQ��;Ѕ�l�ٖܖ�L���h��|��@:c_!u�)�=���Çז�0���v#�r'܎�{/�N�m�=�h�N2�{&t������mM�=�4gu���]V�S>ɂ��or�}y�:�(�Q�N���G�0rW���j��	4���#�,���_{Zb��k���*������v+!1�z�x�y�	�y_�����e���Si�#^��!����$��xR�#4�x ��O汑�]���e{Ζ��!	�Ƞ<���o�C��'��dl���OD�C��eXeë�:����3�y���r;m��ٚ��D1�7f]6h�݆���v
 �Ha��x��u���;E�*%L����Y��o$�	�Xm�1Ѹ�B���i=�ބ�7�@ת��P��ʅ��w�PQl���1���޳A�?T]� �����!��w!fs4�#Н��'� ���/��v[��v��h6�;�4��jp�I������D9F�:����%Z����E>������׷6�;��SҮ�#��2��Mƙ�h-����j��2EG^ܐ65_ܑ'.	�y��;��k�����Q�=����3�lׂ�b�5Kb��j���B�����+���_*M{���k��ڴ��bjp�?3�����_�|O��.d���3�ϡ� d����g=}�pj�x��L���,U�o��d����ri�����1�%��=�T�"]b-l�`a�UהF�Y �U���d�|�T���͈su{I�l)�����IqY�\;�w�I������+�	�Һk7�u���T�-��m@&�E5�~n�7S��"�IX��Ct��ǝc��r�3ʢ�e�e:U���d{�T�^]��.A�%-B��8�ܳ(n�NpQ�*��B1n8.������X�yg�m�\�����ŗ����<l�;��r��Q�"2�ZA#ze̟�hI�UXC�Z�����H,M#De#�v��zЏ)#�T[�R���x�uy����SÉ;uz��m�(�߰����q�eH��\n�`���m]�8����<�5�$�"pL�J����	�)9�nMs�D�����B{���f]�W��̵��H&��1y>y�$���f�M�[~x��{�҈�<�*��o��!I��I���zoRk�O�m<pDi'����G�{�"+i����^���Q-����,ם9�m���N�y������r̯^�Zx���	�T=���"�#���n:j�h�9�Tf�cu��sh�\z�n�tc�O��ސ��� �e+�H���A�J��&pv��ؤ�Vj���¿�A��6p?+��E���妵�>�!�W(o#JқP�BGyH�D�����)Jkj�GB�rS+w,�1MH�@z5jTU=X�BX��#�O��$W��Ճj�t]�U���wY�=~�>b\n�pq�:UNe��������҆������>#��U��
�����L��r;<G��%��VK+c���-�8��7|@�JЇ��̪�<W }���N�ԕ[��.?R����bd�!~�cX�J��Qa�ޘ6��Fi*������.��_�zi���~k�8�@'��aLr�1����"$� �?~N��z}���5M�U�%*Z�+̵{:�s�C��F�k��c0gҟ�N%/!,ql������`Z�bs��:���b�dR�E��a�����'*�v��Gm�J|~x����ԗ�`�g?�;�`�H��m��>��֩V�3�?j��dN̔;G��Ñ��$H��,y�dT{�i�Zd�d��}r,�a߰Y�`��k�U�$��W�`x[?�h�ht�#�	ث� ��s\MPR�?�-��c�����ZU_-��8�
�#P���匜W��r}�r�f骀�1֍�``h��,Д�Fr�`�)"�u��u�Q,O�*7o9�3�D�����h�mg2�Hr�&Q�^z]�8h���`�[;���*��[�"�ޠ݁gZ�9d^5��:|��}�����x��)L�g��o���f�����~eU��<�D=�؇���v�RWT~[D�/��N��U���D��y܉�Ҭ��:���t`h	`6i�����(���#6�����Ո���|4Rc}���)=)���<��o�cT�K!����[�l�=��s�$�!W��4��ՙ�j[h�%5՘c(�|�#�o�.�0W�2��u���W`�x��?�����G��ͪt���5Vr�V�<+	V��v�1��|�IG�Ll��#�n���F��Ӓ~0=~o�cN�eS��Y��ۙ��[h�R�2n<��?+���d���q�y^J����)��#ص�jjL �Hd�Ye�~��m@�e�<m
a0�d߻T�m�'p���q�1��h.;���9���՘�nc�Ur-�v��"�5����f�b]~���ֻU8��nP����ڰ3Y��ݸ0Ư$���t=r����zx�D~�\6XK�@o+��8B%Q34�@�����m�\C�]۫"/bX]�@�P�Ȅ�?nVGT�����J��6���f��<Pǟ7
��y�ڤb���=r	N��-��-�7Ԥ>M�w6��#�k���7��^a�kdr��W`�vY|7�ן �[��\� �S�n�{�P�b�����Q����ꖜK,>@�e�/T�����D^��,h�xG̢ i�7D&��	����$-ٗ��<=��[����!�v��ݞR��m��k�,nb��wŀZSs�������e���o�� $S��l��/.�t�?%�:�(S~�:h�fiR\�'*<>�Yje�<LmN��(�䆡G�:��A ϝ�v���P���_����1���+�X��*��B`�߽�l�v���?�P�D��Đ��>��R��ވĤh^��*e�P�ܢ��&:�I����Jʡ.�����"���]8��A|����nf5�����D�,����௽��r�"�o�E��]��|"S�&�ę�n�+ ¬�V|R;���q���s�����t5*�$�-P���!�~Wp� �`A6P&N�tTN����os����ښt��2V����w.�K�
��l����~���9�g��uS��8��5��۝��?A�^
�����{���FJ���N;#Ӣ����k��f�X�"|"�`�6�C���=����]��ۇ�C��B �;q����� �]U�������� h`�����U�|�+4sd�GtxyVAOQ-�ܟ$V'
����=�M�b�	�Tf�o
8�W�PG�N�,g����Fz�p8�M����>Q�z�θ��D����]I��2ևæ�-�|�4T���7���b�l>��Ӵ�Y�`/>|�����>�6�\du{YLQ���}�Ӷ���w�d���J�9�c�fc��g�X���@�I84��RW�R�?�i������R�p�έC�뤭��3G�5�2Hz18�aɹ|�������@��6����g�!��#�=�l���3��vm�${Y1f�k"˒��^4�_��p���佭�m�V<|�ҥ�6��|��_�B2��*���!,���!��������	�ɶ��	��RR�(�[���.�c�({�R����i���u`x46�2K�%RƙS�qc�<�=���y��Iw�5� ����V�g�W?Pv���2���U�ڡ�|FSH�̊7�MH���i�Y��Y��b�͡�w�W�a[�}ٯ�};������\̾:�jٱ�k���+���p;��)l�i3���k��<�)=_Ձ��=�g�(ڰi�:!T�53ˌ�hia�S���<͸h2 43�d�}��l]?B$���g[V�1�X���A��Kݓ|0�z�G��4R����F\A	�=׿�+ݤ�K�Ư[��K��<�Hԑ�̓B� ư�9�VT�x�!��VQ��ZנZ��ТsUs=�kM��g^fy5\��w�_�r"S��0�OjL&����+� L�N�/�$����x�o{8JǙ��2�NEU��-yB�0���*�Ò��Q��,��>d���܄��T��X���&M6�
�RjY*��zhѴ�.��>��q>�l�r�W� A��2�K����G�o}�s�w =�	g`�؞y�����Ҹ��o#6C97Ǹ���Y�B�KA�OAn�c%ө���аEs����bRW�����:!^v �r} �F�Gv{
�<�aqo��L�~샰|жj,��P*��+�י���{!�z��#�1������� |U�4��F�8��; ��"\��_~,8�6z�9��1
�kE�I]��y�@�
1D֎`��(�5��} �z�<tP��i��̰�Z�"T"���Nș��2b��ċ�𶮄T;w�G� �Ҧ����V�w��$;R� _���_���݊۽d�gڴPJTz�1�`��#�	�ح��p�/P�2��SÙ.<V�v�@o�0A��h ���f�����mə������$Zx_��H��-%8P�$r�qm-��W�6j!�x[�GGQWJ�F��ǖ�U�l8��;�s����1��&�t��
���8,�����N��x�14��l䰸��<Nb�#I)����:�Ԙ�)�;f	���M�#'�MBDҀ�7�E�b��'-�C��o����$�5&B��[�i��U"��rP@ҵ7��O������{�RJ�",��d6���P�';�|aE�A��)_�R�*u�%5PuI$79��|�V��0�E�f��2ؤ��͎c�/�\'�(���Qw����w�s�u+)������HO��a��ȑF1iw/����P,������������F��v��GH��:�C��0�X07�Z���E1U���?�8��� �����rBI#ޏ��1~�3Vck�	�:�?x�G�,Z`l�ڕꪹS�]J%Sצ��^&�V�����*���a�g!��6��W�e[L��'[PP4,�ҳ��}ז����kŤ�g6J�1|6�9�]�B��V��n%���mR���:��QpS���"����/S��Q�N����eI�^ЀS���`b��ZAvd�f���T�Mv�Ȣt���Q	������A׿3!�a����Ŭ�QES���v�\�����*��wN�n� u�]�o$�����.Fb�J-U�,t��߷3Y�ar:U�5d���4�}_#��z^l�փ�u����W/�7v�G�-��o�YC��/�����.�������&@���ڰ	�,�4Iamb����?��R�c�cemUڲ}�]E-@ILI�vk֤H���d�����]ͣY�zG�-���M(���:�o)~ᰋ�7����엚�{G��,
v�������Ә:�X�Ɵ�ֵM�%h�!:���m��\��8�.��f���� 한�%k-a�JɃ
:]��q��*BP%/�UJH���Q�e��K
�1Y�p��u�A9\;�A	�v8�����`��װ(�w$��3��ө��}�і��}��.��O>�����֒��}L��Bځ>'0�l�aeWr��b!�V��z�Ղ���I�l�D�G$ȏ�ȲI^��jF �$��Q~f8��R:EL�*����z�!ւ�ci�<)V7آ��Y���OC{D/Z�)���%�4�9�Af�` &B����0�Q�h�p4���1�dw+|6�)�Cj�����T^�t��q�a�DH$��hF���+�������V�ja�i�a]�����ȳ�Gq���X�y�ĕ'Q#���a���a*�@�4���{�ᙇ��$��1�Z0����,K�ZQz��򈀪�K��*�g�u���t�A����E�I����۷�ra�㙀t��^��?g`��!��o��2:F�T4w�9w�T���-��5�vPɵ�U��yL��5�����J�y~�d߯-gtJt���=��cݴ��b{W��B&v׼bWS��?D��"��URiHb��%�<��<����ѥ�����m�1�	F��ߵ���+��*��;j�O�{Z�:i2T�Q�n^̩*B{Z{�?��-�Ԏ�.#�>�dBZ`"�ad4��5:nD������79=6���K3n>��fM`����NƵ����� ��?P�~�J�� T>��1�7���<~��cO5ؖ�=�<��?XM:�c���X������dS]'���)�`c�T2gd�o���K� +������`��א��"m��	�q�vLF\9={�Ip�JA�{��,�=��=�� m��u�z]�,y������q���C��]������~��� ��\�.��wi*S��L:cR^m%>���_nIo�����Z����,;v`��O��-�|��MK��7o����E��!KfUq���
*| p����}����i��d�
�h�������ˍ�DnE��UY�iOD$��&Y��MkSenK�Q�bQ�93��gL(y����2���H9	���ȓ�}/�՟��1O�(gf��� "W���b���z����-S���,��t�C��JB����+6R�g���e�����@�J笶�xOKwtz^�=#��rQO�`u6����@�C�(�}���`����r�憱��4�ƥ���ISI�Y�R��~�<�m����tmLR�
�#�?1ʡB+y�\�Xl���]�(؁�rUC
E�����q~J:��(2~����)�`�B��V�$*b��k}�m���
�yN�-��U���8fc�����	�_��s�����t�5�^���tDd]��v���;/ȐW��2�.DT���k��y�@ac/�"<�c��U^;Z8��w�{�T[��ѳ?�>��:��d�Y2_ڄ��PL�I����_��N�l��%��S `�R���ք��=�J�n�������x������Fa�m�S�j�q��r��ތ�*��'z�d�*�Oxh�A�_�>��C�q�K*gvl&�T�Olv���;G�O�T��!p7x���ܾ?@ӓ���pz߇�od
�����0-u,�������)B��s��O2��q�a��6�1�=��Sؚ� �y3�&^AV�*Pݢ���Oƣ�F��Hv
<���A�ЋU�r��(K�h�W[�]��S6��(|�R���G�:�RA��:�~�C�y6H�"6�{V�I�Os��l8��Y��u`�o]۬\Ly*�1������������,��$r>�� m���{�)�&�H���称,���z%��^��u������"�@ �	Z��V�,�Gݗ��:,Wr��YD<��8B�{�/��	���9o�����Oo�Rc:����Vr���t3`q9��Q�7xf�w������E���9��,���]�H�̰NS��̶�PY�����D0
��l"�D�r��=��#( F�?D �ҰM��������śLf���K7��=8e�z�Fţ/ww�[�:��j/��-֮�-�%��Z� �P�~~Ҙ:% � 8G&8_��#����z� �#���D���TQA�e��G�3מ+��ǐh�y)]5+v�󟄅�Ze H�m!>S�[J�u���gY��`L[�)���:i�w��~����0Uk�/{Ɍ�r����.�
{����^m8��s�И�����t�8���>"<}���T���-�j��e1�G%��Q�$Bj�r�B��?�4CD�|3�9{��������	3�e����X�`8��cV�Ӵ��yÌ�& �����i>K�P�]k�[��d1��>��`����U�_@���03N�g�� +��(�*�F*My���X�H|���	�ڛ��<�FѢu�Q�4kʔ�u-Mh�bK�(5���s�@?H�ܟ���'�����4�Ok`�w�c6ʙ~SN�����0
��b�Y�Yb6�jk��/���f	J�3�m����KJ��ći�����K�������y���м��|h�ǡ��;q�n��;8q��=6�l:��F���X�n���Cj;����x��� ����>"N�/��0��>�`�=��x�P �i�4x�Hʯ�ڠ�,ݦ����#�����D�����ĀU*�@!ʚƸu��e'�˺_+n��Hw��0=��)�ZS~*(�ƈ�R�@(��n ���dШ��l�07ޱ� d��<E��zR�? ��y!��=���o��9�j%8����,�\V����;�p����E?vY����&���(T��;h���d�,���p��fqc�+7�G�is��k��d�g}ܔ�E����-t����S���hz@q�R9#��)p�%>�B��[w	��kɔ�tB��R����������D�%�( Ш���B�u�H��䌫nׅ���k>������#Z{�v�۸XՓ2F����|��QT�j��]�r�����/�0T�yf��S�#f4��9�Ύ��&�M�$'�'/�1`�B��&'ڙP��H�7��eFGr��y��C��#�H��vҝ4]��k�o� �b��u�y/z�Y��%0&��BN{L$�f<&��9p>�z��#�&����M/`Si ��X��}�w�W�V�&� 5^"�5Z�|Ɨ}*�8�w��P�wY"G��_�q�g�/q>�ޕ�j�����f�K!�sjX�A7ӟ,�v���B��1�`�������+�C�\�W���2�2��9�eu[R�-U��8�}#&e-���1� ���wp�v��يX�8�0?X7׏a`X^{qnjV��k��J�&t��a�!�$	]�1Oo%Q�T����hP��s�@b�ܞ���&����#���&b2i��e[b�~30�3��w� �a�BtA��v��&I|��~�n�q���k5n�.�X�e�����>�8��G��i}�ǽ%�[(�'X�j���L����/��'����ʓ����.H����X��qg��O.�>�L���>�w͇�Ґl�0p��Ͻ��8��������5	sMK�8�|75�(/y�F�(*�g�Ԑ ���H��8΄e�-]Ժ��<����jӥiZ�<��z���^x.�b�
�����~�j���%��?%�评�	5:�/�q�U@�Xk���iz�ސ���d5�+����[�>���N���\�t��6��"���VLA��l��Q��9m�+����P]~��g�՟'��^J����o�L��@`�Q-R5TT�#+�LuTs7&���",Nu�B�x^b�cl�Z/�t&|D'ʀ�-[��uA���a�W=ЛW\��o��$�$�c)�wj��m\냛��t��u��O_�o��|Ih��K�D�H2��^|��(�$o��Y��%�n᱆��M�@����g����0�p�J�#.����C���c�Ϧ)Pٳ���&d���nv�uR��2���N'��%�~�JjX�3��G��C��\��B�,׿'x�)��+�����%�i�(��ƴ�PBB�͏�ܶ��\pSՋ1P͸G�T����G��rg�?�g}0�0a�j��ڗ3���&��]��cAP�1�z�~O��ҏZ[�-�s�L�@��Z�Ŗ�9�&+��7�Յ���ޕ�j\��* ��%R�
5'�����7v�9�S	����B���X
���w��8a�n���*�EK��d�����~Ա�!|#�W*�^�i�����rA��?Ӥ{$)������Ǖ�s�<r���u�F�����4���4�k����XA�H"~��!O�٫sl��0���~�.-�� ��zh��:џ7Z��}X��@����^f�9xN��-�=	�����|�>��C�ډ͘y�b�,q$�ڞ�gv���B&k"\q�w�QM�߶Ą�ZUq^a���vXAU��.К���/I��,/��� =-8����T᜕xk�"����a/Nm``(��K��tT�ݓ\�m4t�7ŭ�fOg\�̓K��0����ݍ8$���BG�8W=��P��=���vD%9� It|"��C�`�ĢB��F*��d��������Z�o�$u'����"�w��C,�o9 i���RE�<�8���$�~?�?�r@���
���bV��6
R�d��f��)�0�Z�oS�
0VB4�8ˑӇM��2�Rh9.�B��6<cN͵+8����ñ1�~�4E�2Z��K�Un��\���Q�,��A�0Sft�����+���BIG8�J�46q0��Nr��"b�TTX�f����D����Jf\�K}_��J"&���E+�!�jÑ�V���/�Mo�qK,1|�s��_���fb�>�,�r&Y� -H��0$�H��/,��^Uk����g�&Z�Q������*�xiAհb���YF(9���߭��Heˍ�M'|L����x��-�a����e=�]�S&i�X1"-Mc���|��
�Fչ�����0����Y �`1�Ɋ8��E�	�?��Y.>Δ��k���\�l��Iy8+��|!��3z��̹̀�"Ʌ%05ʊ��#���"hq����9u]�s3>��z.B^x��+�)w}�r��6�~^9�����vpބ���f�1��ۈ{��w�h|w��|��L���4b�?�!}7�L������&�}�IB⟚l�K�ǁ�}�τX� =��MfW�YX�ɒ�JX!;����*�;�iD� �
�-�ˬ��&��e0�;�E^y܅� �d z'�m	*i�E�7�>z�8�F�w(���pY\�[w�+T�������6�R��" *>Pk�Y< j��ܡ-~3&��"��Gr1���$���uJ �R	V֖H1�;�Q7�������}ڂP��&l��ҧ��l���)���8�Y�o��+d7ܹ H��H��/�!�Ш�ǵ�A��D��X����n���dN=���X�6,)5���YD�0q�þWp/��e�!�oFW�e���$;m�?���!Wl���-�:��3Z֌z�t�<8�	�*�,���G7m��CK�5�4�\�a�I�\��MW�y��N9�k�/�h��偬v;��I���d��W%ERO�\�R�����65\#�Mk)�m�i��;#o��&��,W�!�Ml�B��%N��9I�Qc#��t���WY�zF�>�#I����[���=6�b��6�:Y�0ghx�C�+��
V��\�q�}��!�۠ !�܀�5��"q .)!VQ�]b�R���ʿ����M���,�<��iApf-��t�@]o�4 �@^�@�M�R�畦����\;]�Rl #�	W��+}���v"��ಌelKs��)�\��3��8濡���'�Ӡ�>C��$�\�҃~��O'}�Ȯ�
�!�W��!0�T�q�{���כ�u��Mh�Yg�21<.������Ϻch�*u��M�{�6�K�
�%��("�u��z�F0�Vj��?�����ut��b��2K��;l�e	|�?��:�	�76ެm�jó8��#�ԟe|ؤ�x�� ����t}z���_�<�{\���ȝ�A��:w��$�Ѓ���Y`����SjVЕ��V�<�C�P��P���Y�1C��<�� y�� ��]K�!9{nbe��o5�ٴ�.�}�:�n/�-8k��lş�DnD�v�v d��bU2�[%�Yc*���n����s�����_u�s���#�';+ʪ���1E��N�@x�4��B���������D����#_7� �?�悀��-u�@�S9Jؾ9���?��;�>vΘ�ZXݽ(&�f�P��U��L@�X�M݉�@!>��,q	?� ���ᐣ��ﳮ=D0I������U��ԗ[�ױp���\R >+����y
/�o����Ɛ��}�~J�<����՝�'����Co��+��aɈ��l���<�$R�
�������>8V��^i���Ҧ厫+=�'~-ٯ�[���!�ȯ�-��k���dY�C��t����X-�_F�����B���V;噈o�_�?�.�Q�H:�������~�mH�i�g:�l� �G�1u�#����<~gW��%� �u�W����5?���(A�4�O�|՟�4q�Ui\��r�Y�pE V )�0Ŵ5ݿ���a��3���@�%ɼ����@$=�F�#�<�5ta~��d؍��:��f�]d��p��o�Z��Nlk��/����C,NA�͉W��Z��ԇ��w�b � *9�(} ��d�V�p��k���mj>�]<M���D��o��#
��Tc�N/D�J�$J�V�!+��O�t�m����	�D��T�UQ#��T�2��*I����A�q[�uw�e���k?�;�f�I�Mn�؀~�T��GO��@���6Q:ď�x���KG�ư�p��3��ſ:�u2�ou�zP�i�%�`,���{��2�l��3���r�I<�R�\f����C�r�1
 =�Bi0(p�b��i�*�RP�c�i��wb�$�*6z��s�ۭ�S��1�AQ?�fP�I�=述a�N�jNrN:j�f"٦�~J�S�a��"h�'"��9� �7bK��3V�u�¥Y�xʫ��j$G�M�q^/`,��-C㿹���tZ `q<=x	S����= �����7���k�)��c(ᰐ���\ߤƑmՑ��u�(���=�#�.K���=+"M�� �)�vź��V�$ \�V�g%�N�Uve�(L�.�B���%
�)��KX�MM�!����x�WI���bv�m-��'X[�S����( M�_��/��&yw=�T�����ofA����G'���[��:ڇ��6�k���_�{/3��lWU��+��N���>5�fi�]��;f�/�"�&���'���O�j>9;\��p����*�p� [���w���*gg�	jIW��$v
�˫(��T��%���8�LE��	x�MEu��p�A�*��1���PӰo�u�T�boP�r��|햢�X�5�AC�8�m�����>�-���A�DQD@��*���؜n��w��W�b�UC�-w��:�
�E1�V��>�Ƹ�b�F6C]�����R�u}�(=�Iw�TP	uTM%��y����8��m�b�?LL���|J�e��^��nc�?��ʼ輈ql6�:���`��w.wZZ�-km��(���O�u��*$�q�����bԗ��6}������3�S�4YH9�bN?��-9;G���Y_P4���9�~O�Z�L��8M�����R.C����4c���2p�In�b�����eD%����6x��K�O(�F^��＼�8�H�3�ߋ�7&���2�B�<��Tضġ�Mj�������"�����9��H�E-�C�� {�ѯ�HB.Hf�N�UG�eT�z�!�����=V���fW�Q ���`(7v�}E�^4��O���H��~~�D����q:} '���k�*
;�� :� ���7J�{��vxbL��}P��F&f}v�*Ⱦ_��t�@�<[k�*j%�lP8IhKN��Z8������G��Ҕg�.�?��=�6 �|W�E�n&�ΊL�۳�E���Ğ��w�i�'�a�|�.N$Mt k���GFR�����/e����.WI��Pأ��֖���圴�{�:�nc�>��S?{�LjTC���Q��U�)�`J�vYH�.�ܔ�:A5]t�n6�� �����z?G�f!ު[ݿ�z�C}ZAU��IM���~�Z�++�pw_�T`��NrR��r^>��WV�o���oZcI�Hm���yX��=��J6:e$�	v2��� 6g+�L��mҜwl�+-�G��pN*��yj�AbWNC���r����\�9��*xS(����?��f��ݜo`!;y��rb�Jxg�-��{�ȋ�C�p���{u=�`o�P��F�I�%��o�o7��l�qxt׽m@�Mj"�>a��ւ�t��5�4Y�P��Q�m��½a^D���Sc��x�{x^�3��jzZ[Wzj�z&S-��"�b����Xk��aJ]*��D�b4(��UB���A�^�tMK5װPѓ	/0D�"O�ëpD��d��4��� ,)�����%\2ye������E�$�/j�߷��N ЂiI��cL���C�DPB�C�l@�a�Yy���u���r���y�(л�+��N��L@�#��լE#�N�6 �E鑹�c�S���J��r�rӖzk�k��kD��{[��J�Pq/˰tN��R%�-⦽X��f2��� ��V��}�T0q� o"�W�-u����m�= ?[?C׳g"5/ǿ�i�K+偕hId�VB�旃H�m L�=:,92-{Bj�������.�K4OT��_�X�B�V�fY�w�c�p'j����o�l5�!��5�P������Y�o���t����B$i,q�(�au�����z��v,��M���}��:�C�]���F]7wĊ�G5Hc�r�>~,P��vX	�� 2�T	��Q��]�(�Q���"$,����� baVD�i���"��{n�KWσ&��L~ӱ�	�5��d��9�F�Zc���J����\pH�8k�C#��M� n�_/E�y�w�ǚf��!I�u�����2���؎^q�8�M�e�,(���ܪ�W	n�&�i���3!��j�C���kM �� ���%�1~u��;��IM�=��hj�����C�t�#�)�
�V�2�B*�����Q�`���Mce�w�}����\��*L��O}����'E$t�tI��&۵�/jE�-�D�Z\�M�"�^�0� �Y-W^=�_
���pg/*$�2�dkG6�.t��^l=�uRR��>���h�/���bOhKc�V$/��bE�6�~_zR���95����M$9Ѧj!�xn;0�ˢh��ςU��1�J�G����w1���g}�ӛ����������;VMlI~x���c�q����:�e��=0��s��/I͸
��?�١U��	\,��JkG!�a�����M�;P�;\a<�.�n�s2bDQ���(Nw�����E�;t�Rp�S]Ɏ���֊f�P���x�B�f$�	�[&���%�@�� �aB�~�L~Jr!���a': �kyX%O�ȎKx[,؄l�~����|����)K6� ԟ�K#A�n�|�^/�Ժ寑�d�^�nC�d*��eC�������Ej���#��tL��
s��}:��ݺ׃s��0$�/f�q�P��������V�[�cv�㆚�@T�Sy�J�\N�T�Xl�O��=e>9�Է!P�S��a �	Av�i`�Lӛ�E�����U����!�����p�aS<�ڔ`5ڱo���� �UxkT��Ls7yC�$*�>�����=�饀y�O��
�?�-̾1�����_R;�;}>������W�A+PH��=Oa�Q�����e&6	�y&�. ;�aaD`1$h"�j
Y�c -#C��W��B�� N4O�BL�;�َ���V�E4_�	A�E�MgaϑnC��BM���q|O���z�N%[l8Y���������{Ā-��[}�u�?L;r#�5I�Ӳ���	I�.ַ$����Z�-�۶�L!�`B�c\���ö��Dw���E�f�H(����v�e�w�}<��L����^����T��]Z#�k{�ס��RX&�rcÑ�hG�LV}�D��\�-�!v���[EWOh�B�C��A\&���ٶԷ>6Y��0w2�6�BՁZ��-�������g�2Mo���]n�|����n�Td�y+�D-f��<��)av�\?af�kb�m��c�k��Qs�6*�?x��5��&3���� )�+��S�FA�T�FE�3��4��I���l���Ӹ�|+������o�l����?{^d��2I�C:u�^7
U�����n�͒Yp՛�ma�����@�f)2S��.r|I��k���:0��A�(�r�Z N�gM�~��i�7g�)�n���V��i�Ra�� �a#"�o�KX
��<ax�7��,f�А�v�T��ͥ���ԇ+	�����n�����"6l �c&ʝ��o5֕�Z�X(��9���<��*��ٓ�+0��/���(�����T\�؟����&"������ �˂H/~2��е��Q���,*�ݺ�O=�����)"{���"��sm���� 7�_PPN50������L�Zt�Li�M���k�k����\g.���L�=Ϲ;1%�ȼ#���p�Uo�7X,��/1|��	�BN�]�é,!�*����X�mW?�jQ8#��Y�����{}nϞ�2�����}�-� f��$����#�L>��ٻ�X�����l�%v �x�PI봃�]`ʝ�"&M�[��^�h�9
g>d��x3m�IQ��&�L��^���0&}�?^�x�+B�E������qQMB�R�+�|A6Ș���X��h�.B���5�xĝ�����A�>gTEY��U�ncR7�}�=����~��h�E�n[3¾m<��:���jm�oD��W]�m��G�\�%������6Ń�O7�{-�����J��~�B�g�	�<�;G�����t��I>1�p�v�'<pm��V�ő.�߿/�8l�V}�m�pK��s뉴=V.3�����뮔"E���e��˚~��aA����r�dm�\q-��Y����V���lʷ�_�SAY�^�����HL���B��s�J-D��^���7�7"
=��)OI#�R#u��ی^+����RW�*��̄4%����e��z��F�Q�VAr�;Z$!�	�3��{.*0a_ �|�m��-q���0�E��Gw�|����թ� G�b��c��|��1yʓd`�� Ŗ�A$����(���<��$D3��';z��cWVV�U�4��.��y'����ɚ�]�F����o�åX�3�u#U�N�Ҝa��|�>i(�ͼ��^��w�S��70�js�O������½<��v��'�-a�]
PS�1�nd �)������$ �s"�2;�5�i���0�8��N���8�^�!9B�&o<��O%�x�t)�%c���9���D�52�Tb.���_�����o�G�@F�}��h,m������O�B�ŗ�j��=$�j��` +���2���k y��tj�ڇ�j����
R�ܷ���01��C���G=� Q��BS1U��YUdn�V���OC��T��4�K����o���uƄW��m#�uo���n��E
�I^�Ք��� ��V�����΀s�B|�4
�s��e�v�:%+q���(���[�9�|��:=��_Dq�����%�:J<1I����g�p3{�i��z	[e�m���SH=����4��i�{(��j���ExLr�8�:� X"�3��E iT��gq6$�ev�/C��O�uQS�p���=G�a4�p��Jh���p�:���Em�Ô�$���vH<u�=K�փNm���h�	45Q]��x+�f�vLy�d�Ǝ�h���AR��^f&S��\:b~nn8����x��W��b��h[����@���,��?G��yQ� ��u�	G%s��+��?:�8�;�	�b�^G5j�=x����َ�1�5j(V�'�t��(B��:|� �;�����h��?��ۣ�&�i[�>s11����ߴ�P&C{�ـ��'`����0���v�dm�|��k�ȁ�a�`n�WB�u�����!�5
U��K���n����{ك&��!��Y�����U=	9�d΃f��M||�B�*� ��i�� ��rي���A�P��#��)�,NM�{_nܑ�������
��W�h�%�RG�klE1��/�󾩽�x�l]ҳ�^[;V��|�k��N����>y�4m�$���c�ř� ��5�|��#��D�t���Q�4��i�8�[烰�$)�TMM�)"a��c�W�.4D>��2P�,��i���(J8����j �о��@���wW�``���=�y�-(LX���5��X�e�K]�)�lތ���kVG	�U\��^�z�r��7T~!�y�HcK\���Y�J�:�Ռֳ�1�kН��,���Q��}1�JO�l�@5�(�H��$�!�~��m�(w��O�\�X������6J �m��mI +xl�&�^/G���<Mh�L�d�X�@������Z�P�
{\!���å�0��Z�AH栋�F͌h�|VK��25K��v�y��E������i5.�-�y�b� �QX���Q��,�2�$$���vzqr��pB$�~�}t�2�AB�1~iX�o��s�\E1oJNhH���9 �@p���!F��ya'p�
Sk\ w�:9�]�ـ�3������n�p�/�� ��eZ�}C2A��k(ʁ�\~��ዑ��>|�����{�B�1J�P�3
QRyV|G�N�p���boT���4 n�_��ֲ�aV��,L���J57��1�~�]�wB�wTzzŽ��)g��tH��wY΂�j���*�|��"v���K���tP4߭�+ɖ'?��@@�D�  ��N#�Ǜ�M�`�j}���a�l�|� ��O��*�:�p�h7Ip���nx�}6X���ش���G�Di=a���5��uf�L�i�a'���&�i�B�9B����W6�k s3�I��e�(1����!B{M�Va���4t.]��=�R����')�/�U��(��b�Ѕ���Q�Shp���+,7!�t+,7KX�l4�"cq;�k��}E��f>���l�K��,e1x�Ui�°� Qt�����I�or�.�M��"�����G���]�F�{�D*��z�Q�#�ho[�g��-tW���U/�b�ԫ�'��>�;%9�����v8��%�$^b�B��aFwC]�_`��F��n��"w���7� ��q��6�7�� 	G��T|���Eg�U��^J@����)*��i^��e`W��`s]��Ǩ���L\-���M<� @?T%�u��(�:�	ɭM�(*��{�3pQF.[0p:֡�(5��Gk1���v��{)���>a�g���7_�6� �7�s���'�j��z�YŖX����7���'����#_No/�(�JQN�0ײ�܉r`#��@�&q")�S*fQTǾjnÖ�놋b;���:�.�pF�K��:<�Rk��O`#L���y�rԞ��rX��G!��4Ҧ��ĥl����a� ��;���)n� ���ƬE/΋ߪ�	�I7�@��hi��w>䞾.6' $d�j<�z�'pV;NP�!m�!{}Ӣa0<�_��B�PH��S��b��/���U+D`�3MD���Ii@���W���`��2׏�+<cC��m�ʱ��챀T���V����1�S��\�ge�#]��sـ�b���@��7�AE��UTH%{�:N�U�������`�Tf��	��:���-ex$������O����WL-�����=z���dk�$�=0}��k>°w�T]{5�	Zy��إo|-�?tN�=��&�on��W����,�9�[��	d��="�A��s˳J��E��Sc�R�(��\y�i[�;48��
uɄ��0��9C�r������5�z&��f�7Mo�[��J��#��&\�g{�9	�ƷTN��ۊiI~^�-��0���;>Y��Gؙ-IN��?�?����Wt:X�����V�F��+��`���!�^�A/&8b��۬��(y`�g��`�pnr� �!iw[�xep���H�iamXg�a�*+��P{����ΥOU2#p�A|`��a��`��p���W��E���v.T�:��ȋ�����x6��Q������bʉ $��p�#Y�t�B�QEbY:������̇YBT�?�rW)(~����Ǣ�4Lk��ʖh�A�o�!GjzS%TXw���� �ZW���ϙ��
�.�A�7��kL��B�� �6�R�d3}S��"�bu��X�
����R.��7�v`���R�KoΥ|�ߖcs�26�uJ�;�������6
0F��ϘP���U
&&��;"<u��Y��S.�p�S,ѭ�/�Do���� MX��b��Z� ��1u��h���D����b�Q�\W����>�P�8��7ж���Ga2�����
t<��^���~����0*�~g�{�~�ܯر��s�����&�Ƨ�Ӳ�N�ȁ]�"�[m���D+��A~VAh+���\��BYac���oN�.�V�>GJ+>��M���IzU��i��Jffˊƺ(��W��s�Q��<!O��#ZU{(�w��3�Ҿ��1� N�94$�b��3�ԏ�f?�"?n�[�ç}�%Z�) ��%TӒ� ir?M��x�v�F���9pE!���!'�ų�L,���b�~r��.u���9�h��K(�[��j��Nrܮ��C� �B��$)9-��`ՓE�-�{]YqjB�6Z��̚NEI��h��9�jxln��1f���γ�.�6��.����a��7����*]�����Sӑz<�������X:��әf���tEW^��MTݚ�����@�mJC8���R�`�63Zjnq_�!oU��\��*�:@�h���:.�i�f��>��p�9Ǿ��0i�ErgF�!���9bl*B�ݢ�K��7ˢ+��ꮙ�h��PU��Rq֖��ǈ7��#g�Zx���W.B���ݵ�C�+ц�s�	pG"�P_,��!����g���![��=H��"{s(�n(��OŃӉ���-_o�I����&F\�kL�X*����e?�4Z�<�Ӟ��ݗ��d�4�zoܖE�)�>s�o[R�n�YY��YGF����!2OȂЅ�6,\��S���e����o[���͋�H��
�`����]JbT�C�D$����n����Nf�V��~Kl�sa�0�>�V�d����j0u�6��$���>+`�ە	�ܪ�]��U���1満��sq�]-��胤JPHM�Ŀ���Fe��Ծ;&��/goo��O5�q( ^8����`��#�����c�+]�N��&���YE3�V(����5e�YO]<ŝ���XU��z���Ef[pK6����U呃b}8K_�+��g�=o⎋��	D���͵�O+�H]��^O�JAm��PaB��:mo�HT�� �����p{LૢO���h{���(���ȢLp��K����G:,R4� q�N��:�}!��(x��#�cV���'�<z�>�_�C�h��A+%��WCq����C�Z�|#��*(���M�7�b�I�>6�O!��������зN��L���K~��k�G�6��Hs;} �|0*�G(� jrp�>�N�8�����@sy��B?����@�\����뗏�E��S
^Q��˘˞�*�;�L�/A����=��Mu8�M��]��L�8M�����-Qu�/1��L-�$�x�2������X&�}�{j�j��2�~�e�qq<������dE�ny���`[�:`Q�i���J.��wи����a�RްM�l�B��J�����"�e�/�+�ꂶq�oM��Ȫ�计iz�IZIch�\�AGi1���s�$t���"Q�V�a�\��U�߼�]�%��19����ٹ����r:#��m��#��e��e����.d'ǽ&|�:j��a���|�(K1:ҷ�z��:�5y�_{�/:��o~�(���-��͟3��1#���A��\�Y���Ɖ�K�`Fb!�o�n-/S8i�f��T֯�F�D����P����N���҃�Y@#.���ē�Ogv��f�J����]u{\�}���Q����s���-���8�c��K7w1�����!Tn~w�e��V�Jb��� ۏH�NRx��ԟ�y�{��IG�7���}f}�R�=�aq-����>~��0�>X���x M��?@𤋮��Ƈ�1N���f����x����w�(e(�mI�
�fL�u�hѽD���c.��~�nna�wd��*���a=�v@���x�a�PM�n���{A�qn�����s�$w�BP�TX��|ƈ!ú7��\ő�uw+-6��$=�qx�~�H��'��!Q
�P�lǿ �E#������:��-��G����{j��SdK��w3����Y�k��s��Mu��L}�g��Z��G�H�9�=�(\[��T�������)��>I����0��̏����b1ϤWYy}�*. iؤ��1f$5o\	@�$�I����,��sn�����j�((�b�g�a�����9<P{�yw�m{O.���xF��Z�ocwD�\�⬶ix�f�������$/�����UV�V�3�g�2��V���q�O 'B┕���D"��hkLM$��P�p*��šl�V���ܠ����(�qU�����
_g�˒刳�_P\�ja�No4'�&}�>.�O�[��j��t׶���y�O�z���*Mș���	�q����N!�Ku׫�gOz�� 2g����|��L�βogQ:�w��:Y��ؽU����Y�*���|�A��M�CJ@ F�,CBC$=��P��&p��/Xy���ۓ	�>�j"@��@'�^�������
�SK���y�@�f��u�Z�+���T��u���0j���A1ڡ�.]�#��g�?e`�U(��\ۡb��U�� �cvv��_���ѳH`.��5��g� w�o*��@)b���0.`�U�k�5_�����닑�[V���&��٫� ۄ��m㫞t������&6���.г�
~�E���)Չ�9�G2KN�i��dY\sWL;@nw
���ߚ,袽1�H�+F�{�:��V�hEr�����I��z�H��vMN"�QcD��{�������?��,w�n�f����~��rA����"� Qɜ"�*�$W���0<�O	.Ǘ���s�_���Z��Z���(5O	���E�@��0i��62ʭ��͛u���A�w�,km�sZ��Z�ZkBsA����u]n\���m���� "�E���k���"V��Xk��W��zS�,Pnns��>9�Հ\2�>Y�u����/U�#p��]\��o��^+��	Ő+�[�Ӯ�&!߼ʨ]��>��Ж?2��2��:SKx1c�C�R�YC"���M�.�&��Ad�x֚�%4?=:��h�� � BL�e�6��	�_I�wk}Ө���m.�lr�7�y�V�<�@1dP]��N/k�;��N��3?�Ǿ��Yh�Q�A�J%������!Z�tփ�`Pһ�X��t��S��#�V'�v:�	nc�Ku����9@���6�GM��k�;� i(��(�(�Z�>c�r��nӸ���|��!Ƶ�����]<��)�E�?�a[ޯ�z���۰Jt*�Z^qt � ��zF�Kq,����1啉e�uEG���'�]�ad��@��#o$�֌A����毼���'�,�fG��/;�+����Z�F��%8�@�V���B�T�&,=\[ح��� ���R{�e�y��֌�s%��}�ǽ��ࠠ5�~8�ڇ�qyQ2o0h��g��9@��Q�D�c��7�	�I���!�ZV0���0�=D�զ�yQ!U�g���!ې�y$qޔ��>�ݦY���Sa��jD�
q�;ts�u���r��;�r��3�n�ЦNF7m2�5�+��������m�¾y��_���9<�DB6��|߇N��6���K�� ڭ'HxQ�Ϣ���I��|^�mHJ��e�h(���ZG�]ꃱ�w+y��-�)�4
��aU��\�\[k�͘�������(�!�?�^�й�k><X'���Y���䗯�)W������K�`�˲��	�D�ܛ�H4�k��s�~�^���P/�ψ����� iU��в;��rF��*�A��R0�UֵS�<>���3�d�gF�{�6���Rawu_P
���/0 MF�B}�	���e"\j5��8>�#���
�6 p ���&l=�K��<3]�.��AU���h��x�vǠz��*ȣ���cu��L���Q���U�~4!�Z������9��V��rNtn0NR��lA7�B}����_h �PLl���?}��ubN�����#�E>�%Z��Q5�S6s t��!�m`xd�Lگʙ�+�,u��C"O_������0��]�aԳ��9�s�䊱��ߞ�6^�^[c<H9$��2��;�9�299���R�D�j��;c������4��+M3ū����0������0`5�ޅ.Zߒk��'��F���:�`=B$�{Lz����}3B��cB�&���3.�`�-%�~�i�=@L�~`�ޝ�$�9�!�c�5�T[�b&��
�����F�G��Td'��*��|A`K�8�l6��w��I�ȉ�|�hG?׷e?( ����|���ӗ�/��ǮwwTj3R
�
_�Q��	�T��h|��L�4����Z�$�����g"�i�+Ħ+T	n�Biqܭ����=��Kv�fl\v�Q(u!W�գ��=�l���	��j�ױ�݀��� �g	�����maib�۠��W
W_%3Z�H��)y$?tن��'��#�-�>��R{:�X���I�7&kbΈ*v�E����+ʐc�쨰lr�]��5��۳֡��R�{��<ۃ���=z)�I�;�uM���q$Uע3ifz/�8R�6?�^�9���㇌*�s��C�l=K�1�qE��(��8���;�="#��~'!7�j9����1�!�s��a=)D�ߞV�w�Sōp^��_O�|7Uĵ=ۑ��:�}�G���=�Ȍ�f�R:��;;Y�ep?�9�Ǹo�,A���a_1o;Æ�`�[j�Sʌ3pJin��_a��rJ~���Esf�1(�;/��x�́!d�z�Z�da��mM�4��$��-hȼx��rE�y�}��>��m4�1�H�&�)b"	wR�Z�m��<�wp�	�V����eҵ��r�p���n�1/��[��Z���M������KB�0�;s����8���e�cW�����k�U�h7�b��y��pn��Aǎ!ް�H�8cx�Ӓ�w1&�Zh��|;�o 8�]��l�u�(�|%����z�I���Y���%�I �`���l9>~~q��D��E	*h,%�>Pp �6�wn5+	�Dǣ	N°eq'��[o�;f�B#�mcX� 2��ʗ��
�vR�]�fܯ_�@Fo�����H���w2?�?�9��'!<�c�ل�@� 1\V�c�7�ݹ�ɯ���eC%�ݥ|Ju4�������T��H�+���<��� �w�d"C$o������wO뻫����P�0Bd�R1l���a9'�C�'�$�ץ֦��c>kہg58�\Z$K�G��Ο=�PMř��T�!���O���}����#y>�pe��?6�Gj7P����3=��*~By�J�Smta�_}�d+$�bw��.�`1XOć��n}�����5\u^�
�&������H@��(���ʉ��cW�6�P�����{r���d�8KC�3��7+ ��KAaz��׊zs8�J��;L�_�BH�8|�x{>�\ϥ��0�bVO�����Ė��8���|�/H�u�|h���P��xp�$&����\�����|l��jV��u�B�tj.���F�ھ�ʪzo����X|�p��S.E#࿧�� �`�?Iα�� o1�Vi6���ގ��,���P��E#T����m%�.�<�v�XoA�$>$Hcg{�ࢷ��SGu2?���;
-|�sJ��W@B�Ľ�|GEpbU��=;��i�A�8x4��LH�K���4y�#����xeV��b:_�B�s$s��6��R�W�-暖ʜZp���{����O�k�V@��9��8�[��[/w0�9�55�黢d�����g\��4���D�ƹ��qqYu��(?x�3GBA��kb�I�e�_>092��L. �?����y�V-��.�����^�^���&)��]^15<-B{_��D�����.`���dݛ^�����[+�K>	D7M��H8���G�������0δ���٨u�yߨ��*�r�]�mF��a�<=��k�U&��ϙ6y��B�]8��Z�iJ$��Ꭓ�v�Jz�p�X�y�F�,�^�.c�[�DKJ-�hwۛ,�S��زMl-v���T��j����'X��'��c����F�{��	�2�q�Z,?v�Χ9HZE�������o��Q��(���Dpy��1#�#��2���4y�)F1��r��Yo���ᒉ�5|�ɞbn��eW��1VV� ">व�B����{��|�9@��X�WzJ{��襲!���a�6el�gE\�\`�8ɷK�ꔋ͉�$/�{Jƞ�*Ά�p1<e�92�x�����lb,T�R��J�'z4�]���e�#��>��,d�q����Z2��!�z��*;j�}�{/��9�J�X��U��'�=,H-��r3�У[��T5�Ȍ�QJ�<�5	��K�sї��Ɗ�������`y���Y҄4D(7}*f:u� �*'�L�l�4h�^ �Hnylv�����`sR�Qÿf��'����p������m��X$��Mu�a[!ۆ�������7��*����xl�6`�tS�\R��B����GΣ26�֕X67�Yj^qqU�Xمy�3`�@,��O����Z��"����f�>Ù�����ͻ���p�>��|�w<%�$8p�ek��ҿ�|H7!k���c�Z����7�^N+�d��z���ǲS0HHۓ��+��[��Wޔf��@+����E����ٞIK	p۹��U|��0�=a�ׯ㬘�[<�H[���K���-�9T����2��w.AB�~��b�h���̂����%�.�R���U��j�.��j�S�hy<{��B�խ�ʹo�a{~�]D���-�� {��"m��*���r�Ф�������z�(�爎��ON{�zfVHp�;R�8�!i[@���$�tf�B�E�1(w1,��mʽu���$>�ԃds4I]O�_�\�r�^m����8L�D��1KR�]��׵oqc$j���fX<AԌ�*�U���tm�H3��������=��	�+���+@N� ��Mg��'�k��H�dڹ����ߧ�񜰊ib��E?S��T�3|U�ĴDR�9���C]�ghK���I0F��>�N�G��c	\D,�2I.���Q�RԊ��HC'_����q�ؾm�5�����nHck�½ԌT�{[���E �� �K���4|�Z��sIM.fۖ�.��ܤ�rRvWd��e��j�
���]� ������̨���������_xM��<�
����j�
y���@���QB�����ŋ4�1"?�=a����ω��5�M���b��%0�p'����'�2o@�{�ƛ�H�]�w�7M�K@v$4YfY�ղjx�W�	k���ʲ@GP�l��2�5��־D�;���N�-M�O���*���@����|�M�n��T��h�Un:�\ǖ�K��&�#1~�@j��y�������7��%Z`^���9�:�]�3;3���4�6]>�l� �L�~����,�X�}<~�c�̬/r�����0��4����P���}q�~O�ŞC���v���������B�2��-�����3T���w�ѿD����K�T/-Ͻ��3c�E��W�/!?��4�$|[[	�T���3�� Z�3y����h@��TM�`��GT��I��6_>�W���-6sV�ł��ч�R.0�<"�qv�ep�v6B@�,	�D:����s��>�mkBί�,v�U�ސ�t;=~},�Q��pG�+=������$lt�b��#.5X��Ӭ>��Z�&��a�|rN�&u�nM�c?���W�����\P�c�gi0�
ԙ$;��G��v7K�ՃE�������2A&�� 5��񓩤�u��}T����.��y��{	=y{�ᦽG�9�fk�@)��*����&2��H�'C�
r�*֓%54D��LI�Rhi�ԩ��0	�v�1��X~V:ZЃFK��Ϯ��>��g$���G��F4���[X�f���;��P&�C$��B�X=�����FT�bKL�,hXo;
h=WgT��c��CM�wu��˙�E<�WCt�g�Yu�]��j�E�5��b+�!l�^W^�	�I�Ѱyem ���+�8
~gȱ6�V�`k+����{B[S?���҈���� d�#M|���U`��S�����G�."9L�(�4">��Հ����������D����4g�V��7!sn悦V�ٙ�f����Q��?�d���z�r	lz47�<^�OŨ>����YB�|�K��t�,���3��jPz����[<H�GHm{>�PL��kLbƹ�8P�[�Ȝ���n֍��&�QD/�Ű���Z�d*���j�!�<C��BY�M|~����bB���B0������t���I�/����9	�=��d���C�(Mʍ��K������q6�~1E�$aU���mh�75� "�8���:X����o�B�U��۪�V!(q@B�wT�(�#T��i���SA˗P9Z�L�NRWm��bvT?����͈��r���]��6` �>�_�|��x7I� @�5f3'I����I����L���A�ſ��Yg��x0�(��*	;��M�L;�����t
e$HI�jV���c�R�]�F̹8��D�1�>Gq6��O�FU��6�`̴}w*X���{�<���OkFw&[W���A����Z��w�1d���Q�W�d^}O;��9KZ���Z�$ M3?���"﹔p(��;������o��NF��#�;���
Y�
����"�i�?� ��8O8�7,R�r�	�o^\��W��@Zy`�����j��@)�3��ƥ�<z'P��6�s	3�w�������d��쁜�v����jU�V�]k4K�ܣg��*z�3 �NR|��Ƕ1EQn��q�t-Y�|<#p��[�����2g�6�/�-m�[I�~r�t���A�D���4��$&�H�2��D�E yS4V2� ��"���Ԟ��X?txxp����G�g�0�G�a��;��� �iP�������%���}�
��縜͔����]�E<m��GJՂEI ߰Us�/�T:�醧r-���Q�k�u�-�����gL���G!��\��+Z "�ţII+&�u����5�M���طe-@Gﲠ�4(�i�S� \�n����ώ2�f��b"���]�2T���/���:�I��`�pR���s�k���H�եv��9���hg��]�~Nh�� ��g����>�e�E�@���6~��w��{AeU�1)�D ��ёr�Go�0�5Ă�*4�����ІB͠Y� rT�Zr�Zmx�A �$�ߊ3�,�d#�F�,^�b�td{ɖ�	sj]�6�t�>��nT�G7@���.�>K=}��!� �0��|�:�ИV�#J�>TE��9\&?��$/<�Gʁ�IC8�.��LgV�W>��~���Oq�3LC�5Av��&#͚�������yX �_.�"`���ʴ���=�֩>
O��?���%��(��ju���ì���݄��F����&���b�s�AR�_�����(M����QU鋛�&"G����ޘo�?�r�7m�Q~'��s��Vz���m�5.�!���Ϻmz��#Aa��Ԑ��R�{]!5�q���E�� ��" Ӓ�3�"+�q��T���?=d;��M�g4����������I� ��n�XN���?� ]Q��SRܨ�j��=AfcG�8�3�x�.�x]|0�,-�K��5�#O���<(u�l}`*>�7`�[������^�z-Y��-�2��W0�'A�th	J9��p/0�ڠG,��M��4�i��� ��REG ߊ`U\���ɶ�H$�;Z�E��H
:?�YW�3o�-&:��Yv����o�4����g�)�pk)��Ae��b�rJtA�6j+��]�Y�A�7Z�FHӭ�}{����֚��>�?�%�p6��TV`_U��9a��-f�zb�N�c�FC�r��6r��<�AY�{�1��p���j�w���Ǐ��<iS���A/�0{��ޫ5�D~#��)ۃ��_��?��w�/�m`g���)�bk���,��KTP�D>ŀz��C[X�i"�v�:���\�.����]����m^�Ҁ��h%z�q �5����X�-�������"��3�&�`��{M���ՊtH6<#M���-�[� :�"��(' �5$��B�I��>;�T�-�[q�UЛ�%&P���S���S^Գo��i�H���`.�aM�8�өVw��?D��Ae��'��1t^�f��$����,^��X��(2]�"�J�2�쏕�Kv��v��T'_g�� y��XP��J3�q�(���q��C�)El]�`�)��:���)�X���G�(}mA�N�5
t�*fgLޤ-��O�C3���©0�g�j4�hJ��}C���4/�5�e
�'�9'�X�E���&C��ْ[/M�"B	��<� '�Bc� ���S�}�Ow��?�����U�ʬU�2ǌ�D�
�����DE�-�_Ŵ]���ke&[J��^(����ɈNʚuκ��MX�ڗk�[��
����h�qu��ē� �:�b���Kl�ÿt�61���H���x1xY�D��	�NV@��1x�Q�On��A$*Ef�؀vZX�ʘ������`�r�\�(�u�?��Z���F�Ku&�AF�%���9w���7�L�:��kM��ʹ54��+���E��K���=�X4�����v!8��r{q�C�h��,��0M�<�@Ũ��X�<����ge?�jYiu9��l/w�����=� Ӷ{�*(k�V{�g�!�����.�s�1�%$d�|J<�1�7��IཀྵW	���<����:� �o�DX0��ũ� �ҡT~��5�����R<����(��z��Feno>�҂�������u���Q������2>L�o}�Gqm���]�ʃ-7+�L�a��8����қ�`�+z���x��ź+��#��x#r
��nD ���߂�k�-|�r�wi�G���LH�d�}ٺd�O�w�+��[Iy����{p�S���C�����q}.n��`a]X�h��~�ϵ���&c;������I�� ��nds��_��c����Z�g߆u��r�=�:4V�Ƽ�n�.<
-�8f��m�\�d�e�ssT��T���p�����2V,S�Vw� ����d�l��y���3Ų�p�G�7d�yw�ffq;X��d��	1��c�|�zyʲYx`�M���×���z'֍���;����W�N�s6�6��E`5�G�%�,�i�t��"���3ۿ��׹�Kv�j��-�ƻb\���_Ӽ4m���$ca���K���d�H�w&/�}+=A(�*d4!�䀢�M���t�ɘ��$�F��)`�H���ݒ V�	�xC��'�� ���ʋ�3|�bN��,j�a<"���uƳ��W~�h�̀�Elw�+�����'��|�f��'���Ϗ-�� <�d���b0a�L�i�C�H�i�ق	��
�ǜW/i`��"��q��_;�jc1c�h�ʻB��C3.{a�I�Rl%6��m4�t��~�XX\�l����8�m��$��%��̩�.���۴�����A��b=�̧u�d��m�"���G,�ps��LQ�"����X�ZX׊��#h�h3�G�tv��!��J�n�oG�A=h�"�JX�vd���NsH��uv�"f�{Kp�Ӻ���IL��~�BX�]2��l�k��q	���Mǝs$VcѤ3c_0<��b�c��]�&��p:g��J�W,W����{�ϩ�}���g��'(��������A�ە�;[���b,t��H�$�/��\Ghu��6l�O&�Q1�j�,��شL�$X 
	9�E���Q,@���|����0.a�f^7z)&��l��	n	K�}�1g�Q˒�p{�y@q����@�*A�N��8θ��(v��c�j�V�Y��"W��N� ��Iۻ��C�5�1CGzg�]�����PpHS
f��K9=^�+�#
�4�6tx���H��f���G=E��F�Z�2��};��
J���<���QlӞ2��WT_@��_�r�w`c���ơ��d�uQ�$,/����V`_j����!!4�*l��$a{h��,6�n��Zf0.��!�d>�?���=h�8d�LC��_Ul�� �=?}�j`�e��1��sE�4ρh���+���#�a"�EՀa�xgM�c�����3�Gӫx3���UMFK}�uCe?����q&�X��:�o H~�m�w0�'y~uO���DΠP���&Ż[��)����fhVfM��L�N�@8�J��V����mD`+ّ�+��}�J4���oY!�����,
�䯭b�(�CD��O�N�"~�o���(�qQ�>���V�@����#nhOO��6�w;�IdT`�$8�[�'��0'����O�<ڎ�<�Z=�"��7��y��s}�O�xw@a�*7����W����]�y�'+ig	ׁ��!srz�c��)7G�]v6�èG`���)H�q�#�o�&��7~ړ�QT[��Y/�F�����@�bҦl<�B�:�,浏��Uͩfj���ƎP��,h=(�`v6:��@���J�� q��_�@��ҶZ����ƅt���$���B�Q�5��	�% ���w?�%Fo�{�e��AS���&KreXU
ԻDG�����?VGYR~���T���?�B��L^����
"�KR٠F��9í43�L��t�;y5�$�;"��)2���^�ǵ+Ϩ.q�ۍ��(��Ȍ�k�'0:����Zk
ͦiSPG��%X�6S++�/�w��JЭk�l|}.��-�oy�C�ɯ��#HqL%�\4�^��c �&�J��Z?��I�6�y7���KJ�Ǚ��(I�B� i6����4K5dQ��q�p}�>�l��Rt��z�,���FYe�������5��#���mIR���J�|�5���c�A�c&]�Db�F|��S	� ��S�׊g09�'�V�#%=�����j9�  +�kx����,��ݮ�rע'h��L�؁�$ ���V����A}&�vn�Ѯ��UU�DQ����!�M坫č`�|d�LTsK�Jl�{�s��!=����咍�+z��M7}],�B����5ф�@|��+Ķ��~N�^��a1�+�Aj�M�3>cx���ܖ�f��K�5O/㮖��E�(S#���'�A��j����I]�V�\t��M=ɮ�n���a���m�{/�~���e�Ǽ]y`���iba��R>~�Դ?Y5�̇�=N�F�6���k���*�H�K���s��^�7l�He��>����!�� 
n�_�>tJM�E����{:�'Rͦv:r$�L�ׄ��=g�a���zX[�kS�ye�GQ���(3�^�y�����Pg31\���r��-��X��0{�Q͵�W�{�����ŌJ٤Q�wX[;��gC�oD#ϕ��	?����x� �e��5�/����e%�c�K�m�T�`����.jZ������PܼG����0��8wj�V;`p��	�n��0D�&nʋ_��S��Hr7�̫@�f.�}�E���E�6C���6�q�Oѯ��}CEG�^��`3�����C��V�w8PN]'��\cĴj�[@f����cB� ���$���T@K�)�0�b��+�a�����C��Q��8Dz�$f����hj�#�n	�B~�~C*7NM�^Q��z���Y�g��ƃu��\�&8�LZ�R0��l�cm�-@>x��!7Ҹ�����qu�]��J�'B���
�b̄p��)�{�z5(z��A,���.kX&1�1�������}g���|�f�TSP�)S��W��Ǘ)egU�D5D�F�&39:��9�Ӏލ]��v9���>XJ��;��wS̾O&m���{3o��ր)zmԠ%�?��oݚی�#���yI.,�q�u�a��	�P����6�g�>�\�;YV�|��s�(,��z�We9\�7{��%��[S�>��m����}λ�Mې���p3;]�pM�K$M���^�Ё�Vf�o5�~|f�<vx@��!���o��U����76���&d��N�������y�.����~P�G�k�O�0�Ƃ
��yW�Z��{'7n�Ȗ�2?�X����/�.s����r$Ј�"R2�u޺mA���/��?o�mF�?�1y��I]�Ac��b�0��h��rji��v��\��-!��7diofQ�BuU���.�vA+r���J���,V6���2���v%��ƛ���(��=`���~�}W�v�A�[C�V94k�5#a?zH�^y��
�3�������&�5����gÿ\�G/�+Rb���*~&亂�L$;`��S��׻�8`�-��pl!�_^�!��Oǃ�7�8#J�
}uRf�7�	=f�MV9���)"bg�ȋ��<(	��J�ٍ��$Z�-���Lb����f4 ہW����ns29��#���B6�I�Yz݋�H�=�au&�g\u�oz����hhR-v�j|+�]��G�p3��i��N������4��@��s�8A�<��w��`�Lb3�g��\l���%94B䰴��bGC��Y�_��Đ��>4����sYTC���ev��D�whX%i?i"�8VF��0spu��d�s�s;nSI���cIGT�ļ�}�Qf�J�����{ɥ&�P�%�r�b�X�7��ˤ��M�/9���UA{���E�/�ɰr����=�-1�q��m1.�)��.,Fʆ�6Ʉ�,f�\�a �a�J`E���=��iFiԇ��J=�`�Ff�MА-=�ḆaU;Om�!�o�p��xl0rZ�����k�h)n��hN8rx�Mv���[p��{���~^(�|,[3{M'e'W�
�P��aӬŭ�2{��Ұ�K�i!�˫��wG�x�k��,G�H�Z���8��D(�ܵ�>��&�,���������zd��(c�����݉x�l ����K�}������l��!��0 ���qU��q0>g��O��^��r�VW���zr.BK=���3�I:���Pk�(�.��ƻ�i2j��4����{��"`g��z�ųx��!x}:`U/��`[�B�0.���ޥ��б��P�Gy�U��?���QI���=�
z�{|�Q�Md2��IoU֑?'���jS�;�&���<٫�W��Û�ӦD���R_/��n��A8�6�}$�N����܀������}���m�J����N㚓&��.��
Qv���<��Z��kd{��=���M���Ѐר�<U���D�NH?�^J66�����v�&ȳ,ږCZ���Ԥ2H�\��4�7.��P��Z+d��HsW�x�u�4R��b�A; �*�=�*�X�����Jq�՗;	��vP�����n�I���=j��e�hu��=���(�G��:�^����U��ȿ��!�Y��4�"���Ս�E��"��E�pI�w���m�C�fE=$��k���7(����F�`3g�J��oT?873 8:��E�ϽE֘���朽r	-�ijO����[	�,��U�F+0��f7u���f��I�A�g����2��dm|O��w�v/cx݉"x�&���I~V�t�r��ӭ��l|�U�/�YT�d�Gr6�AZ�.]��3�D.0�nK�Ǳ�)"`�n��T� zw��1[�"�xJ��S�2�3&ѐ;�oWh]1�I1K�z��]#u7ͺpy��sb�8��0
�\���xe�Nz���Dk�İ�{D��LO�XW&9�?[|�b&n�����Q��P���+$�/Ze���LƤ��\cfv�z3����>2�ў5�ƒU�YC��o��҄�xR�fs��>�x�p2q��%#�m_;֔��8wt`-�TT�]��h�HYg���]��-T>�X�ݗ�H�V֮�'-.^w+�r����p����K�Dg�x���J�1(Q�vO1��}�U����T��3fz��3dv����av-� �tK5A��d]�+b�'�����/t���à��H�H�8�JU��K�)�)=�R�i��r��	]�{ͪM=�b���lWT�ww4&�2��J܋�T�վK	��P��dG�k��� 9UɌ�G߸��w����V\�ޥ�q/�ǰ�΅{)}�@Nۈ#�Z�z����.�����|#��n�t���K�$�`lx�BjO���	����q��IA6���W�ҍ��H���[K��E7����'ݛ+Dvr �u0I�p}��茵�
�I��NqV��FO�QP�,&<Ƹ����9:�B@����{%vI jB�m���ο���f�dͪ�vq0Sr��W�S;�{�4�u���|��cjޭ��}�����P��ܛ,9#$�VB����e�c���h�i�	�Ú_R[����q\=̭;1ň�R�@(
$��{���.>��Qb���Į@�n��6@y_Z�Gΐ��� �*�]���"A�>�u���}/>�S��Ɓ,�5!XT��*�0�E�2	�W%jL�1gT+������v�h��j�Q��4�7��dڤ�?�ң�g1V����� ƛ��tUn�B���mq�Ɯ�闢�,�ð�ÜE��)��Z�>���P���J6�w�ҟ$�FQ����#�.RͲ���x���*>��D���|MO��*�aeX} �RN �r�QuV��� ����*�y����@:20����.&�SWSP1��k�n_�!y�ud��1�	5�r����p\SY7���l:�Q����9;�Dȟ�策xTQ�3�/�p���a砄��	����'Zk}Gđ�&Y�	Y�W!g��
	���n2�B2�]?��y�ȍ�i��˚J=�|؄�	�+3r(=��~`o}C���%	�3;{�χ���eފ��<Myk#�XR�|�Ԧ�w����� Qd����[��%��ͫ���Cw�I��!��� :��>e�Ī���������� ���FB������(]�j�ictۥ�	F��ob�=�5�[xOł�'�	�'.A��t�n�f$8��8D��dz�U��<vN{L`,H� *-"k	��"��ȁi���̡!3����'�����P��W2��g�:����'j!�\������S��:!��݆,1�gĄ���W�(�غ�ۅ��[�.	�硫I!�����7-&���K�x;	}��&��F��3?�Qz��S��j�Wu���$�Žk=���9Rm���Xރq�uA5�h������bPx��,{��4��B������V���R�r��Un��oH��5U��o6�1�tSW)-G�,� ���&�XX8��V�_����Y���zQ����풥T�Г�@e#n�`Ә}��[A�����,H���h�Mm~��!K��$�����w��8����hgjBYS���*2f����8�0�KA޲�0vת.���|�VO�$��Eԕ��bx׆��Q�m�e�7��:�<yٌ��+ ���|��"F���_X=��wY��|��pD4��ɽ��u��e�v�����uB����Dr�����OQ`�Z��M�R#��2k8eƧ�a�UtY���
h�Y�%Ʀ��`uf"g�����/hS���G}?,�J>�i�����Vߚ*-ִ���� Ҟm��f���>ƒ�h�rw/�Yj��\KvxeaoA����S��p.kH��ڋ2v��q�f��(<��w!��sT�������Ȭ���&ǳ�,�gۥ����F�����&��L^�(��S�bo�G���8��7��3���I��G�NS�L�)�J�Ϧ����&���l)�$�����/�W�.]Ϩ�;�c}�$q{������7��65i�Y�[���Kd�/�+C���H- :ԁ;�lz\}��o�oG�L��a���O�*�`���(�I��|��c�o��W�����k[�]Y���"�����N�����1�����т-=�=.4Ovg6�(Ek�T��~��L��j���7����e���Nf�<��C0<�d7ht�H"c������m���v�*G T���{�M���8 ���:嘛���c��R��(�'���:�V��]�4`M�-jU%��pi��x�<#��9�R5/ U�`X���Ns�Iͅ�#$��Z$���[l;~� � '���1T�v��ǸѶ���[��ݤ�g��F���yÛZ��� �2���N�Fc��RAs�Y��D�.k�ԛ�\�:��X�M\l����/� zLT�]���:��Ia���i+e���р�M4G�|�H+!�Ɩ��K,I߻�_��r�5���:-3�G�کh�p��ߪt����g�wV�;O��_H|�}^m'I9�4�����Ȋ7�^�B=��2�J��~k�l"��WZ@�S��9�ʫ7�~8˭��cAs>V���sf�L�5���y��J3?�X�x�Q>������w5�*܀i����
���M���^�s(�_��/��9Z�J%ê��HR��+	P��Y��M�I*d�͓�.�7��w磡+$��xj�.�#�rO��f�^����
B��6w���u�|��~>	�[��}��i�J�y���D 6�@,�BHU�k��%eh��}���C�^��9�_yw/B>����|�(m7rj���oElɇ�$�����!��U���&��Dľ��IΚ��kAj@���ΐ���ΰ��|�<9z\��Խ!~wnCc�0kz��a�g�$*�c�v�n�Ɖ��'kq�i��T%��Z=�E&'�0����Wf.x�hQq�3�qoo9�ċ��h�{s�8+��P�+�G\�+r!��,�OPMs��\�+�H�Nj�=ѥg$-6Hȏh�G�/r�K:��)�	!�1��,^L�S's�j����A�+~�QY���,h���)�l�0�,���Nmߍg�h��B���Z�:ƍ¬��6�ѮY�D�1,nL��1��x�s۲;���Bɳ_�dW��|2��3TÉ�~�Q�v�o%ېmc+�P�IE5��6��%�k��LSdSEbh��Z)mѼn%�P��Xyb�U��$���&M���@'����K�AL��1T�:w�W����%�4c\�q���M��W̝��F�hVS�ƛM�R�����\���K�bv9�N���/9�V����ʅ�`F�7�<>K�Q���?-���e����e��eX�ElɃKi�� Zĥ���g�@%`����gl>�;��Y:$����_��Mȱ�D3��dZ
������<2�<�B�~���E�V��Z������8��zt�B1XL+��H�ch݃�b1����x�X�/�$+���X��yoB�W�{_(�Ba6� �0�b���D
�(N�s�}�4�P��. JJ��ּV�c���!����[�@	vD�T)G�8�
�b��'N����C�����b��h��]lvDA��׈����! �U��𠅧���B[k�p5N=a��hA�� @����Y9�ROwE�wp��h�Q-�Y�Z��t�V���6��Lz�D��e�����`�%��գ땻��ps����s�f�:k{�7�_^�p�����/�NI� $�zY�/qڕ�ڣ �S���_v+V,$+��-���__Φ�MZ�Q%/���D��*�U��
�W�*��S�ȸ���0Ϭx�@�,<�pz��?Z��%g�I@o��pQ��s��[	,�$�W���N��ᴜw�,��%�n4�~c�����Z�\}����c��ҿ��t���raYL7Ej펅y�'-2D��b��F��j)�W���SE�A�ȶ.�L�@�L����L~���X5�>�t���%qh�>Mmg�]@+��|�G|@7)�θ��K��i���FW���	|�}�l�+W��_%f���#Mј���&���{�w�z��g:��W���SHi�xr�{{r#� ���Ѭ��<�1�,��+ ���t�7��=���R�TXb������c�e^���f7��ɲR��n�z�A���J�8��0��	���v�Y PeF��	���B�}��wx����p��ߑN�F��*$F%�c�@��>���|g��'VTrIe�̢ן��-
A�7c��L�X!��<�	�n�0���Q��QQ8��/�ņK���ݼ�ܰ�넩y���LJ��)� �Ţ��7����r;Wf�i�� s��*�X��j���?ܫ�Q`v�]x�,�9g������O��Sg'�q/�g���ȼU��9"�p�׸���U2��<�������O�ep5�7���WX� ������M.6�
�i�(-�ks b����p?vt��pR�����&=+�$���9�!j�w�KY�mY��5l�&PQCZ"5�gM���
�����
=�M�I�/tt����l.�Q�Ϯ�C�l`[�D��٧�ŕTI�e��Oj�,����r�A/Qd�R��Ol��\3<6y)*���،��[Ï.M���)H4 ��Zo-����r	u��B�%@�
��HE��K53���Ǣ:9�1MQ�!I_��1�?+���Sۂ��G>��h��_ˇ}F�"[_]�=�7*(�!�7_dR��m��S�����ۧ/V���b�R�ɪG�EV�ɾ:�SrNڟ�.JTT��-�j5�L�Pp��Y�h\_�'�Tn�^��?ʐd�vX }R�m�2�����`¹��vEH|޸l�r�0��3��R���Yz5v<��ŵ�
�%�?�n��`_�xŴ�;z�R�_����~Mwd��Õd��Db"a7e��=6@P�aS�aa=/Z��ʃ��i�wª�#��k>��oY]=��/;�y��z�Y�)s�Q�2�9�3@��W�����	�,U�n��=�I���W^@82Z��T��?�-��U��L�V���f��]_%�z�ʎ��\xYZ�4�݅Y�&��['N�E"�9�v��� !�a���Fx+�e�.%��)����I�"�;�:�����v�8��M���S�s��q�R!�-:h)_7J#��ʊ�`�[-(�a���L�
��GW�GKg7��~����6�\u)�(}���@���VC(h���I���B�9	�U�܃���v�|]�{�̡�NR����V�3�J���R# ����5M�|S��KG�e�Y-��NgA�������*�P���:yٖ[{�q� p��c��+����F�]�7��:�X�����<���4#��-x�tb�O�f�Ӗj�x�MQ���L�!׉c5� �?�"h��3�l��jc!��{�:H.�.�X��D��k�=s'���C)	D�����8̥S��$Q1 |��6C�i=+���$�N�l�mҦ��}�"�.p>��|*�;��T�[V<8=��b$���ʞ+UO9���v�閹�ؼ�Vk6���N ��M+<J�w�	W���#��*x���A���J�_��b��� ���ݮH����v筵�����R\_^&����J.AyM�᤮�ٚ��?�h�#�#��r�aG#�ȍ�߂�$��ޘ��ύ�~A�Ye�ޜ�O̯�ā�̀�-�1w��N���brD�D�O{;�+$�j$�8��'GSܰu| aB24�z"&��h=��ҁq�EW��}�xU�tq��(�:�-�G��,i�q���PJGӕw�*И���VR�_7kV���z��E@�ذy�t���}Cg��auQt����s�P]$�5���[��W�φEQ��U䛻����C �$������,���%X��Te����o�Q��λT���ҁf!�[i��g���e��4�M�K�oִ!�l�%2w`�R��6#dV��'�*u��^(�I�P���J,����L��O?�r����A���Kl�m���ɷ")r}�|uI���iD"c�;�g�r�@`@�p�9�Ŕ]׭*>YR�sȑ�^��Zxq���2�,Z��EK� �/�F������n�,��g7@��G���NQ/<��R�NW�d������x�4q�����M��V��xܶ�w���r��r���k~+�F	�T(lG�t��Ҹ�>K>{F�:vNs8��](���gX�'Z�p2�a;C��ޝ�`&�U�����,�	A�2�	��RK�!��i,d|�{ӷ�qR(+(�њa�F�WB�ݶ( �|�*:�ȫ:j��u����68,a�fZq�b&� k�����^C-��}dz1-�k>�q�z����@�BMp�J�e8�*�KV����QF�Qk6��s���f�'�l�cĊ�a��5�]	�x��|�q��|B\���{�d;�M�hVR�;�N�|C��q]�+�S��0UF����I�R�u����?������.��E�ĺ;�ǟ����/�t_d?��*�D��f�J�5�]\,!����$e������u��n�R������U�M�؇9z��
w�d�����#�g���;��Ɣ��y`��	b���>M�f��2�;C:$�b��x(׆3�h��S���Fy9�[8����NA��z[�b�%��7{j	�ժ�b���(�m���z L�m�1�W]IK�
�x�p�hN��K��~T9�!_	���[������vb ��*Κ}���]��A7Ȗ�D�o��	U��/� ��-�<S�b}z�"�����A����E��<���d����
�黙'��v��J�0�u�;l����b
�E�+��pޅ�Lmj4��XE�j�H���  ;�;�⡨����qˀm��z��)%���x�4���)�+�Z�]�{$Y5���.
}k䏑N�>s��p�/ە�[��4��wPs������hA":��w/�/Xr'�v�b��rTm�1Eiy2|N�M�B����tz���[P����J� c�$���S��#����gs�����ok����-
rK'ʒ���� !_ϔDw\�DLI:5��fCa��wJ�V�.�-�f
O��f�Y"i����n�ڤ�{�{GZ�
�$B���<c�����躼^�C�|�y�Kk�gc�u�u�X�x��<�T3�c�.B�����?�؆C��4(I� �*跧Lc"����č�c��xW\����Xw��ؔW >�#|��zW��lή�wX�^�:}�,SJ�"��� �łLR�cc;c�9����:'�7g�]OZ��a1��@�&DČ�Pa�^��`"V�~O�x����t/��_ 5�n�o�[c�ZC��!{�#M�w_���V=駇F�:g������x��L�K,���a��T�J= c
t���Z��d𢹰9�2I�yc�\,�z�A������ ��+�J.�"���qw���%��{|�k�R����bI9D{�!�_�f�m�����?aW�3z�'<,��l�m�����^�.�7]� D����
�uS�����&���J,����n����ur��K��x�٥+�*;��î�w*ќf"�7�޼���IЩ�Yh��( ?QiĞ]\<��Ɔ��${c�
�*�\	 ���L���9��M �Ax]eV5������O��w'=H�'�0_	ieBv	-, ���p��j��il¡�/�;��X���I��n��QcRI�ȢfLZ��b��c�-'�3-�B�x��d�>F�x�*=��儔w����7�ō��(��}�b�-x�(씸�l�Vpg�В9(E;y�z��M_	c`��Z*��:�:�O�]�Fт["��bXQ*�Ȁx
>ޟ�ϧ����$��>���顯��!����&��W(8�g��ĵ��k������r��S�Y���5�/�F\�J����}QL��J�"5)�_!܉�p��q�����de�{�H��=J��8��@��0V��U&@9��j�~lo��-�9��K���n�r1"�0��9�^�3��ũ5���_�sc�7,;�wʵ{\~o=n$%ۢ�k!��:�l�����?<���F���u�pɄ�)ᮬe���)�a?�R'R�R���J��ܤ����kF���ЅP�\�Gӵ�U�>Rޗ]M<S� �bW�~�w(�	B@Q��M� ��U�|������j���V�|܇:���co ѯ��_b����*��N��V�㚚8k���+��7��$-d�2=Ц�m�2A܍c�N�v@6�<FϭW�嗸�޺��KW��|�ۦd�Wp7@�����P��2]�]�K.���z��#�#��nd�� �����m�^��U'��G��ύ�r������?#_����j���b�&��;J�)C~?�8��+�fS�?����N^0,�q����p�6{+��_J��@��荟�Oh������40���]@�b�NY=�J����;��X&g�]F����
���:�4�ǣ3���:�OT��`�b9s�w�����!��i�j��Y���@ Z��f,BM���ЩW�EJ�yOihVC|����
=����1�dDi��v���4�0ƥǵ���Vk�����۲����#��������]ݤǫt�JiX��"=�3k� ��#��Ǩ{�*�Z�*yd;�{���Ĳ���d#B�ϝA��]f�Ȏ.�KSf!=�.Ԩ��	A����.3/�ƾ��.G8�
�GZ䞚��s�~A����X��B:�	)�t�_�OS�ȁ�&��9Oh�g�=�lkY��� ןu����5o�r�G�����DlHd�mUu 5�yB�"�u}}�hTEY���("'x):�Z5��3?�T�� C�W�k.��ǝ��)<�{[�Y9���]گ;��%�o�/x{�O�T�����v q�u�d��Żߥ�(s#YI���tT[�,s ��e<�=����-,[k�d�L�8�`��i��}.��v}�TW(_�hĤ�^+�����\����$�Ͱ�^�n�_P%�s������^�K��k̀�/j��[k%�\�h�����ёY {����:���yi/Dg��N��֎����U��Ða��	1iP�a3b�G��t�o��H��gW���q���p� �j��J�Uٝ��S3�O.4(ґ�T��2�4A	
�=E����4��7O<�U���!�.��Sԅ)�紦��k�E6�Ҍ��1�����l�S�`=ȩht�)-1��2���P���������G��
�	�@�ހ(3��ln.֍0�6�J��e��w^�	?Aye%�Ÿ���2�9��+׼��i�]�����u��^� �b����,`�4����	�V�����ه��!;�Gx�+����r��z�b3�>f�w�?Hsۦ��8��|nx����-CSGA5	���t95�oC�����-o=A��љ�Q�pb�;z�����U�L��x6o��hC��Ngi����	u#�?�t3 �CI^��[�O������1����픭�:/��]w;�ZC;ו�'��G'A�!�rJ� ����G�l��e�:E@�d8��t>fl�J��+���x�����r���R*����s3�%�������le&*����*��K2��E B!�k$��;�tn���?5�}�{����3E�Q��iXd�����x�^��n��o(�Y$$}�T\ 2���^�^�иg:�'��ؐ���Y�d��s)��SjW�+amn[���� 
���Vpu����s�+1$#g-s�j�V	��%�S�U��u��pk?��4Zه"�&��1r���䮼��Q�.���!ׯ��~�����<K��6�>�%[�x��Z�I��U
#�k1��玃\s+���-�[v�<��zt�LH��&���0��ũ���]��Ҏ�s���	��E�:gP���S��0� �MH	��Sk_h��0���z��L�����k��Q�:7�G�C��c�]�C�$p�;�kPAmē@c\x�W�����Șc�ſhz���n���+^?
۲�&�\Ҡ?���/YB��X��9k���,g	�>ꈉ���� �[ݼ ��
FA�r݃:H��%�+��NS��Wγ����4���Hp+³�X��q�EZ����ǐ~!�C��*_ݫ%"R!����~ȫ���PX������v������l�O�P;.0���� te���K}5��.c�d`�/q�i<���D]�z��Ba<݄� L3-�<�2W��H��![j+��q�S��u�X�f7��źF{.��SBz|�+����ېS�q,�qO��\HM���g��"��L�glom���+��󷌁�"���|�@���!?�a���Y"�	e��oq�v%���ə�J���5 �~���X�V��(/VQ�k�P[n(�_߮����N����/��؉ c��}�bO�-{K��DeZ�Y��g0� ݖ��K�;kޚ�ۨd#��z�=�aA���C��	m"*���paD��2'�j���~��<|Β�t�A����o`�ŽC�+����!��`���Ɋ�@+�/#ju��9����άu}��K ����j����ʎ.�j$�v��aW>�0-J��`����	wm�I������A��.�ƳlQ<��ړ��3��9�Zl�E)±UΟ8��'��}�)g�D}�Ww�G�Z�
��L`M�\k �����z_���C+D@����>�4���Iׁb��~�W_6��������Q�\L�q�we�)��2I^��~B�Y9���p3A縼�Ɲ�cL�"�#qװƚZKF7��Z �m�#��)h�:8?���L@�癆�soȎ�h:~�}��������/P��������H���0�:g��+!ܤY�ȗ��w��lbq���P��(d�Ǐ�dT҃�g�'5B�r��M���su�	��#!zG�rU���4��Rg,�[���:�J=8�|�i��:0�g�Nv��-9&ڜp��!Y@����M�������b�H8y�����4y�q�!�[k؉V7�J�F��9�d�νj)�6P�\.+��Mئ)wn2.4��Yp�Wg�Ґ"����L�Y�`Uյ��c�|0��b/���W��y��/65���5@auE��0%�O8�iT1�!ZG!�3`5�D�t4��P&[����U[�9N���A�M��.D�3BU����3�7�L�W�jP��ߛA�ޕ.}�7���_�b�$�
��-�K["]��&]6��I�˅�`[��(9��暜
�֢(�;�Ԅl��6�Ȍ�:lu�j֨�o� q�c/�%�Е���>�?_�s���Ia�l���0/��i��9s�eh!F
P�5Q��Dg�����n�O9����cT�ɱ��$:v1c^G�J�>��z.x�Zϐ!��=mV���kӶ����F���)�]U�V$Oֿ*��� K��D��.��Ϲg�q$�bn*��]S������&}��X��9�QF���j�难����(��c����uȾ"��1��Lf�yN�"��;i�7��t�1ٵsFc��H��}Ǣ�@��"��xE�O�(�90n Q�r��Q�$�Z�gJ��� 儞ޣ��wt!����pFG����HV3t�6���fHQL���¸��22bb������;.���ܨ��ǺO�g��PJ�D�^���/L����1g�M����Z���,�5�J
��ۥOq��P�~����	�8}N8��(��*ϗu9�Z 	�����4�p	�&��&ĻIE��^��%:)x��ݺUMj�'"�2�h��8��"�B�P�asxMN�^OIMmq�AI��7�µŋ�z��,�������ߗR�<A��sKPZp��e9���po}W�"��'v�;�$�:���rcwc�?�o49�o�8i2�rZof�S�CDAl�Ȼ����Q��VƧ�%m���3��Uy�������4���>K6��4[vp�[��&|��-Y/Q�_�h&!����@�o��O&M"^�ȆA��9q]zI
�������^jsyQG���Jz~�߃�+�(���L�;�<ڬ�5��K�Ƈ�Aa�&��n�a��^�_-�r ӯ�]�#�w�DU�#51��k��0	AC�D�&߹�8>C֤�VȃR��f9����R�ԎuG
GQ8�x%�bb�#�����7G�uW(�/��Zr"E�� �g����#��0)�o�2�� �{���z��H�7@l���K�!Me�i���Qa�k5�Z�ωm���[�~,L�(eN�	�����;,O���Z�&�.z��nR;�P��mF��o߼�u�	Mۨ�¥��G���:���:gRę�8*�U��W�Q�����ר��o�3?;�f�%vλ��%��Q��$=���P�Ӽ�<4[0��،Nb���{��� �f��#�BGP4��
R���Y��	f ��|���Y�/��D���������\㨊o����JE�6B�5��+�"0p�D�Bf^NǞ�S�c�X�	���C�&�K��?��V���$C�|��_�PWh dj�]�vQ��51E��#AXC:)}���[�	�Ov��(}s�^%
�ˀ�^��z=u%|�����i񌞫]�\9���5��^��[jX{��³�7_:JM���H��+��k����G�ǩ�Mm%e;!�@�#�kl���k|m�0�0qH��f_j�4�9`Ő2y�d���1�A�؜k�Ѩ�VC�� ��L�n�6	��4U�6���AV�S��|KɔS0,�[x�N��t�i�	:��2D�>6}^�>ݨ�����Q�3����.�f�}�yM5����KN4+Z8N@�p��[)T���>�N�@���}k��)JS&��m�u\L�%N��<Dd&L�^�$C��g��IMzb�����/����I-�%�^z��f�fW��L~�qr0�ͣ���a�l��mW����B��&��JuREs��RbV��x<�c��񒀷2T�!���y%��p�(P�O`W��*T^/�2H�o����M��"�/9�=q�9r<g��f�4��&7O���X�)7H-[�Kj�,���L.�`�ƹ��0*t�Z����,��4M�����O�*�ë�GG9!��{wȬԌ*E[V�@cdV��I����=��K�p�=J3�e�VMkΓ�H�	?Q���L1F��;����Ԩ�e���x=�GX�^p#x%ZEb��*���e6�(�a,2(a�]K+D"�3Ҥ�5���<�Ҽ:�{�;�5'/SLpu��0ԛ�orْ�J���V�p���;O0���6�'�G���lz��X4�3��8V��-]רv�g��c��@��G�6��/����؇�@��-�/�:�^��R[�y@{L�©g��Mb�h+���XaB��(�r|ʪ�Dz)�מ�՜+.���AA�M]�gw�K�2��n�6�?�L�S����-.�1l�	�nkμ+�g��AW+��씄ϴ�2|�>zK�{��et�J5�!���V�G�r.�)!l�Ǌ*n0=[,|�
Ē���W�Y��gv9����jK����!�k�����1���G,��phw��0A�ͳ0v�Gl��7�d�e^�lF�<������S�H��V^�:L�E$Y9\�\[e��mLNj�Ԙi8-�wx���=ڜ
��d7�Mq'x�Q��,���*VBD�?wk邗Le��3\@_J��Ű�E\��eZYϊ	��U�HȂp5N[z���H;N����1�Bx�N�=�Ț��qޜ��$�N�W��dp���=a��D��*Z�%�Q��i�urgw�k��:S &f���s�^2:��c=A:j��$?���M~~��C�JeM���_��;Bq�&�u�)&8*.���\(:�{kVיn�թo�~Y�#- �E��[�|����v�W�֨��u����]�:-����%O}�k>�� ��z<m9VD��2�2�ć.id*Ή6d��G|D��K<��>��b]�sQW�s���
�<��Ue�rUl��2�R@ݻn�z=�@�0c�ҶAaa|�,��Rݯ��$�-����W𠭻 4!�`N��@-eU�,Ra	�J0�j	e�iL�~$��<��,^�HNշ�򐁣D ��Z��M�Mݧ8��o#Ns�gU瓄���E�s@�z �6�U��9C�q�B'(04[��$֡�
�wLJMmln�]�j?P{�
p�������J�{�'�ba��)h!��'j�(E����l�+f�nW���]KӜl@F�PVj����/z_l��~h{L	Q�j�p0��i���YGn����ͬ�_z�;A� E8F��k��r�����%;��:�YY��p�0�0��F�8��,M��Jk-�R'�1N^\��'���J|ϹZ9�1kج?��"5��D��u�;�|mx ��7�VY2��C�����vëզ�B�ջ�� ����y���H	vb�����ѭ��hW�ﴲ��2��t,�At�QoU��w�o ["�_|D�D���F^,�|���z)��P�ۅ,؃�ђ"̿t8}��`a���1�!Lz��"��"I:Q����X
�ā�0V���;TK�Nu��1Q��S�e2�/��a��z�)�b!�qB�5E�ÌiBs��1�βn�q,�|qk4L�����!�_i��̞�m���~͹%6r"-u�5	�[�uy�M�d�E��m_R����k=	:D��(KWs$.��;�%K������N ���:��߃�UIFt�&����O�_R�G]��J��F���ĂBp�ֆ�d�ů��ވ��'�1\nY�e�'��u�,=��w�|�8U[K]��N��y���ֆ��*�Ѫ�1�*��ZEm��_s����V����ƶNz���2]xb��\�q��	�cd�4~=)��@+���˒�#=IWќU[�:���f���*[xO,���o|�Λ��k���t
HH\�i���޷�oK�T��Ӈ�d��H��@��'�����7��l)Pyݯ�m�*Cɕ (qoJ��b��G�I0C�t)K��߉s	vp�r�MT�~�s[I���z^�ƊߚCT�^ͫ�_��,W�� }3Q��F:�]ZU?-$4��=ސL��	j����Y��n�(���09\���U2*�.O�ɘF�V�=� ��Z��o(q��+.��#&��d$��IHw72�Y%Q�0����^���|NA/���W�6� �B��arV��_�Q�&篱����)`������
��c������eSX��XR
SS�����ti��Y�O�o���h�m�C;M=(��w�c>x��7�m@��h�� p�9s���z�.P���4'հNJY3ٳ�!j���y;(>�$�Ćy ���n��[�`�X.����#��*Z~`
���}c�&*��>wK��}vK��>T�o���^�h�%�]Ƶ	���Þ�v��/m���� ��;x�����LFE�.�6 �^�(sFP|�5��_Hh��z��&����X�ԕA�>�(��ӹ��@�H4��\�����?v��T1�HX$�%����W���[k>j�[?J�\����>����2F�U�~��U31I��߶��p��-��jəT�1V��x���KwF!�k�U5���\��Q��ߎ�'�}�9s9W֕t�Q��8����ų4�$�����}�G�(5���n���%�'eT ����s���混�՜��E@0C��sP~c�5�q�u%�;$�A�E�#�{2^ݷ��:��F������W�'�lA���c>rԅ����g7�-�8��X�4��5�E�~IT�$]z#��"H��-�~^�����$�D���0����"-�ՒU�?�o��Й|8����Sz*Iw�f��r��U�޽F��S��[����b������;���B3a%E�d�N!<����c��0x���5g��Y>��v1UW�]"N�֐�-��<�O���N��ƧG58Ŏ9�|�ۭ�,]K.�sa`���g"�B�%�"E=
<ϝ��u�V�{�͂�"XL/��x�zA9��w�*/0�մ�F�d��i`Xl�vE�r�mD������qi�샲�`׹�meݩÈ���'p:C����ܨB�q�=DxWm3�e�V�<
��L{���MҸ;!�����'y/��7����C���0��Vf'��ǖ3-A�&�Lj�(���@}"m'�k�߰l���8Y��d��o��&k&�<[H�y&af������>�­�c�#?/F;��Y��4:�5h5���@(�����ђN�Hz#X��[p�Cb���Fb�E�iNAؙ 7E&�V�?���"B��C1���l���[����r�6�����I�l�,z���>�&"ċ�^ǁ�N�I�;�t���yx��'0&�Ѕ�zU��Ks"�:���*��
���F���!l��c!��������~@Mq^�F�Y��Qo3��M���^�N����N�OrA���gi��Z���AE*B`B[�Iep��ӻ����ۂT��KKy'	O��M,D3g���`Y�}U�8�OG��\Ŧ�	�׻|���C��X��+�IA��c�Zv�����g�Z:I3�~�/���Z��OJ��9�zBz�eY���AdU�i$[�ˋ�m;]���{�+�^��6Csn���HPE[�'q���_H*���A{�N���2�P�~�J�-��EA!��J&�#�N�$7����oD�!����rp?� �X���<�u�(�"+�4������}�R��q�5���b�Y����&��t�U<����ٿ�:,�]�?���C����`�:��Ez/W_��G�WS�[4�P�P��z��$6����X�\��BYO8b8��`��>b��+:�j�R3�I����P����|Y(7���R	nW9-Kt2.�O]�%�	���'�|c�Em.On�9H>�HD=<L�����N:��Q�$���z2��ށ�6��sWA���$M
�NV����X¡)z÷�T)�]�hj�і�W@v6��I�Ғ�7n�XD{-՞�QP��V[��lC,/$P�O���Fd���cd>r�<�Zmꑚ y�z��H�	�ȴ5�Nr��	�WH�u
��B���1tt��N��l�X�����.TEu!����H��!��8*>��HA:ь��cޅ�T�}�~5�;���I�6Hz���K�ӝ��#y�
����"��[��t��L�wk&�K2�߿t�sX|>�&M�����$I%��"l���KEoo�V�X�Un�0S�i_C*�/��""��7J��v��h'j����K�`��rX��д1M�׺V����'��LY&2���Qe/����.6/�����SUh�Y#�x1�����OYI�����Qg<�VøZ+8˙�8�]����rƿ �a/L�D��iB��ea2�f�V����6��@����0��ݹ�\h�1�<v������LК7e=/P8��H=��'��A~�����Q�Tt���2o��gM�(x����؉S�id�d��+����lqd�d,�k�:B�m�jh�PTYY6E(�l;/����uhٙ�m5�D.���u��S���~V����,�'T��=�_v����}k�(���v�P8�}	���*�5�� �a�
�ۘ���;�N�3ߪ�~�bF��nk�gG������e������]�*��[�T����"e�}i�V|��p�)w��q@*�b�A����xɒ���x�éW�x�Q�%��[�a���hL 	�4g|��;5��U�e�z�6�xtKk�+t�z"�t�`E��	?=���^�d)�>�I/�q�����a�'��x3P����l�����
�ywfxd�����w��lr���5��H�4۾��4t����°�ǃ��u,>w��� \����J�S�<�cKW*�u��K�c��rH6Q{m�w��e%8�s���-3ZU\'�<+���S$N��c�Y����	ܥG��������`(����eX?�e���Q�(W�ܯ��8)��>U=5�&B�%��:spQ��r�9��/tT�:�F�Y�Bs�d��8Io�@&2���U�?�Q���],�(���b78:�f2�\S����a�55��t�r+�2l�la�C�&%�Ąt3o��Ab�n!�h��~-ڰRyy�<�6	�o��Ũhټ��9W�1���H��8(hUo�}��^ �5G���j)�������Gn��q��J�,�?n�0T6�A���^2(o��r�3�=X���7{i���7;�[���`���.�bf_�	�v�A]��8�e�C���M�`�N�^�D�p�N<�dݶ~�m��:�x%��RBq�	�+Z�N�R�"��a�I+(4>�Aف�L���J+����; Ƀ�N��Rt�>o&�p]W]�md;��з4o]s'S���w�&�
�!�(��� �	�(!ۏ�ta[N��1�m�%' e�z֚�j� ܹ�H��T�����`�1�`�X�Ĉ>Z��e�Y'w�&�3Y�a ц��&��q��O�~
���Ȅ����\6yM��I��?�aI(t��S��u�}��xrTI_a�gp�Ɨ;����B�2$��<�P�Vo휙����2�Rr,�h6�����P����	�p����(��_����J�%-z������U�%����@��y�?Xa��
�;eA�=lJ�3��� ���,v����I���>i���68��?���8p�x�U<���G��vQ��U� i	��ۛ)�ܙ0�L[{Y-�1~��H���&��?�rчS�KM��Έ?�ߟ#`qR"i^]�Z=�j};�ɛw�Sv^�m!_���yZ��E�>˫����p�N���凌�l�?и��G��A,H!�?I��A2Ud�EU ��x��βN�
 (�&hMCfE������G�r}��ț֒��؞7t�lu�#���z�,����Y	c�z�1�j������[���S��ܵ�ï�q%�hhSW��U[X)�	{�KC'�1��7T|�^k�!a1��W����K�;P[��-H	Nfe։���ͶE�'?@;pQ��A���w �*)�c��m®��K�3���R7Ɉ�ژԚ�aB%n������#ǪS������
a!."�Z-�GS-�3�WnBqo;�z�Qȟk��K�Dkl���� �3�gГ�Yܙ�`7�z����Vk��#��[tn�����]����C�b�+�SEm�1젭��] ������ȡn�R������o\��S��v�������9juEs�Vl_�)���A"�_�����8H0�����ȗ�c};��[�r^�S+�S0����*��/ES|m����xx��F��W��+��UvL�	�3��Pu	[)lκ�	q`�5��e���[��G�O��S�����D0�d�(�J�Q�����9�`>������~����0��& 9���QQ۹�?�b4m�WI��;�����n�1ar5��r�&$��2�7�C�*p�x�c���~	cٴ4a���ݩ�u�?��xE%�	0�b�����n��4��gQ�}φ����o|&�f�pT,���R(+�×�V��t���,�̌�i�g�B�$.Xލ�2A(��2>��nJ�t!�"�B>m�ɂ9�y4P N]���E�XH�W��� :7g���925��d���
�a�F_UN�9й��i6p�\׳%�[񶗚턾�	�~89�ȍ~�a�⛪�d�l�����)7R"����@�$)�`��kP)�/�V�N�m
���0Uf�^��s�f�!	a8�$�q�����h(&<>�IW���*���X�0���ͤ�l㵱-R��}_~Ry�)7���,yh���ȀN�v�e��ӝH�PbZ�3���,ψ5�SU�!�T�u��7����.X:JfhF�Is�~�/�i�fO�?��8t�>U^Å�@�7U�ty�����z���E[#�5��QRH��z�.�a���K�y����~�Y��[C�ܑ��q��q�\Ur��o+�8�0~�&��J⼤١ƈ�Jnz'�E~g�Yy�2].uV	d#e��DPyU��FX�:L���o��� Մ���Y�)���=��9G�_"k�*�����p���-�~���)؀�p�!����ű}]_*}��Ly�g�˕On&5�7��v.ҭL���(����%�f̃��{i�\�ґ\������W'�%V����*�"9��A��0�%c����G�ʔ�'�e8y����{2-{��G��H٠�mY�D*C(E2\v��O��+���;B�D�J�/Е��܇c�EV�Ս����%
 �߼N�f>@�ɞn��ޢ��q��2�G�?�B:E�G��!f�ii�X�EP��.K�L� U��L�R�%�6���D�^5狁@��-��6k&�c"`z7�q��hl�Jn��WN�6�.I��A(�I��Y�x0��7���'P/|w�.|�ɟ�Y�O�C�7m:���q��=�	%���:���B+_�VxO��s)�����ʜ	�~��2%�n�C�0F�%J<��R�!�}�\��8Q>i��f��D�����s:7�����g�u*- 汦]�T�Y��C�t�A��}���e2:�o,�Ga;�Y�4�2}�
�<����j/
9ɐ96���c���,(]}	�˾�݊�3 ��~F!U����5�v汻*=���$�4�~�@�%T���L�<K}_�)�.���S���Q���B�ą�
.�3y�ܦD[����\�MG	�S�9P�߷�Znٜ8kH�r���N}�9ӛ>��n��\�.�3lgy:��C�7��H��!n�#Z�	��6�Tk8vPߌ��A%��m�����o�r�SA�B�'b��À���>����FZ~��^8!�w&�i��[�W���3,�o�P*?A�8
s�'|�M�w�ê����U𩼥���v��܊ZaI��o���7[�q-k%����P�n�}�wj���T�3<��#F]́{�j�^'�Xp7B�@�!��5ך��s�˻Տ�-vw�*E����z[
J<A������V 3ǫ��H��O��a&�O�c���KU�����-�ފ�����U��m_uFyvN����������b`�q�u�Y�(�҉��_�'"��B'>��;6�2���0�n�oIzG!훕��ĉ�%%�i���v���8V�{|lG,���I�åްTZ_�;"��d�N��>��"<�I�s�����v:����w�1��L�#��X���
 ��y���:�=�k �
�� @�Wm5{PVy�LZjNn�0��}zU�<��O��<Q6���)j��R�+0���(<���~�}J�wh�oV��
3��#*K7�k�W�N�]�V�B�^A���4�w@9g��9Xbg���/���hPp�����$Ӫ�Gi�b�H8w�$��n�#������Aߎ���"���,U�*��f\X6m�����=<ǧ'� �%���J^�#{��A����J'�>U��s<>1�#�b9�d�(��c9��܏e�1/��U��z�&$y��(�#���jw��Ƙ�`�|%4��q�s��4��kp����N-��S~�hk57T��(:���͚{�ͫ֐�KFڤ�A�m���d=�9
+M �|_�;��v���r�?t�#Kx>�>�s3w['^�g� �k/�Q�Nu��q���Un�sVW9ʭ*>��q�����H�*��X9��VXz��Ț��!�}�g5���I-�FC�A�"�\4�;=����������-_��P�|�^��7��M�I���Mkr�]���6M#��͎������n����[/\y��G[8;������-�،L�:�*E�3m>1|F�%e�gL$���^#}�ݡ���	�>�q�D�Gi*�������$��L��(h�{i� �(X>��w@݀�Kg6�o�����JSI˳B�7wW���ܞ�[����O���Y�NOMїݥ��WR�B,��J>� 2����qzSJ雐H��_����*���m�&U&� �d-���p�۷��g���,&��[d#<�Z��! ���h�)cO���`}��JyFi�� q�W+1V$���v��[)3�����:�K3�8���+�[B_)���Jw��s�8��M�li�(;f�� �i��q<�.�G6U��pѭG�a��$�����BM�]�/�K$��e�Em�։�^�X�C����O&/���Ė�4��y���PM:�lhH� Mb.k��ߓ��/Qi��B�r���ҁjU�L2�~�����b��,�K��
�K-@)o�[����^v�7_�� ��{�����$1�*%}y���r�@�ǸYS�x�*�G�YK�pz(ux��h!�W����?ۏ�����CYscu��%k�X���'X4�W	�k�cQtnÉ��C[�^����/ة`/��su��#C�U}6��xYۺ:_E�l����3l�~�S*��j��L}�'��Cw>�$*�z�>�U��i���y�k�����cȺx6v){��4E�/}�E�Y�(w���9J�EB����.�;-�)�"0
��.���g��
�J�Y9m�-]��&�z��Xs���T#��hM|g�a-����s��`)Ji��r���<"
�h|&x���[�@��˺�$��$����h�=% �^X<��KJ�"�aF����"j`ȷZT%����\���܄�?(pc�j�Z������#��ށ�͔�y��[b��� ���vxU����k5M�[pe����|/&��DD�`10��̅�/o�ۄ��!�q��N���Ǜ�#L.$N-�)9N��7�()�X�w��q���BJ��Q���d��W�Y.���rzb���+-$*�=��ϯ<�0k]r���}su��~�H�Y���R���- ���U}Y,�P�;8�§]��ߢE�E���b�o��0�����.��6�C�*c�1X��B],u�'���s����na��-����>��$8��7����mx��e�̌o�p�yIK�U�bu�,�,K;���Ub [s���,i��Ÿ��=Z揯+c�ڡeU��0+ ���[ڴ�g��"Oq�r���z���%��8Ta�sJ�����5�C�q����h�
����c��{�y�H�.W��QދP�ڢ��ǧ��(7�
�@���s�<+`�6;V%+�y"v�e�d��4A�������&i^!���B������4$������� ���B��
��>z�:��щS~{Q��3}agʐbɲO�T��qS�J]Ac���f�ج����e�����S��w��vbn209%Y�,9.�����T�kE�Ux`L�=7��&_ɳ��mM�k ���o�/���^~&T�NU~Ϗ�]�����rX�U���Ć�9Z��ɟ��?����Co���fEFL����o�#R���	hڍ����ٙ]��t��U	�>'���z��6%iĳ(d�{2'�����f��_�j!IڇTc��+)&}��ɡp%pz9 ���=�#�B7��M�̽Q�yc�LV�0��;^˿@BK��;���6}�FbV��.���k��Ty˾�kHYu�'�{y�'`.��U�x�w��0An90�O�G�⺤�x�31���7�K��L����vvǙ���w|�T�V���6&@�3���-�D����D�K��*���͘+���XI����X\ *e�|�hz� ��t�7��uXAo
X��U|s��³�8�X()���;�V��$>-/��h(�{H��e'�+?���vŦ�r�<��k2����4?p����pL�����Q�U/��jY��*u�;���?�^�V�\��%N��������{s�z�H�L��V�Ϫ�5�H ,$({��\ݸ�4�b
�.΢�^�?m�見�U��fLW5�}Rc֔ʕ��j�qsS'a�b�L0�\=�rr(�T�lܨąWhP�'ؼ�<#��Ef�r�����	"�TN:h�]3름�-�/Ʉ�����	N��O�LO)�*)vt��E%�ޥP+��&���K͔�v���&������� |�'���dT��M��"���#���wO�G��_��>�M��I{S:-�h�ͬ��_?0y�����;4�A"�I����iY���Dү��p$�� �!�O���ֽ*��k�����j�����Li_�Q;;�4+d�R��M���?����9�[���#Nݣ�iǵ���mO����O@�z���D�uf٘ߛe0T!Ɨ&Z\��5�qYS�[|��m��wȭ��s�/�W�V�-���b�%�	�g�����/�kpSgґs�ʈĞ�V-�K�|�w�NMc�5���C��u5��k?������$�m��`�j��?B�5f&��g!�S��4��tq����l��R�B�D;�ߜ�0�������G�pQ%j9ւAPV��#%@7�7�������u���(�ە�Ky�����	!?L��?9K)���,I47F<$) �C^Q?�a&D��z" c���4��%U�Cɗ5t#��
 ۥ9W�"=�Y��/�ļ|0_�:���kEFL��h����c���8��9x�9>�ш'� �*���_D����'��jPk���Ji�!�2�{�c��E��e"2����Z�Aq<q�	��#CU�MԼE��TK�c&J�w�L�����Ur�ܢ�`=���}�%�D
0�xol� �UIgSv���8��sKJ��W�w�7�d��ߑXj�I�݋���q��8��c���,���
���p]�`�fRtB�~N�cS"ji4����;ԏ�c%�4��|�wI�:��r�A��W{�u��O\�K�o]��Q\��0堁�OR�H��=�CLP6'*����+�*�aHK�7ʊ��/�x���u�M� 9��-}"b�A�r�J~�U�I,:�kTgW��,yu�>�o�����#�\�Z���<O�5�M)����ݖ���ٻ�{���·ں�P���V���H\e�!����ƪ7}���<Fj�����,~��+�&�����5Fm2�>�$@ �;E����?�q�(iU�=���a�Ȼ���r��f|�<�����d��ۣ|d>��вR=�k?�w�x�$K��_�Qg1Y������c�H����ݰ����M ���H�$\U��j�3�����R��qժŚ$���.}�t�M3r���|�>/Ϲ%i����~ʸ��������Ed�x
Q�A^���	�� �I�b����>&���^t��U�ą84:�{���'�7�3��tb�x��m���s����%��u��'d�	�Bs�/��S�ȣ�J�7b�n�w��Q`2�w[/P0�0g��kI\����7`�{��g��1
[^�u��&LƳc7�øF��zw��2w|N�Y3b�]���8\�u�UvT�<Cϰ�F`��:Ɨ�5 ׼7hL(����+�/tŵ�M�.�W,-�5Y�+7���٪�T�2Mv[���d�0)M�9���7N;�p[��E��f�M���w���z��8�*��L�c&��0��曱:�Oȟ"��u���YS&�;�B�rN��?v&��Ԯ��y�����9��;R�(Ԕp �<�k���wE	lN
b�x�E��m�V�O����!���%�/(y�6��<��f���6!���bC�`l�5p���ݔ�f���:->��q308э[�8��/'�����Mt�vD��+P�A7��h]�!��}��, QJ��p?�J���m>�O�f��ks=����]����� 0�j�C8=���V[//-��;V�I��c!���[Ni�v�t*��']>j��Y1W��z�\R��D�Y{F0��SD��6�G����Ҽ���򗯝n��i�n�G�O'	�}��ub�Y�3�����P����o��yc ��z��� ��_�l��Z�g�a �q���_�o3�[����o�۫��6�ӌ��8��1*xWa�h�W����:l�L��Xg���t�s���[�=�gL��O?UTkRF4)�`�+��TJ�B�z�]����jC���V�w�M�'G���ȡx�$w�ъJ��O�h��+\�B�;�d8_�����	�3��
=�d�`�~}��Fh���.�s���@���%:���3b�R�BҢ�6��]z�jn�T�Ig'��ԗ7f*b�TJ	���݃�����znZ4^�&�2���(@��Zhh�8?�x�⨫�Hb�lE�G�M f��;�C˸�iL��'[��ؚ.�V`�b��T�N��0J�ɴZ����t���Lh�9)mK�y>�l�����x�H��d;��۰��*��!��<��	����"CY�;<5���7f�}6�$QN���m�
���L}��5��8��!��L�G!�T��6]�ajޗ��\WL��NO��?5G4n�2cI4b*���`ٲ!�V�^�v���Ɉx��Q���Sb��G�����j�:n8��j��E��_F�]'OxZN^���(��	��Vr���4�^���4M��<e)��]�7��I�;��]F�T�f�eb�3���״byc����e�'�C�w�Д�q?�	�̀r_^�'}�ޓ����2&��!� \��ӷ��F��Q��˒k?<�I"�^X������b������t%��.w1�2��[ࠟ��[��s�fq1mH�`��6ďx>!hm]Yq7�5�<��?]��y��F;�PX��lɘ���Z�"���R̝�Ŭ��d:�7dP G<U|�ku�<��up� �){%o�D`�T�(�;6�m<�Un��x8	�񢣼X �}(��<ϲ05��a�M������X��Ґ�T��
l=�[#�Ʊ=~hfF�p�_.:<vm�����p3��n�� C@E���H�b��r%�HYI���Q��]0��90=�}�jBc�仝!G�P+�)�ש;h|W��b�cV�}.Rw(f/���
�ءM���\T�=���l�=s��^Q�_'��-�'ᐄD(|D���5*��ćuG9�L�ʟ Q������tc!;Ȼ�e:--ߟ�箼:5��U7���7r\���@��kW�}z0���A��bׄ������	��R��3BA��"�+���\����s�*倴po��6 $��ә�"���U�H������6G�Vi]���Kh`.VLu<��բ섂6��R.q��78j��E��o�$�~�k�:h�D��4���1L:@����>o�G�V�+f�L��{21��l���_�܁b-wV���.):���[z	�P�O�I�
F�r�_��Od� �(�L�PF����-y�;��;8�w���a���)~������sjc�?��ᵰ�'��-��Ϻ�
+�_S�)7+u��bh��4�i�9t���aƳl��-m"��R���=PEUIl5"t���]�pm�:֥ �G ^�Ղ*�L�U0ȇIx��_�/l4��#R�@��/<:�_"{%BŋU���?%�M��Ҿ40�R}�_�������a�C��|Y�*5�=�Ew�Ʉ�B	S �S�{�뚤�_#��x�f;�����N��4�ϩz͑����x�^��ǚ\�|8*��Oc�o�/ $�B��4�]�F�����3*�e��{�Wb8�nV���i�5,��'�-3�}@=��1�gwṄ����!���|����7h7�牼:)�������Sv�׹>��j�Wq~�`�ᮩ�%����P�L�6#���)�QS��TF[H��w��<��7��f8������܄���C���1H�i��0�"K�M>@����@!�9ĝ�Ah|QƠsOX�F�L�G?ݰ�|�2��Ñ�j���S�:��t�Cb����£����aV0���d�Gl6����L� �-$\��y�߹�9���<�\�2�Vs���=�-RzV8��p����ɮ�w-��IS�[�=��	d7��1wC�/�_���*R�&����$��Mj�fR���:��-3f� �n�!�7�έP����)D�7e'��|�0b�km���n�����҉.a�����+�$u��3��s�H�V)����m���������iﮇ�m]2s��6����a��NҶ�r��=�� �(�ޑQ=�xd�w��%��׾-��G�w*0���6A��Tb�(�C�$�X��7�{D�O|wj��/�:m����O���]P(kD���l�tdDvrȈ���XqI`ʉ�O�ʗ"���:��`js���C;+�������&����2k���CK��L�p����ԓ����$>Jf|�&J1u���沔�mӮ9�ҏx	:�A��l���n%���3��gy�!��Y���-K孺ɂ[��"|Գ�ΐ��^�9͓︞��Ç;ȗ_�sӰ%�/GT�uq(V�t#u��B����/"aq=r�8��oF{V���������ښ1lh���FAH��i���L�&�v�eW'@�9xME�F\56��p������G�0�C@��V��R��V�	����a�p%��k��l"`W��8��a�%�K<�;2�ܷ��f[FI��JZ�Nܐ@TW0�ؚ4�A�h�Q�yAdxx���t�x ����im�	h����spo�B�f�;N�7�����v�lW,�(�a�_t����LT�5�Ɠ�o�����۹�#��m�F,�|UP������?e�o{b�F}[�����F`e=����Ǟ�]eeZh�H�D���=�ש̈����/z��xl)�V+�]4u�*$�۬S������R���֏�#���"�2]t���#��P���iZ��ݢ�1�_?QqW��w6'~80Y��[��
,�X�3>���t��v���O{�>�q��h<�g�T`���3u��-Z���!�U�0\x��?��[�5���D��
�n_ұ{�=�R��d�����"��P��f���e��z� 4;X��H�?���?�0n.m0&��5�d���6�i��Ĩ�a�w����AK�>CC�<U�?hke�qI�D
o����CO���֒d�&�dy^��Ki�{�a�㘩Q���~�V����V{�ېD��ُq;Xq�K
�F�r�m�E�>y�OwI�4�;(g�5ՙ��g�h[�&;o;�O����|��=U�&,}j]���v�ՋWv~|`w���4�e�
�� Hn���ާ2޺r��I���'�%��N���D���@�!�s�9eo29&���z�h�-��=��&�aR�F����s�A�6P1�}N�x��į����Ƒ`H�#��9�(^٤ ���+��U���9�-���(��g���͒$��H�j��=�M�ΝP�E�hvyu��h�z�jE/z�i�A��cyJzRATR&--�L��̶	0Q��?�r#ꊂ����'6g���_L�s	���x�(�0�\��DN�ļ]� �O]�?��cA��ojL"��#6��&I	 \3�IAb�;��5��0K�4y�L�&���޼��ݽ� Z=���U3�����7�Z��8 V*%� $L
��[��I��yX����_���P�i���V.�Y+}pp�zHc\�@̌�G�7S_�r�.�7=�}%���<��F�Q�p�$�MۗѩS�,��t2:<�O�@s��펐����UА�M9 b���؄�F��_���|/�"���'L(%q�\)���l"�#5�pߞ����j˾�b��5	���7R��ͥZN��%��LA�@̑��-`jTŠy��x���k��
Y�pt���u���@C/�I?Q����&9)�Gk�p�O��ᏎW��(?px��*��d�5T�Y2���.	��`���85��KM��e��m���v5�8��¶M�".�qש�P�F���K~��e��࿐����FB�)�=:�z̵��t��3y[	\�z���bQ�ҦHYC�RԠ�_})���Q���~��e[����"ˠ�>���v���e�B�gM,�1��Bل�˺غf�JSe����g�D2(���!�m�U��5��S���i��]��ic��(�r�5K�)�D�	jT�-�㥕5�Ѣ�d�a]���)EK� �{�>�N��9�cz���*�{�Q#�';�vZ�f��pէ���X�x�#G��W��̝�v-�տʣP%Z�WC���{Z�H8������������W=�G\sp�B�6aqѤ��~s��4���m�!Ӟ!�i#Ϡ����"���e�uu"�<Z���W���s�hktF�,�.~u�� �Vi��- �&Mc1` �&�,�����?�<�Q��Y�y��Nw	P��4;�?H}�In<��Tt�}
qV����|RJ
�7�<S��1k��_�x�
�.���%n���M�'�{�Oj�pVT�Q:Z��Kp�k>�[oK���l8�#��"���\���4�̨,�������������'�(�1�ލ
ԩ��(��'�.�̇P��.s.�W7�ٕ	��#�U��/��h��l��9/f�ˢ��^P�K)	�]�
w<xsE��)w�0�������ɕ��ʰU�5�:���08�� JH~Đ8�j=N��؍��Kw�oG/�5	���%�g����c���P�ֲ��	
�����
R�.TiU8���J/
X��6��$��P+��H�A�i�/��m?8HSe?9��Xţ������e@��k
3����0� ��� �l�Y���y�w��'@�����hр��(�{��~D)	`θ�1��.��hO ,�U�y����_,}��3o��à��D�P�G9q%���3!u|�C!|�U3zc�f��C�!J�P���U�1� ���*���0YFY�5H�y�Ѻ����@,O�Psk*��p_PN*�gN�X�]1F�6{�W��mQ���	�h�dvN7j�	��)C��<-:7��Jt ���kj�5d��z���x{S`�AOCld�']�dn�ꀵ�'B��oU�d�`M> �?O�2��lj4pYhN�����(�`�9Q]�qG���qt�pvãMWUl)ux���\�!r/�s�pΏy���9wߪ+���v֟��d�����"��}>����I�@�@���e*6w�`�ʪ�NƔD������	�t,TX��|ϑ�m��r���R��6��O�'Q	�qn��>�QِGz��z�̳g���Lb�A���=���V�D�6�)Fe^|����Y;4S~(�� :ﱯ�+��b�έ��9�t��[���N�i(�t����c�e)#�D�Ǯ�� m�)a���t��&�T����G&K�ͻp�.E���;si�h{�gn�� m@��/$�:���2��g�:�ߖ�5��\�ēm ��|�5oQ�d8-��+�-�Q��Z���i\�I�����g�@��l.������]F�Mڍ��k��a=�xBt�}-]X�R�T�X��z�2� _�C�C����2k��c�"].�fA� ���*]����9��$?�����Mӓՠ6P=p<�f ��XZi$�z}����$�^� �+0�7SK��� ˁ�5[��h�V汣�^�Ձ��
'��:��[������r4��P�ui�nmy�h�.��c�	I�n��.�Q�|�x�d��q��ܹ�˩X�ʕ2��+q������Ž�͸��
G�4�-e�����?�A-��_S��'a}�$��d����ɜy�:��p0�Ƞ�X��j��Q>�=���a�8�*�k=��Mu�����3�U��N�9=2�}z��M�"��PX�!�Rr+���D�T6�u�n���_o�0�jl�-���������~H~�~#��"�*
o�&GZf}��� �6�7]�~�LT��&���3�X��4r�od+|�)�<<6u���Pd*�XAw�m�
��Y��g�Y�I!��~3���U�%�j��n@GC\[$�ac�duy7�~��k��Tq�ebKBJ��\3�ƁR9���H��x�O�[��3��ق��Z�=��|.6K:W#�~�R������~`Ѥۘc6ɩ4�,�e`��v)Ӓ����d��8o+�����v��)���GG϶� ؅�(�Y����~�ݛfⴧ������+�CJ?W�|�V0�Y}_�C�g%G�)ۏ�qAh�Σ�^	Nv��$��]`��m�>rN��]́�� �a�#wlC�&܂��w&�e�<�|╄V��r�aҾ�P��zz�Jl	�ߥ��5�
�=�嗒���.}����e�
�����U�h��AJ�+�Z�M������4�_�b�Fic��#L����j�a���s
�$�;�$��9~�:n�낇472���Ly�x�^�����L����Pac���{x5P�*�2u�e6=��I�։�h�c��eMC���d�[w���%,������s��K�k�M����������`�������諵_D�{�ްH�p�cB�!
�81�һ��Ã��/������n��o�+�����,e،_2F��+b��D��hއN;&$�wa��e����9�"����y�t����qBQT�Sj�û㠤K��ɑ��
�t����-BǱ[��a1��k���f�i�I���	�99Ԯ�
�.�]��6~���nخ˷)���;X���U����=�8�^�����C{������
=!�T|U"��{������h�K�,�W��6�^�s�8��)��[�k��|���C�ώq	��2
G�	C�M��pA��hK� �6��g��J�i혾��i�����?P��|]�QUn0+�����&$T����]`\φ�ZtC���dE'�]Q��zᱮ�D�x��Y{K�s��t�e����+�$ӂk!n���I*��h���r.�t6HcXK~���Ą���6<����zQV�=h��%A|p�e��]���O�w�ؤ��J��y.�}��˪�l$��qmy�S��3z]�1�g�6�((���Q��w��W�0�UE6�Wq ��xV�����Gֳ*��p@��<�<'s�t2а�n(�>-��͔�3��/K�m��Һ��OT|:U�jե`�)��݃�k�]�8���L��sb�S��Ɔoy�w�ꥥ��mtF&�:���xd����hz;�*�&�EQh9 X���0@&ˀq����!mh��I� �&����>Qp�O��&)7r���`'=�݈\�d���P7X9�4�^L�h0�)����${�c�h�F�fMu�Pg^A�+d*ΎS��!E�#L��G�a%���Si���L�������Xt�˘ e��(80�Nv�E�P7�L���}]0)YfqE�x!�����מ2��S̖iŸ�`&o'���J�5�&w�������XT���c��[� n�\vG�N V6��Vo	@���;�U\t�E�m�iz"�aju/	0���@ȕ~���!�tź(�&���!�\}X���D���:/%J��xҪ�Ti70v�>����+M�T�=�>Z��B��
ٷH����D}���l���ȷ�AR�9�S�A[�@�.���{��Nt���!MF����Nj����T�INz΍�g�g�l8�Z�ΎodR|�I��D�߀��sN�&��5�,~�9Ye^<��CSj�7LlG<��F��u:�z�v	k��c�+I�)��@����=.�})<G�g�����տ�%��D��PF��#��9x��_1�8Y���E�l���<�.J�1`��3�Gİ0="������G��&	$t�׿M���݀w�U}	@l����zVE��۳9��˨v6�w�U_�!�� �$�=� �lih"]��{b���	�q\��A��J�<�����CU�z-���{q�r����C�"c*m��gN$�0c��&��9᠂�t�������$̷��������,u@�m@xl�&�x�L�f@i�V%V�|.������Nɇ�G��=9��K���%� �'��d��� &|(��'!��!`��#I
�= ^��x�%���jI�5��MY�}��J�0ƾ:�.�>�o��A��6��񅁄bw�W�*}܀5԰Ñ"%���Ի8���4��q)�,��8e�{d^��p�M4�B�3�����Ye�_I$0�j�=`�8���i0�ٜN��e�e�Ҝ����@�w�E���0w�'~�t+�#�]���F�QZA��ޱ��'�����K�V���c��ͺ��ʳ˸���uqJZ�����,z2��e1�=x���.W�J���Ш�e&���l!8<�*g����f0p��.,�"�}�� �E�օ�,h�Z���F)ٟmY=�������63���-�Awq~Pb�6B��5T���Q>�h޻A%�}e�N�3x*��C���N±�Bp������3�X~Yp���9H�`�T�ad����߾�(̉�[�93���J��lI�	l�k,P0��
V� \�6�wRP�:w2FÚ3=J��D>) 37~���y���&8�󏣌���Ζ ©؝Ǆ]h&Ok��E9&J�[S�Կ#�D���^Y�����R@j6�-�̷^�W�u#�?,%@��v�"p��!��>o!��4&�ը�5���$D\^:J������
�R�d��� ��<&��������U'ic�wƝ�5�����DL�͔J=tk)mӇ�1+;Q<���,�[^���<'��TDPY�Z�I�R�z'�=�����<En�'��ടR@�"k�	�<�_I#JY�B��uJ�y�D�o�]A��0Ys�t<�F��LmNtT�I�Z�Bы����X���
����d�P�h��@
"tEB��[e��R�s�I�p�k��:�2H-�#���]��2LET�,3�2��p�
�����f;�|�Dߝ�_��6�[^��ƃ�[���r�6�|��n����0*��-<ID]D�i�u�|�K�M�Z��J@��j�<��r��<7;{n&NW�a���Vt�]��-���)+����IX�iZ_,ʑF�m����W�?�͝ ��/������B`~�|�Z��yt�6�P^�(������`68<�G�;g�E=֍;���yX����9��F�A/�(L�n!wF{B�3Z�-�{8�쌈D�
�f�$l V�T�㲞k��X1$!-�c"ӌgX��#��jgK�]��.�\:u~:�c@���A���{����7h���"|��C���+���WPA�X��n
c�/�,�C��������s��}���2�d1��,SỈ	؞��K�tB�UT���Ɠkok�'�u'�a��A���I�R�j�������n���KMڨ���;�dp~���a�[@�&\�z�������j,�_o��?�:���{��� ��c��S%��-i(���=.l�/i��Jx��y��q ���MWΕ9Bc&����e&ǚ�d����4x]Y���g�}U�N�c������� b��a�mʚ��m	�k����tc��w�M�p��gZֽ��<<����x������k�|7B�$����=�)2�-m@&(�ʵ�C�f��V�W�g���L�L�:/�������.��͜�]�����y6Ԕl��y~�0�BҩX�͋S���V�f�HH�ˠ�,�4�m�uWy����b�7uMw)�/�_��I�r�J�Ƙ����f�O7�J��3�j0yQ�����J��8H��	w�qZ{���f��y �*zz+X֧�t����a�o�_�e�--�E��>s59&/�W�T�1C�BFufii�HN���\�os��ë_bD[���Wth���5K��)����m�������Y��͘D6>�
(���6�-4iV^����,g~w�Br����1�O���}�&���I7ar֛�c�ț����qq��	tv��C��`b��u��8C���9ƞ�?��X����D��O�1iU�Crס�@��(�#D��P]6�{/$�>��)(�YN{��Yf<L�?SY�'A���d��N���>/�y�3\Sª��F�*-	��WT@�����D�ڏ�R#K�?h��W!P�F �i���gDC�(�e�=�Jvq~�O��8���N�*l��;�n�9P�
�teS���D���)y!�z&)��FP/��m�h2�t�"
x}D�����ag�T�p9y���Ӏ��q�������ډ%J-�[�RE� �U���{Y�S�qЅü����H7{Wl
u7�m(L$�k��OG�a9R�r�m�q^|��X�������lX��X�tJ�j�����P_��ė��e;*�S`{��*u�V^1�����Ц���j_6d��g4�������Zޮu�yq�B�FJ��P�V�+�q޽��~�<�gƻ�&�	�r�d��*�Y.pI�ȼS�3��҄��M��0du�@���(��ˋ3�laL�ۈ�д~{!Fxu�������A9@�f�h_���Qi޺G���ur��|L�*N�^��� ��Z��6��;���Jma�� 鯿kɲe�kz0�wz��RYd�Ntȱ�M#+3���=�9�n���p�{�v�d�#��It���0�L�8��<+����]*g�v<���)��3�)y6�/��1��5?����cH���v�ŵ���8�Xu|�k�$�p�x������RY�5��^�Ò������l_�]�{t	����ono�ҿi�T�YY�M�����e6^����2i���2!7�x7�?�[��!(����%S��F��!*C���u��~����E�����^^C$h]h�$��w��� ��5�����S��NR1�]Tơ-B���d]zO�c�p��4Ф6��Ŷ�\tZ��&O�Mp����~<ϧ�v�ǚ0a!ڳ����j��	̚�ó��������{�B�fu��eiʳ�
r��D+���N�+ �p\6����Ez�3�E���J=J6��Ov���&��X����׮D� ~�?��Č�X��9���b��:�{��S9����]�4���qg�f����I���1eg����o<X�0�d��0���X��V��&�������C�4�A�b�C��$��Bƶ���dA7���N��5�AmY�[#k�|Zk�Z��26��3(m�;�om����C�y*��F)�cK�:4crc����G���R�o��!���=�r�Q��ӏ�^��s|<��!�ԗ���|��(69������/�����d@�9�{*vy��/���~T{t$�#�I��i-���8 t���,o�
���b�L���lJ���NXغ=�4���m�U��Y�F���YO��\e	��}�b"���x�F�>_��'�/
�D$`\L� �7��7�3�s�ϹO����,~n���0i���A��MRY�ch�+��Y�sV7)�S`�NW���(;F�N�9�{�� �'�ܯ��D&�_��`bΙG����m�My5c�I+�n���m��=ݕ�+{�T/���:�D��vP�&��"���o��W�x�q'w��:x�0�� ��6��"�:iR9�,�sƢ�2:��Ԙz��6G���G��k�|�V:���#i����*��׃ V������n�_��Az��I�QlX5��4�\ۥ/D�A�N_��'��eB�lrUA. �S0^�azQ�3%��d7��HV�a��;�	Fɓ��d�cC �L����3}am��2k'��c �fa^U���j͕Rҷ�:A�O²��coH��f�J(�o׃�
s�l��4���K�C���p�@�5�0)�j��o�t��2f'��������b��)h�X%��q�fO���vV|�c(jJ^&��=V��c_��)���/��P;B�[�ۓ����+��f�Ĝ):. �(���*~_ݳT�¢Þ"`;Mk}y�?# l�`��2E�����d�8lP�A!��sjh�d�.�2��Ԟ.�Ma �g�����߻C�Y%'���B�c����2��ȮC9%��E�K7z��!� �n�������ɥ��B�A4��ͯŁ��xj!����y�����Ϣ�w��O�F/GN�lnߕG�2(5���j�ՙ]Gy�t�m���QGn�INt'�V!-��I�I@m���F�@��{1Di�D5ioĈ�?���6�+!Lb�U������[+i���v�C��
� ����������F��S%>���ȑƓ#7|=���mL�"bv�]$t�l�V�\�~��J�	�~�j��F#dת�����ɇ��.<`&�Ib;��@��q���B�����c��` ��DG�6���D}P6�4<�މ�>g�Y�8�nJ�B�NҎ��v�F�#�'�����-���5���gP�:�h��??<jA�w�U�>�G"�Ɲ�g�	��j�}pP�Z�0�[���&ԡM�H;v�0�^� �4O:.�XI1�Ș�ʮr"��촂S����%�����wYC=�/�ᥓ�t�S�D�������~�� ���Z�S ��.�xv�HlH
}HRՊ	,���J�/��wR�\βtʮ`2}��,ɭ��D����xk3�<���4�  �o�3`��eN8���xo�NQ��D��2ت*�I���)�+�m���6����y ']�nk�P��`r�J��,��GCsV��<���e�iM0d��I������"�O�A#[76�)��[e2iE�=�M�g���:�LF�o���+,�K�o��	��;G���X��/���@Ҽe<�ދ�|����T��3Ǡ�����JYf�Ek�)�o��\�3K��k&^�wm��0��Ϯ��Zy�y��[?W.?���]W\�`L�z�窈h�3ۜ��f�~��c���Lh�d�U�5��f���S<��F����u�z��L�2mɎ�������m�(��!�*,2����1l	�����/�q�Do��&}/��J�/<H?��{-��mG� ]-6��5�MO��8U�;ū���j��1��փ`�E�h/gҥw��Gd��K-�s,P�)�������?0�H)���Jh�AAZ�"���謹�߾����}� �9�������.�H�VM�7YC�d����k���N�h��x]��� |�Dg��/��8E-��|A��\�,�Qb]�	
YU���q��ƬHϭ8h����g]�^�L��t�p���������}�{e�T�W�⽲L�˰H�<H7y�f'6z4|�
[�!`<.@�,P� x�0r����E�G�l�����)(t�^��[�������D�N��E�Nڊ�X��w,���,�d�&yg
�gg��O�CI���>FC���Y=i'U���'�3޳��+�6˿]ApzH���.��>�<S�\��LрB��&y\��5-Dc��x�0��T%����Y���jA�~�@٣�@���� ����3�#�T��W�
oj��3�N�p�����S�=D9���yɵ�f�voD��� /��@' <��wGI�OV�X�%8[�����͛�%R���3,#w�O�D�o'`cJ(��bMX���JR�/�ߙ��5'B��6<d}g�J��5g�f局�êu"ÁD���i�i)�Wcց?��N/��K�N���4���̅$LB���>UV�>C���e�\r��/�L%!u���KG��Ǜ��)�6�:D�GT��W���!#��d-?ގKS߇�>%6&�S�k]��fB�⥺�M��΁.��^�2�;���d�p�ZT�;���W��H��b��а�h��K�2=�̀��d���J�4w���u�$a�i�w�k��MT�|fIH�a�W�	^Kdǌː0bS 2�5���	�aNy�ᡂ)���J�Pކ/����lbY��EcM%(e����U����\�G�c~{�w�_L�Rm�!˿2&�8�c��ϱ6O���;���:�OqT����v����,�ZE�>֒���8�Yp�SK�@-�ζ�$q^�"\wO	��<���5N��QJ|h����ֶ�`�p>"��BaY�o��b+�8�j�V���[�7�E �=�T�~���t�ɖ���R�Ə���͕v_ο��6�>];"ꌁ\	�%��4_M@R��?�s��Q�Њ�3�����F��`J�>��΁>R7-���cw��G��a]�M��p�#DA��D~��K6��9FvS�1{���w�-"��� ���Fx��mq���u�^�&�zF�@_휮<Y�2e��O�\(�-�b �c��W�H�|6�7��}kT$6B���6 �4k3!�������W�p{�@��)@�BH��g��f�#U����ǳ���猗���͑�����}`�DP����|oeP~��Ec��Fk~1�>8c���Y?� W!. ��� ��j��%ᄻU�Nk�����M��#�*ш��D�e\�*�O��	�+�׽y�Y#�|4i��f��9��'�5��t�yn��p�"��$Ӣ�bͶk�pW��g�h	�hk�M	�;�J���1]���tS7�[��1�ߏ��1lQ�6АT����0z,��('Uf~��K �o�4;wy0HIa^�N�&w���I�Ш�aywp"�Cs5��Ci��)?���Dvğ�HX�z�I��Ԥ�r~Ya�P\q�Z��P���o0t��&`9j)>�썋�:��z�dY�JS�W;���&������ ���Ko���3���nh'��ކ�5�/���;l>���g{1'�`��&�@-�e���=�Z%a$�V����A+r�i^p%f�����é��t��g<������{�Ć��3s.����Z����5(��P��}c��i_N]���b��Wܭ�E���
����Jg=��(xI�wĮ��F6�+�0��/���h�e�X�+����/�j��l$ГT���eKz�/�+����u,�'���|M['��	�ͭ1N!�G)��tcm��P��_l���*��ջ@A%k����Tq'Cw. ��Pe)klْڐV�]����
�G8���R�D �~��������%��;���@z0�ppB�c�)/�L/S8�� l�/���a����W�1+�R�K�(h.3W�Mn�̓�6�y2j|ֱ2�(T�p̻��xކyg���g��4��{4�Z0UʡYU�2V* _^�C�a��vc|+�6χļ]�Uп o��]{X9��t�՜���b��Q���\L�z��~��� �wF8�?i�?E0�w��$������xc��4�BJ@��ԩ���$t�����E��Q��k-(w��QO��!�째ہ��k�Ug�#��������nNZ,�ex�"���ɞw%�
�94v�q̞�Hx��U�F.-����3��֣���QV�XEj �C����uT�=�`���� R�����dz�� ���k�阂92�vZ%c� ě�8`����_u�z��u�E-_��' �ذc�XG$�.aĥ��)�r�S��ڦP��9�r�/�K�7"�K-`S�'�k�D�9%��1��%�+�O�]�'V��a%��aZ��9�"��|�ze�)ҟ=@j߬���޺��mYqRyC��Y��Ki����cP��'�Ŭc�-i���7�y���Gb�nc�
���P�2�4TY�`�@�¾�5Jh�M"�6�ʛ���{�1�V��R�*�@"�5��ܰ}��ªd�������Q��f���ӟ���5��$�_e�J( 39�M�f�̘3R����ς�oa[3w��	����_Ո�(��p�ږ*���b�w�.GQr����d�zƯ 6V+��ܴ�jq%8(�D����/�.�0%�i?�0�}��y�y�uvj�`W�wݦ)[�<`H
2�ɇb�x��PKL��'aف�9d:w��y4;*G&�O8���&�ᷴ7��fl|��iܑ���`MزC�7��pl��"(E�7�o�TcH��d�C"n.�TP�5������dv ��>[#�'��k��@�[���X����$6�y��
��L�pX�?�3����I��Z�%���̵��.�DxF=�������-Vɇ���vx�`#Y����~��JrJV]�u�0
��r�n^:D��#�ݼ��Uŀ'�r���T�aQ~�z}r���.���8U��t�]�]���4Ѳ�0[���`$ي��g5�u9�Y�c)B7<����6����Lj���w�a�4#!��x���!�R�As^	�[�̸�6�"��ܙS�1+��v����bXvl����g����׹4��d��K�͞{C@��7΂�[E�j��c�".�Sv�I�M�5F�1I5�J*p��)���
dzd�5A��>cVPhS�8���ҕ�X��s��Ku^V��9�z&<;�B�4-O��xP�ޞ�4IW\b��z�	�VC�`�(�huR
�;L�h�Es�� ��;����2]j���8���o��9��ǫ�"��y���O�Oh,� ���~�_.���Np�І���-�Qwa�,$l	f���~аyL����[e �wV��ْ���6��THj�+~%o��"���,��!�8�-'���yπ�%͒�i袖��>�������d��`���w�B�V:��S
����ry�S0��5y�9G�����! ��//ʕ���������wt��\�x���F�3����ؿ�0�BVa�ۉ`67��G�iU�t���P��˞��F}hY��(Tk�,��L�4�hwE������~��J d}�x�GU�j��F,=��rM|�>Mf�_QXl����6=�=Br�M*�����tc��$�z)r��,.%�}u��WLvP��^�>]��D�iu�%S4���|�"�A����MZ���e(�Q���E>nZc\�Ʋoh"M��?i�̀��ˁ �}�[�f�0>�2����ؽ^h4�%�jֵ;W�j��M<Vk�CR7�I��.�Gk��җ��Q�v�ԻN7�8$���6&V���2���GƩt��|Ť�� i��8Ox_4@�i��-bk_��"����9�43���Q
A�1��FK:Ā"��S@���3y����䳅{�(RMw��H�X��ķ:�NWJn&s�&8P�����X�Z�ƳiD8C�w���S$
��j�Xm�To��֑ �*�W�g視xaր��<�Ϡ�Z}��al�*L��OG�&r>u�<[r}U(��.ĺ%����=q��[g���X�O&l/��A%�f:�ɸ�p�&��Om�F9�}�=?�p�ѿ��s��k`�'�R޹m�L�g{�B�}��rB��y��`�xUt��y���i�"]��A���R#X|I$k_���3��}1��:k���"��b;�q��u~��l
HtkY�tm��#�o���YZ��%�Nd�d>��HLK7�,`j/�3$Z�:xG=g��MW��ld�N�S��x���h��ҵB���c����xM�g��1���*"P�}��l�j���%��T�F���>�"e�^,�_m�:ֿ��6���!G*z��%k�ZOP�S��ku�N�t���&��.���R����9����P		��G�R��	 Vw�(j,�g�@�md&j�m�2-w���G��z8�9-�4K���<�Bx��֨ޙ ��m�ZϕP�g����.x����L�܆�BI�.�7Ae���H�Lv�z�͜�_�"��-ܤ�)��ʘ4�1b����W�P�@����q��6�~P(�kjn?��龠���߶������J(v5�k��|�/� �f�o�aY)��&��w6¦:/��ZSE��4#��j�����S�}�,�q����5���f��하C�
�O����~E�k{������O��i��P�,�x���7'�oN�Uĵ�5����|��EB�L_y��b��I��ji�DR��"лg\~ t������Ff��ܒ���m�� s��wj�r����_���Mp�M����;Y��jG\��D�e��XR=OL0��amϘ����ّ������1r}d,zk���ضTy%�4��5�!����@�۪G�RTql�ji��Qd�� TU�^����CA�Wbb�B��G�{� /����r�vox!��M\~pKB��6%1䬻{
t<�L���^k�{��Xً�aO�X�+�CI�b�T�+v���S�R�%��K+"��bS���<�!n��������ڰ&Q�h*����-"!��)߰�����3��騫�o<��?�*��X �ֈa2�(.�R#=q�~��Ӹ�klnM�]�/��q|�� &Վd��x������b	�4Y�J��"��3�*��u�>T�#ù��=��i-��)=I*m�<�0��7Թ�8����xmD��UL�'���"'_�Ӆ�2� x��,n� �c�N�p~��>����]~�����[Eܷ�%`wz�=Z�%[���[��w�B�^��^� ҮFN����˞�f��5�j�
7�+�>Dw��o* �T�ԇ�<��0G��+!�O�i@�3���J��:2y��}�~��.s���z�MqgG^�yaQ�Ԋ�t�����6�`���3Չ�(��a���^���J�؉��M$_�7��q���d$
4�vd�߆ҕ��aip���V�E��.�Z�v��������!vM#wU.4�s��W@�j�^�f�u�Ć�Hpa3��_���IK}�E�FCUM���6{�1��	�S�h�>}�����C7��C�c�8)pe9Z��"�k��:��S7F�?7�e�H Y(+�줂�}�Q�Y�/��������&�<毄�8�v�"Z�gN)7=��upl�뎙�\r�N.xOh�����٧t�Z��l|W�*��H�5'%!f �4�&�g��MϫN�Z�]+���ky��E���V���u���^`�� e�h�`���w��ik����Ql�Q��3l9�Vfe�Ыs�B�=���ᘮ���Xޠ*�:lgP��d����y��d�$�w/N��x��
2���/G��,s
�GՀ3�E�Q�؊c`�y����G�� �ʌ���ہ��;m�Dj�G�������1}��y0�u��o~����+�_@���N^D
!��Ҕ�H6@H�h�t��:d��,<ʁN7��[¦��Y�G�s�r��`�O]=��>�[:ō-�%�b�q+�tRh\�A	�6��,8h%9�NY��j՞���)L�$���A��	�}��A�\E߯"�T�W��Ak�O����a���)�__\���+���`���EwXk�
�7̎\�mwR�QՒڴ�Z;�&�T��P�X.*�
��s�j�%�'B����;��Uĩ��\�v^jf�V�2��^����Y*83����a	�;�[]4�D��)g�Cf"�Jy0�Lq��7�mu2=�ځ.S�Ϥ�>������g+-�b�-��9q�q�)�ќ�{},�eM�[
j�N��f-ީP>	���#$p��C��2;�!P�W����d���T�����I|�w"%�vc�%#.��HV��f��+�Z��A�tu����|���4C����ݱ�U�G^h��y3D��4ʩVf%x���˪˨{��\���ڤ{�D��{�pY�{~U�W�z9�j�b�6=bɀ���zu�Y8�	��i�y�W�#i༝Թ
j$0����&H���
��F�ͬ���`�5I��T>X�x��z�lNq%���J������Ÿ��#s[�f���Fp��^8��1Θ�߂ur�l��j���N���T=�Y�;d��t�w��m�(��L��'�LR!n�7x-������+!4p�L	�N	)�vW���(|�����`��/4��wxr:~o�����h��B~ӱ��Ձx�Y/�$z$F���%�H_���މkD�D���IHR,�x�E�Jd��pMl�Q��i�4��!�ɇ���,�1/�oG)VU������؇���>{+J6�1%��<�_����:i#*���.~cU���<q��Q��l"�,Z�;��~��y����Q^ٗ\P@�lX|i�>~7�|4�+�����)��py��8/c9�0A���ڼk��L
�C�x<1�=*3+� ��~��q��`�N$��W%��9����յ�������ņRI@�Ob{>�oX*"*�7̦���ܵ�A������6F��h�i�� ����DX���. �'���7�}tz=�JZ�\M���h�)k��欅Q*3�Ib'���&i������:8�a�A�O��r0�������5�⏹W�]fgZk�g(��-� �ɰ��<�ƻ�A�F� ��>t�G����L�١�f�ݦGG��c������Ȋ��$��ӿ"$T��J��ڙ���������an�P\���.�O�-�UM�<&�r�V���t�.�Pڥ[)�s������#S��b�a?���wG�l�3[�NӐM����W��\+�d�.���aW)7����<�#ge
��3<�G|�Bz����Q��%���Pǿb�T�+$}�j�`�m�g�)��1�x�[�z��a�y�}sn�-s���K��L�ɟ7�~�W�Zv����Jh$lB���|��$�/ck����Қ�LK`�{���*�w����3m>�sU6�X�'Jm��vO��/6���W�gg�O/����Y�ާi����6�e{�r���K�%#���������8[ 	��h������i�]��_-�^BuGH�g1�gT��$���g��o5�?���x�9��w��9�h�%��q�@��3�Q	�8%Xs��&�*��˽�hh��gյI��ݪ�]*{;Fq~_`Cr���oü�����@o�Tl-A�Lg�����嬞����̎���.�n���(�L���!V�\XQ}�OP���i��N��n���8�h�yI�⨪m�%�.��juk�)��.Q�x��s�^<��'ר�a���N"V^�g���,����V�e���t�7�gߺ�>z�����Yf��\~5ΰ�j�6�)�K��L����$o������D!����(�𺡭_���$'�˃]�Ewm��I�G�^�	_|GS�f�v���=��*@ՊI�z��8�Ҁ�^M�u?��H��1{u�j;c����K�W�wN#G7��>�GB��p+N,�UP�������MY��6�YÉW����E�V��v"�?�i[>S�"���z�	�YyMZ2��*M�[nʃȦ��=&�����e��������e3"a�t�| ݜ	c�Y9�%��N�ޤN��B^���G�K1���!}JK�2�%�8�����s1ƎX�Pkg��⋖�t"O�R��{-@
�����h9���KV~R.�+���,=/���7ƋZ��]�OCv˸V���q�J�F�(d$��w1,�� �Hֳ��2U1�a�K�,e�$Om�6����Q�%G�`���1>��|�>��7�L�Քikm7(�j��s�l��E� �L�v� ��S�Cr��H]��O�%lhP��$��mV�Y�����a�3��t��w��$c�B��.�a���Vxq&[����J��(�����u���I�/D�����B��+���+�ΩO�m	�rv�_�[Z7�F��'��1�%�Ks8qX�|(�Lw��tAJ�1�O!t���Y&b�m�H�S�h��M���|֏��p�O< �W�T�].��K縥ih�Ձ�µ��O��!.�z�9:`���Kc0����p����Sn�7u+�}�
*K�h�d��gz�ۼq;���i涐&��+�^����m�P��q�(� ��Q�m�)#��;r���=�o�a�~w����^�����W:��A`9�(]fz}8#�����m(�F�\s��E��cVkE�ζ����d�1����m1�\3�����0�݃6%��Um�Oӄ���i0&�xj?� Ȉ���ǪHd���e.��4�jf�o]eR��o�-��{�%���?��YYڨ�������}�8pb�o݉�8�8�ˊ�}�V�פ6�i(;���zTW����W^�W�f�p��i��kp�Z�6C�Ù ℀I`d4y�+vp̞:	y���u
��D^�LjM-�͠U���{�BY� ́���6מ`�q�RA$W>�Ֆ��Kf<��;z�ŧ��B,�{n'�3��r;ґ{f�"�`�u��&�ث�-����9��x� ��ѣ���V��ݱ!	�Z&�Ոc��퓨�lY/L�q
��nٞh|��En5D~
����رl�< ?2�́��B�@�H�`�UD9�-��a҄�&qa���|� A<R� 6��s����`+5�n�2�^*�)����~�a��Kv������P�r;&�Q�O�>�N���0����$5��«��k���?k������D���#!XZ�)��p�ç��!�8�O�?��&�T#�n.��&�)gΞ)�P]����m>Ѐ�J�T_�;�`�}=f��(�:k]�l��覱��G�B�6�D)��:�\Lq��E9~6�]t�P4G�T��~n�rZz ���^��]pb���غ��׭�@�:g���&<t�����X���m775n��-�I�5������-%���T������C{"Ǜ�Hj|�e�+aO��%i���R�!�]�;��$$e��)�&�{�t4_�c2T��B�IӍp�te���c@�YH"���*�:���ם�-�߽��W���?l	0V�A �e��c��B�u�ZUk�t�x8�B�آLV�-ZH�r.(L)^4��B�K.I5o���|/C�); �"k�΃M������z��wn9Nn�~�$;N�$��q
k���T�
�U�C���%��:�8<�<�%�p�C.р��AY�[�"&uCEKA0�QZ`ZB��0d�F�k)��xG��$	���{�BG�I��Q�^N�<� �d����X#��;Q��H
@d_� �ֈi��w4��?L�D�PIC�P�sV�rlځ�{��/J�Yya[��;����/��$�K6y;�%j������nl�M��y���T��&�e�����������k&�3c�e�ȗ�N����D��*hwo��>��6'� ���!�����VUTس�;���)�����VT��'"����i�^
�n��9,R�dcr�S%�4ץK{���g��ǌ��W��lQp���	Wa�����˻�ur"��*�'\�IǊ�_��׌:�7�zwZ���xz&���[��~�F�|�t�b��b��l��R��&��N�)��B�%���ɨ�g��Fצ�Gۤmp�)�G[�O�d��͛0K�����E|�9���	�k��iO�vL��hp����G��aH��դ�J���F~-pֽ3�&���5S_�{��.��'��KB7�_��]@����'� ��g�iG����a�y%�el�/����F��9�j.���fQHg�y,Α��I��ݽ7�G�2�0�=��s~��*�5�x��xc$�xfz�(|�4'Z,"Kx,(�*K(W�̘Q�f�ŋ�?��`�)�F#Ԕ����3Z�7��gӒ��/|q��~�]�+@��3�,tW�=̔w���D���Y{˃��T�n�c' ��M�&�S"9��,L� �9]�Ҡ���;�s���c��7���L�=2e)�%��q?j�)ě�th�����*#�,U�{fBۢu���>���*����|����F�
!Jkk�v3E5�1q���]��������{�M����aq�v��FpQ`9�;O�@!+�7��Ma�M:� �T'E�� �ٶ�Pq�H2���9VO#��L�������A��@8@-�R�6.�:���T�1��ǠZ�!�̡��e���4����g��9�*�#�� <Mv�5'�}��#�Q:�Ç��cM��ƈĚ�ZJ�$���JbE	V��A�1�A)�_%���l�Z'��Ң{ͥ����P��l+�yA��&&4�V�M���p,l3`���K�/_�ߖ�rZYw
��î������B�7_qR�65�r8�gl���UB}���1m���׿���!wK��}�$��Z�赯q����J�
�HgW������� A��R����|�{�'.���!΢Yټ���P�+V��6e��8�(�����z����w�OU���RJm0P�5������hK����}ǋ�y�_��>ʈ;��s�9Gq���U�Z�8���\ԟtsc���5�_ �=_n��rHp�͋�M����7W�><��0L�cTx�s'�V�I8*#�?�T!�T �攳������R�	��ݫU�����w)E��0�\�Ue ���t�^V�ݠD=��� �!��o�{�_m�]��������G�^��u�  �|�NM҄� �,�>G���<4�	��Q���4�1j��v����47�
�^�i�?3�G`�4M���D6n����ij�F�F�>�lP�n
���aT�y�b<���L�T���{��s\�D���4���mQ$��3 \�*Gp�*(���Ř햐�V��e�/
be���oVGcm��9a�e�1q}�0��£�:�Ǜ�PtT`$�L�;��8�iz�t����I��X.3�Ȍ���s��(?�˫o.�g^��
	1�Ua$.e3S�N�ԏHsa�6�i�
�.yBj��@�t� �6;X �Z�{̓J��j�V��In?�.
U��":� �:�ú�� �WW	�Q�M����L����������/�j�C�?X[4��S���<�TI��@x�e���gע !�Ĭ�R��Հ��|�p��}M� �Ƶ��gs��n�	:����V���+��rj_�j��r����V��z}%GoB���al���f��侀A���q���5�K�':��ȷ���Zˊ�Sd���Z�,#��npl���̄!Iy+9>�e�]8H	�ء�pg�β�z6U�h�������VQF�`h�i��V�j[ip�^u�e����'��3J2ݠ�{~w$�W�EȆ����T���~9f�=�g���D�5\WY�S�U�%O�<�~`��/�-Q�FQ��m�ޯ���H����n9�2�(�#-�串�Z�S�k`���'$h�z�=�oyΈݴ����@=��%�I���~���_��$u7lkm	�`�;
�A�v��s(UiT��7�HZ �k�Rd�]�ã��7%U�A���) ��M��S�MXP�I~�%Z�(^��y"8EE9�*� ��2l��M,0LzE@H)�w�Z�'@`FB�.K|�yՀ����l��xC��x�D�Bs�av�}̠v&�ial�=5��m� �Z����f`� ���^}�y���jޑ�
�PW�ŷ���2�V���`/j�NR� ���%乛a��9G\�DT
x�-T��.�x�H�-���˰���'��|r�x��gQ-Q
D��9ܼ)�*��n�1eA|�Z����
��UN9��#5�y�xq�<�������c��e����@�Łn��zX0�q��쯗s�pV�\ef��s 5Q�`��Opt�`I��,�����+�
ɥL���zn8D��o0܉�$��x����0�d���!�]�TC��MFvs*Ao�~�cwS.ͱ�D�����*E��'��Y��Ր�o�x���L6�rni Z���IuЁ�q~��h�����l�t��M�^��[����Y�Hs �P�����<	YH�F)!ޑgE9���GF� �y����Xù�˝�-��{:�t�3CQ�v�I���8�"�,�cr���lsFP-�n�\y�����?q��X�Gs��rya@��κ<�yC.Z�����ҟ�T/�b&h�7��S���q,JN�F�Jeҫް�?f�z�Z�_��"y�?��e���h���r6��K��|�)s�o���7������X"��U>iog�T+�-�-iQ��ͬ<�Ӯ�lg���*- L6G�BLށ[��/�xE�vB�Y=9�9� |�rzw���y��#�OTR&1�z�Yx�y��?P���EhPd)T��ʎ*�]�[5׏��q�����,i���7�$W��Ǡ�9������8��y����TP=*��җ�/&��f�G+���
�CK=�bP2v�3f�..:z�����=�*©l���ѱ�3?�.y�E%}���SiI�vv9��:k��,"<��\\2`��3Й�qk.�����|U6��	i|VK/e�I-m���iЀ�s��w���ti��1���J�o�1���8v�g�ȗ�Oo[��	}탫�k�5OJl����ԓP���4}�|��Ps$Rti�	B�0��k"�2kmw��<���ð:�����K�f�H�S:���E�l!���� �Ѣ��WO�p@�*Q�:5�aj���eJR'�@�'TdD�`XO��Md��K7zB��əM�^Y<�p5�2��4�%=�m	yo��ȪL���`��F7���:��?C��BɅN�Կ��4C}=��f�8����e���#�3c�W49N���O�X��ל3r�$�6�'�� ���X�˚ң���ղ��z��+p��3]r��m��SR�e�f��W,���aZ�.~��$�bLB�r����h��h1�q ��2���[��88��� ��>��z�o�6Á�NՐ����w���>IkBKi#IW�js^.8��CqX|�?\.SY���t���T/u�&�
Z�@�ua���eʧ���s�qb��7�?�����E�<O����Z��!��,d�@<L�!�H�>Z������@�*���wwX\ �J��I�a�e������(�~�Q"�ۙ�E���NK_�����X� �(�j��L9�# {�ƽ��6~�C}��Vd������"���D�D��v�/:M�}�2cW����\Ni5_�&^��KɈm�%��<��R��࿱!���BJ+&wx6�W+�wR/�-�*;w�ο��]i����l�1�a���bܝ���D��g�C%bV��ȪI��H^�~�B��9�_C�Z�2F��1i������C2�0 �ڏ�4���07���3܍G�#Ŀ�Il\���y�x!G�v�|��csi���m�2��F�76�b\���c����ŵݖ�\��x���h�ZL`[RR p�xR�kC%��y�\ȹ��`&���%�T�᭟s�#XdR�Tն�,�]V8$9O��f�*��*o���M,�k�C�pt�IhlI<Hu(�4_�rj^�i��v��EL��Nهke���X��&�/�(��
.ǈ b�>�&8V���=�ڨ^.N���a@����Bh
pg�*��+)�= ��?�m�z���~{r��x'�ʋV]~ؖj���lJ�s����a�����RdN#n�7xO�`��	xqQ씧=�|�������T����H�q�2��%�`���O�������KQ� l��%�u�t�2�Z�i�0�&�����Sev��YΉLө�7Y���;�C��P쀧�Z� ��N��� {S�
y�Q�'r�V������,]�F b̒ր����{�G�v���H�6�hZ�+��GYW�K>���G!b)����������8,h:���x��
R�6{\+d�����05	���D���P�S�l:s>U+��b	v8�S�:�]��|����_�|.k�^�-�+�$�ᇶuD������"�I�N�!���(��b0(�fv35/SO}[;?<v���g!EPR�֌�� s>`�T0@�sܯ����?T�:�(g�3��Z��ﲺ��<,�-P�O+4R�Cۿ�Dt+��ڹ2
���0�)>X���L�vM�}�V=ˏCe9��r����Ą�����nOb���!�.QuG���u����R�@dx��H��!�cK�b۷��c:m����K�o�s��[�x)��i�me�@�eok ��+�N_^F�L�KM�5�*$�	S�P���{ҭ�R���Lv�����{�JtV:��Zu��t$ZmΦ6,�_��`�ᶕ�}#��#��gw܍�gٙ(,���8;b�*����x+�#��.���9�ޱh�׼�xi`{]>���UH���͊�\�2)����9jzL��p��U�w1����8�I�3��&k��H_&�ۄ��S�ȌP�!�w�Π��U�~���vJf��7����
�~��2���~Lz��-�W^�{-���C������H�f*}w+"�ꭢ����=��-���`F���h��
2���Az�ɘ�����ͼӲ���B�>{���M��7C��q�	�7�Ҕ!�c�#�����x�����OK)��	��n�JY�1��x?Aӛ b�l��7M�˦���6�]`|��.d�>:|#Ƭ�8O[+|�㣑?������!�s�v�l��E� <#F� +Bom��8�#�����3��������z�v	��gčj�Gm� �OCk������8�&h�2?u0�d9�z�����C����lG�&��Lvk�jr��P,�C.I@��]�� c.�L;�R�x��k��>r�A�+��K�4J$]�)�$WJ�J艳bC2�PK�
ݲG+pŐ���ڞ�t
�H��b���q�[�&�ĉ tu��_i���/*�Sc���Ƽ�-�vE#������� -<�����3�"��_~��\eb�bcA~p�,�wt�/��f����Qi���v/��j^F�Nɭ�#E����ūN8t�~��y�޵\B�sf}�Xt[�+�G�u�wC�ɄOOD���"4�m�3���knب�T�����.J��	ùz��UηXRo��|�	�v��H
��]�k֚�r"� �����P��O,����ӭ=
��?�I�sSn~��{v��Ҫi�c)�C�����G1']�3��T̊`}tǱ�_OW�|���$�LV���Aɽ4~���D����YD�s�c�N��y�َy�v��y2���T��d��(��ڇ�wA������x<.��;�6Uϔ)���.�c�*/8�Х��,��q�g����2|���g��Q.�1;n�b"�&X�E���eo�QҬ�,8iؙ��F���͋5>���zw�nH��~�	x��P�Z#�"��/�+���waY�p�8~������D����9�0��#�Ϥ*�m�m>j��߉�G{��3
�C�����(�:ƥ�����W�T�K��L"<��pؿ�T��e��B	��t(��6fU�<,�`~����P3��u_��4�D}��x�D8ּ0�@m�b��U�yn��TE7�{�"����V\j��3���|�m�hhe�4�й�K4�\+;;���T� &�HG���Kf�P+�:;Н
���Ǹ��M-���F�C^y���r]�G3���9�c��o�S�?^�Ϯ3;9��{A �?��"<�vJQ�X�'�Q��Yu~� ���F�nWR�i7u�3M�`/��o?�W��#o��ސ:�_E$�Qr ���6�P�O�`	����M=��/��6�$�(:�%Y�ہp�cF� �ϝ���!�|@�@�����I�I�VLJf��(��[׎�W�����a��X[�X�y%�ʀ�_D.�%�YUb�7��b9:��D�	չ�p]�6]���?R��Sx5�5�y~���ѭ�� �_5���{�з�ãV�����A�����$���a��"O
���lXf�������a٘��>�R��CZHTm����b �O��ٗtB><�r2%I��v
]���D ;��i�h�]�4�,��h��[vq�!i�}Gv��z�J�ж�[�]��tU�QϣTzl�Z��W�zK�Uޔ?����r%�~�gP\�oiF8]�К��e��Dʐ\ ������}���A�)H�Lѫ�]J�� v���؋�~Y},��8w����d��%
F�z���I�̈́�'N�OEtH�*�B���;%r[Y��O�(�w�ប�b�R����?�\_��Q�%g���X%�����N��\�q�Va�>�d������P6����&���<��5Mg�X�L�c�C�2#�&�M>&� �tMx��$,���v:~��|(;��XN��2Κ�s	�ú����)�tQ�4�Wj�zĎ)`�o�q3"�|�Ip	WZ��x�~0���&�x��o���-%�V��)�A���j�/�������h��l�&�A80�Ws"W���}�`�b,i)Lx1�0W�6�����NF���m9��s�[��� ��/s±��N���wþyd���\K��5[��bp�3�y�,҅��G��1_�f����
�B��RJ���8L�$�.C�6��㜑�)7��/�Y�X�B<�T����Z�F��'���~���@-V{�������-����۶��L�X�8�!?���!E���*Al�<Y6��7w>��ux*��E
���]"�Eݮ^�n�?�ϩu# ��u8�"�d�+��	x����a3a�[��NMp��$��ܘn����B���\��jp���O��������Z��Y;��w��l�:���-����2��#�ݨ�r0�*X�d1�؝ ׋532:�!6���I�3��z ݂�=?�g�j���6�2���Ƴ�3��q����D�w�~�s�o�ֳ�%��.�����nێ�U�����;у�U���w�0%4"�O�z�[�Y��S�:[:%�b6�����`��9����~��(��Ξ�SW:� 3�5%���2��7S ���"�3����*96��зQ9�'��_�Upu�� �Z�?fm�e}`�.�E�[\�l�	t�2�n��}kD�ev��̑�0',�;IS!P��h��'J�}����>���D[T~��3*V��.6��-%tR#�M) ��I 1=b춝�_���*5s������Z���e����L]'�ə3�A�'AdomҥU�J�.��J��R�?V����!�g-�+�,Y�-$����s��`p捹,O�)f^j�f�$�"��Zrv�r�6Z�}$OG�Ǩ��zB2Áf��88�{M���Kض��(��y�ǈ���5��)��b���O��^��p^Men0tߞ�2��\f2�T���f Fs>6Tj����LT��G|�t�����{�rbǋXQhN�l���(�lW���a�d��]v�XC��<ؠu�h㻚@���Gt��7��@�����(a��k��PW=�BˇxS��io}M��Z��}Z���M��a����;�-X��r+��W���<) ��p�N��+��>�@���g@����l�A)fGA��K�0����M��ԟ����=�����%���V#�M��S�1c�b B:�Oì2^�qHKν:!Egc}�pv_����S����T ])xrǋ����\k�S��0<����GW������?	�7�����,�:�����ߗV\�с��* ����L/Ԅ��*_a��u��K]}��ݟ���4���A�A�����EI���><��茳)L~(���[�&!�[C+��^�K���x
DϬ�;�u�^����PS���`�K��1�H����h�{��I<-@ L�{���� �Ne�I%W�i�������1����/��&4��yba��z�r�>�1߬<��6�ԙ�?%��e=X5�tEy'����>������!r�ge ������L�~���r�u�l|�� � ��N�����hX��S(ѫ4��\�mT�� �,^��U�4�z��8PPEˈ���f(V�=AЁơ9��t<,@�f�H�u�I�7�2��k�p�Pj'8P�{�V��\E���U����d����Z?�����*2(9�-�gJH����Rw�;ll-��/�����H� ˱��O��3���w��"F���TrP��_��o$�4^���R,B��z�onௌ����;��Oyl�<�2�Q��HV ��p�U���/Z�*��KVs���xJ�\�>�4kDO��0z���,�{�P�����4����K5�+�T\*]����]��i�g}�+4ܿU�4<Kv3���va�[e�ݔpY�2mzP��Xun}'(J�d��~�(t{%����ZZ�&yY"Q����σ%e�L�ǝ�O�l!9� �>mQ%�yc��� w����z�wj:k�1�3��-�ë7� ه$S sm�.Q%[\X���Ͷ<*%���b�?�'�_=oK���Jk�4b(������˽~		�颪�n¿vMb��������/"3X5�]�U����M��{���5@�4�>����?�������Z�/����2������5���@��aa�P����`�Zd�wߒ�:}8wW/�3�P����kE�3o��ayMQ��JDL�Pa�o�	6�d#jU��W,�JWTo}��R��������J{j�^bh:��\��(�[MGUmN�R�1{#�&l��v��r_\J��Uk����󻶡^��{���d2A(�^���)%:'բ][⡍ϤNr�V�$gҔL3	`��r/��g�I��M�Ϊ��A6h��Qf�\ñ�Ѐ?�д�Ui*��U!AX4!����+�{� ���d�QT�~B�&Zn�;.PD ��m��QV4{�����ak�HYdb��c�9/Q��Dm�a��\��-U36K��=�Ðn >ލ��JZ✫�,S�Ά��3�Q$Tz��D�$�y�	�������Q�c�V�S������y����#��Oȹ}����ڹPE�sZo/oH>37 ��B�jAd�?��v��85�3���Z�����Kޑ��ZaB�8q�d9��l멈_�QCz�S�W [:Ы]�O�.8}0������串d`=�x�q��oL�=g�� �u;��O�ۗ��5Qf����e�P�3'p�����0o:ѳ\4�J��
�'�H�`�c�W1?���q�h�%3�^u��C
h�$�X*���)����:�����Ni����dY�*��<痺��^_� h�3u�~�.�?Cc��~��P�o��Oh��*6�5��[ʺ���Cƙ�2+�\�6�s(���عW�R~�,�;"�z��V�RX�APc�{�U%�o��/�>~@KS��_R4-���c���2x9�j���Y�h���f�q�jr��B���/�Ի�,�8��_��(8&�}�WL��%����Ϯ�o���N6p&� h���O>�o��}�Iu׿X\�[�t�2�r��:�;��-d1��|/���pQ�ό2K�)@Tɠ ~��Ee��?5��
	ˆh���ӫ� ��d��Pφ��l���W��ڻ	�A�<#���6�׺q-�5�����Z�	Xn���qH�浨K��� 
o�w5-c] �}�J;�F
�bR�N߂3�(y��%�N>(B)�t�~gӹt���S)�%��qU�Rң��+��L�# q���^�{�e�F�/�&Y����qz�A��9�l#]0bIH�k�Rǉ���JVc	^`�єZ�e:����+��A/x���9�T����oE2,��+����5���߀*3�5���̷b�Atl��rKLs���a�&4Y�ıd��}����S������4e
x#O�2Q�7�&���@���/��cA�����k��;.����P���{�LYe.p�W�O:��ž>@��%T�%�;��ӂz��v�aQY�LL���/��Gb 1V�c���t�y��E07aJ�0Ȕ��A_���>����\��j~�;�!���W_m�zm�A0
����"f���ߟ��4�:n�t��xn�{;�+��n|��v�~o����̣��h �)�ar���t�}�5�,�cѭ����\�8���?���:��	M�|�H�~m�E�$ݱ��t�C_D�a�(Ax�G!��(�"��+��>����0�~L�g�u+Z�ed��\���\��	�:7�.T�$'c�U�`��:�ѴU�^-0�,����x��/���k�Ĕ �����;����Sl����m�������c��r��~7}|R�戸ҚA�����U(	g�c���d�R�o3U9y��g)��z��{�_v�g<�2��Rt:O�UF ���������y�v�����T�qq���?]R��W��i������J���餍���a�rɪ[�1]n�YgB��z���y	se�̳��~ ��hE��%c*����-��طM���Ơ_W_�Lw�����a�G�J3{=I`�m4o4�7�w�H���&b, a'��B�?r�'�I��A���PA�\��f���劗��en7q8?4ʒK���?�~ZN�&$�ϫ*S�O�d���gz02���y��ɀ�c=��_�,��@5���~톴鸥:���]����ï�x΅��M�kR`�_�:�BZ�sx��gY�5�7�U�!�*%���ujS�$j�j�f%��ܞ6��w�{�˨P�5c�s.�z�lw󙬰��V���1�S(�F�� ٭�<�-۴ l��M�qb�l��B��U��i�fb��� �+��A��.+�u��zm.lS������-��.�]s�ﭰ�h����L���M̗��=���	�G �_{\�Ѫ���Z�U�C[�Ѕ�l{�\u�x3���]X�aQ,����4Q/�$�x�e�d/��nF������;|^�hC>-w���eb9�f��}�,le���ހ���M���Q%ۅ������()��Jآ�%�/}���$��Dw��Z�Fthߜ*S�c�Q��V�K�p���])�c�� E
��{[�M��˙֛y���=r�NY@<-X��6W��,����E�	^o|��ܓ�5�
����j�`��'��"� ���Z��J)D(�A�*U[e��N1@
����@u?���^;�wD�D<�{7f�ڷ��L�~N1%� :�X3�hv�r��O��ݐ��ݲ[�:���	G��c@��_�ybf����-;�׵����Va-�t���
�A��+�R�������J��w\��H0�<l��� ��I���*�f�"���U�)�|΁f��q��9c��fi��+�,U�*�������� ��=�
�9k��'�q��\�#\z:�>�tZ���P�`���Ӻ���vgt~�u��Z�2hژ�]�G���q�DJ����+O���~���'hBz�$?�+~La���Ok�L�!XpI����#R ~Q�;֡�+�?�e�v�\ewF필+���{�|Ԭ�dB"��m,���@R8"�w�C��>k�H��� ���|�7W.ty}����B��VY��B�,4K	��XQ�`ϕr���U��<��^�k��I�SF&�]����͙��P�ٌ�ȿ��H$��i~�e-U�7T~^-ٲ])�/��^����k^��l�U7��$~]iQР-Q}-�T�N��#@^Y��r�����B��g��L #Z�'nMe 9�W@�3�^�Δ����(cѿ<���F��=Z0�t��`Xf�)D��-����i�m\w��������{a��t��{ƪ�j�$&{Y�<} T��'�X���d��� !�cPf&�d���rXy�6k�V�Si?�������!�Q���<��V�(��V������[�����`�l{c0=!�E�Y�y�ͽ�O�P>+�iUZX���)�|0{�2�cW��_�\F�-k�8���o���`�J��E,��$���%�w�d�`���7���2WL��g����l�kb��8uNK��9;���n�.3�2��*GhH1\u�7��e��1���O�2�B�,�0N��!�y�+3.�v�ش^ڷ�,��q1̉��|�D �/D���(�Fͺ|V'�`���K���>Ma���n��	Pq�L�f�'ő�}�4o�)~ޛ9�,E�'n�F-1ct��DC.��m�	��y����U|�`�Rf��{��ڙO�����I��}p��\�K�Ӊ�@�ފ��r��>a�:|sƶ櫺��ݳ���tA=<���P�*��j�&��P�zw���(װz���!#���Jg`g��[u�F�i��u�<��V�J���  G��c����H��?���=_!GV~�M�g.$5�>�3X��A3����#�
b�0����HpI1��=g��=�zyd c/�����J
qh�L[W�
�4I���.��d��K
;$��F;�r��f���oZƶ�\�QwcTC�䩫,I�jX��H�<��a���ٰc�z���F�p.�Nt2�� ��y8�?~��](�v�G�xܲu���9O��:���w�X%0����}�s��<t�#�Y�=oe'�m����#~��[AL�v��4�3�_�����a�h�b��n�����ꡇ�:�@�d��<�ׅ��m��|W����:�����yMo%\��}�Qq���¡�Rh�倔]�Bw5T��L��}�]�ܶL$�Yt��\�`�N�������炬�B=} �q3
_�4r�5x̠8ϵ|�R���{��jW�LK��ى��#�C�Oo�%�qX�Fv9��4�g�x�"��Y�B�.���5�5���4�sI����bF,yuȈ�٪�$�dp��Qt��<�56²���`Zk��=�bD��	_%��4x����VL�ղ���.�`�=�"�A�q���9��k��C�~�9U�����c�V}�n���cR�t���w'��h��y<�N N���"��67�SU�� �3��$
 9��E�`e)���XJ؀p��sV���r��=�V�A%7�{Z)���ږ�,#���A����)��M��%;2�x�&�o��D;Q��̃3?�-O;{_�=S[��V�����7	C���QC�Q��L�K�Q��vG+���S㴘Ql:�i���R���إ�ۍ�\�5��kI��Z�C���Bov��O�s?�Juuo�v=� -Ǯ�a�ޭh��sΒ��Y�-��~|œk���{�I�ԛ����i� ?&������Я�h�/%Xx��9x���?�ߜ���E�d ��PJavc_L��:Ej�󴂏�׬����u�$�L�W0�'..Q�3�J�:�DIu�U�)��|U,F�Q��|���)n,�֋-�._�u54���Ke�L�M��>�8�l ��QxFl`�UJ�{x�%�(bH���o�l�ټ:�Κ��%l?l��b�֫���a�>��G��?m
c�q�c�7�(�g�haօ!��b���TL�!��N�	�<8&&N���'�wY�Ǽ���<A����Iѥl����] .�W�B�&��W"�[�1c�V�ТR7��se��Lx���Q�op�n�|��]�xi��%�������p��Q�_��B�7�vm���Ik�Dp�)Zx�+�j����G����:�<���t>$�]!gF~-��6�������&8|���t���D�->oѭTM�&����LƧ�����,��ƥb1�0�
ǡ�x2{�.��,�R���(�7\�� j��M����0��hB�J�ȕ𹓱g�c�C	U8jh1 ���X/�hW��(�-?�U��'ǪA�@�c�C��U�<{[�^�YĶ �&����M�����^}I�{��hnp��G��U�2��9,C�I/JH�ǎ]^�,��>C�X`�f���[#S�'Yp��M񍮣�t�%9�-:�;7�F�B��)�OY@�nO���|Q=�|h��=|%�1xd�`B��dmQE���t��=�#�0��=�跱R���8�k�!��Zà����G�����&�
��$EIv+4�k8�Ӈ:��g zK����2�_X���ȯ+�1|>v`�� Z8��p��p^�ǅ�$T�LZ{��awr*���tPx����9�� ��2@w�-	����L�؂�pz_x^I�����ތ�B�=���1�eݍl��1���pĶ;R��W�XëD���{�ʰD��D�2��W�G5m<B�:�R��GǗ��!y'�,j�K1p&�-��$4KJ� ǯ���7�������D�5�_A��	J��U��%��ط�=I�q}��T(�T���*8|�R�|���Z����PU�js���1�T&��ˢ�>-l���2��>���h��#Hb��%B_�i������~_>�<|�4[G�� ?ڐmD?�O4a�ՒW���7��>�Ïz��D�N������������?qn(�AI�tז�f����
��6��qE�� `;��5�3{��G���s������*6�����)����h���6�����m��7��Ih����LH��V�8����<���3�@E�Bn�ʉ�A\ѻ�l�mȸ����Ս�rb��g���^�p�/��
V�O�1��v��|QM��C��fCvX�������$���G�a/{�"��Ae#n��0��ҿ##�ǆfHKx�"Um<��r�;�����ۿ>pI�������W��&m2�"�����&�Hd)���w�1�n�{n5|�"�?�a{Fdh�@�L�Ǣ�p�4"8u�&`u��8~����G�S'����pp8R��b�Io��|;����jLz��^�w�A�k�WDfvN?���`��B�#"R+{�F�l��Rr���4�� {\;y���P�r�%��<��E�
�Ɲ�ݤQ��R��xQ���h��ұ�H�iF���;,���o�����֓�M�a���j�)��^J\d,fE$�:��i�"�!��ƩN��u7:X�a���;������嵩�Ɬ\0m�m���E�Md�Nۄ&ğ�"�'�0����~��m薛8+h7���ۊI73�# 3��gN�.��Ę^��=�J�����\  D���`��G��
U�D9!'��wu���i��M�g�PQC�� l��O	T�=���� �v�s��,\���EcxzL@��Z'��ߨ1js̶�m�V��׻h��T�K�>�)� ��d��<x��� �'Sh$ދ�ȕ�^���⣊;t'��3TF�+#B���!�q<
��p�x���\F}4	�A��=���U���)�̈́ �$�ă�-XFTu�*ׁ�[��"��j��J-�kj�F�2���R{�����֗2j)��=�O��#�䷒@T���h��ޜ4���Q&���\:~y�\��f:�S��vIO�'5��+��Q�Ir0�\O\�W?��%9a��(��r����/�Î���G������\N��O��eD�����2	��!��̇����c�8�9���]��ZBW(.�zd%�}~+C��˛�������i("	 w/��d�j�O�~x�����ͅ���8)�1n ��r��x4�(ÕI1��>�=�6��@&ό�tۿW����;�_�'�:�&o=��C��܍�BB���q� ���97�a�y��� y����9ܗ�.��miY����&NK�B�Nu��2��)2�V�9�W�򰞛�U;¬T;�*��\M�@�K�y����Bw_���*� �<L�$����8q�>&F�t�_ƒ�6���.�8���-C�,�#<:BJ`����a	ӳ�i�л�<�"J�5Ky�)	EYY/�
P"���$�گA[�M?GL��f�����
[J`"e)�-�[��X�S�3�!�+ԯ�,�,!\�萒�M�b������#%8=۔��	�!�p�\}c����t�k�"l��X&��gI}C�z���
K���h�}�Tц��yZ�h����$"7�\̢�ՋE�@�r`�7���L<�NGD��f ��2�D2v��c�[7+��u"��g��ĉb"o�Cڇl�X�|Z�)\/$p�>ɖ��r����t�/z��$!�#6x2D��%�
eRdN����E3e�%P���
n�D�ݐR�Es=i�]K���P�^#�iq�gVRp|\��تϊ�^��N�-<i��{2�0s���������e�&�MB߻J��@8��X�3�=E(���^���-�H6�cפTc�Ù�G�y3��{���.=y��t	r˒�A]��{���T�)��9��́�6�g���	'Ã��B������~�P?F���in���I��������ꘊ�ڡmt)�����9X����A�)�Bbaui��>�+�~�>��<?=� �ٕ��+fෞ͢���V��u�@�{�W��d��-��`^�O��@4_���vW�DÚvb���o�	b4	Z2��n�B�H�.E��ֈ��^�_$9z���6r���<Z����ol��ӫ���Xt�����a�-��m&�;Y=W[ti\����m�Y�j���t� �f}MdҜ�}��W� ��8x����e��rH
e��g<ҍ�������Ni ��1���� e�M�u$�/@�!�z�J�`�ͬ��Va����@�F���^ cC��8VK{��1�Ic�.���;�VI\�LcѿD�32pa�#*	���3ކq��"�ܯ%�X��(�㣨�\/d�����L�r�*��N�U��������a�z3�X��|Ē����B����`t'���J��|���*�r@��J$xy�l��;J�����p�Wn��a)h�f��'���'8%������b������7@�Cy����G@��s��I��ׯ����m�R.�V~#���K�KV�1u{q���E�؈�
҈��)K�8?�Jg8��p��^�1��Ƈ����D�3�퍸5Y�������Lx�$��m�� ��#�WIgG��X}�3|W���G`�F	&���n�}bM.�M���w�QaHpW>0�nYoa$ڙ�v`�Dϸ���)�E�|��"+$�GIB�-�ġ�xސ���pkb��?0��{��if0�d��N��W2�/�G��
���AI����5��bi��!�����qr���~�	��fr���	�e9ˁ~P�h����Q�S�זՕ-�:�#%�S�!�iV�3��" �J��'��L��#�m/; ������i�޳�vCTJo���u(��� �mg�00���实�+ձ%��_�&�r�9�}ɇ@���z+�Gc��_��s�e��/Q��� N[ub`�Z5�/����1p@)��IcN��~��jXj���{`��Ѵ��Qi��:���L��2���
�X9dQ�",�	Zpo��S�/\�W�(�Y����4 �'\���o�~��8�JE�oD���pߺ"X�$$y�ү�<�_�Ѷ�@[\<��Ϛ�\x?�����2ɞ�J9��HM7�I纖�Q:����M�)7�MF<��/%��+�n~��Q4猈ߏ���$:�mm`��.W*C`�.x�(���ը�����!�z�׀59&6в�|f2۸��۬ �t��Љ����`کu*V)ڜ�%B0�F�;EW�^�۞�5��uEB�3\G�7[�}S�)�~/�<�8��Tfvj�L�t��_'�Ȥ�����C�F�dc���/b2�Ӝ�W#�)����ΐ�=1��>GX���m������E�Σ��R�I�}�3mJV�a|�>�c ����ׯ����j��<��D�tr<����b�Z�t^�OTDmʼ��Y�@�YMt��u��,ЉY�u	�p�rmX��#�td���T0!r�.�&	�`]YJ�S�os�ܝ����ls�p�'��1!��<?����[�q��o���5RaFM!��P�s�\�a�����+W�(���P�o1�~��e�Q��j�J�g��gH���1�2�c�ʄ�᣻E,���R{��~4�gߔ��5�bG�#�,D�"C�w1vs�+��V�U�- "H�G����ʅ�NR���Y����a�g,���\X������IcE-�0��kޏ�f�A>�b��:(U��ԗ���D{�"g��r��zꏳ}[���9:���Q)�7,��<7|:�j��ޟC���"H�N_ �v�L��JhZIh!E��Pʕp�K���0T&@��t���0���
�	�)+0�*��M���y�����]��Tסu��:�ބu�]w�����{@�A?�>)�_ƀF�u�S4����p':��i��WD�6��
`������#X�
!2il	�p?��<����
���@�J�O��O��rK�sd��\H)�_�C�F�_Sv��$Q[k`��^�^tA�i�]�����`1�R�#�Nr�<�٧�j���Ǚ@��`,Q�x]-�f��D^��VX s������_�c�7=��1�/٧����C6r��	v�@�f���[�O�S^a"�qL�֊�w]K�k�D���ޅ�-$��Q����Q%�s�����sz9F[��he�I��sX�lb�/��L�y����s�ow-�Nc��y��V&�N�%w�=I�~/D�.7i�$��~I��������W�f���#�����ͦ����46�N�ZN#dJl�ˎ�\'�T!�BTk;l*[�L�5>�*%�*�3)��8���j�ߴ��[���IY��f.����heY�O���Q���g��h7�[�5�B&jf�t�y���c�����Q]���P�<�� ��P�%k�?��r�^�(��e��߿��lV�6ʼ!�tDN��#ٻ�xG���h �����׎��75�AO溫4^�&d�pi~A��K��{{ ��ӠG<n܊��&�&X���͡�%M�������%M���(�l_��,M�(�l!�}�\3��v�S�̭H�y����u�s��
����Z���U]�ʉ���6�%�4�Ck�Á��b��X������9��?�nZ35�=:����x����#y��Qy����)-Dl�b+�6}.L�p��ԈB���G>�w�kO�\R-�_�ȡ�_@��^�W���A���R�i!h/\�=���k��a�'tgV�7�K��%�ƴ^D�V(�y��� 7�C�p��Δ��A�D����k�l�L�[�P��ۃWϐ̮�Y�ȹ�3m��B���	�<�������#���Tϣ�L�]�Y{&��]#�s�B��R.�&�Ґ� :f=M�����x���������k��X����wm�MA��,�U�\��K�Ne���-�,R%�����:�|�s��z�N�=�
�����3����La��
~�	�^me�qZJ��!�t����Ljo<���� .I?�H6X+'z@٭BN�e}�:��5� ��&[�$Mn�=�=4<<@D�C
�[�-	m�8�u)6.�ϟ��;7�#�0\iŴG���<8M� �P�ņ�z�3e9�$�/�Wϝ�v<W���i׌��"��i���������O���}]�VC��f��g�4�~^�<��/��TP�9��t�^{6�%�u����?�����b��<œ���[��g���Z��]6f���^H3aR�7u$�y濼�=�M��P,q��y��r�@@G�-�~�'�Ih�-F�;�ˠ�dT��kv��E�����MI�]O�� [M��)����^n�n���15"�=�:�P�/8���jϣ���w������A�lv�O��ͳ�u�b7D,���q���(�ǳ7��ޖ�!��qt��ԧdM!_��!
����S�_a� �LLE�V��;����C�h�̀�=aS��w��%Q��NK���0i��;3t:Q����Uws��O�b��������y�]�a���:ji&�C�ȕ�(�ƝL����Y��� Ϲ���f��Q(	!v�Q�F�)⹢�?�p��{��~7?Ow6���h�Å�)����V�2{�D*�cɝ#��0�I�@67�*�����:yƌ��$�.�ڠ����Jo~d�A�=�_�=����8ݚ5�O��
/����PL��au�v۞��hb�D�������8�"����K)�,�e*4pU1�?�" *�v�S4U��]|�6SyB��'٥Y/,�{�Nb�0��}�!F)j�(�J���q#���I�˙�U��%�O�(�v�U��L�W���٠�/�U(�PV�F:=gnfD0䉃�3�+�I�~�L�i��F!�8@�]���������}BѪ�_�����z�A]���Ȃ��#����=�!z��N�z��|�V���������D�	�^m�<��4M/�6�� ߥ�٢!��ҞrD�籠����P�_@�ŶC&HD�����CF�2�h6S��
R�
#�e����,}�����c���Y��4�u)$Z����߅�QbgX�M�(~����xT�������S�va��o�X�2�zm0��I���HRH�$k���!XQN��a���<]>q�./�3BJNJ�~B�gp���f��k�J���,�I뿏�/��� ,��N�XY�6��;��Zak�D����ֿDaU|{��i-��~�ԉk�^��D�Z��O��_�Oiu$L���q�=�Ib�ã��c[Gq�>��j^n}��U�gU��̟A�>�����[����l]P�������H,@ț$i4���˛W����I���0F���D�m��N�:E����w�]}y[���e���6�\��{ �b6�;��ě�a6����@�����D��py�`�患���$���pĶ#M6���/ȟ݋9�sE�*��KZ}Y_Qu,R�?��Z����zTy(�9/�p�C�͒Ֆ���� 7����F�3���G��P=B�J`	7��*�1XۤB$~/:�+�;D�X�z�jwaNM�̽भ�y@+��9>�I��H����;>+���c<G�c�y�,4��g�q�!����4�0���:�����P����iK�qu�r>9���4@���yR(=e"ڪL`V@ݾfe��X�!�o�ކ,����vC�����2�����Ů�C�;4mp�.�w��ʄ��]X����Y嬵�x���V���G��r�l��%*�6Y�*��+���/�p�� ���D,���Z��LU���=uň�eZ�ُ�%adc>���EK��*���{��S����>��.Q\�V��L$Atm	4��R5ߜ5�ājo� G%k���a�}���.��f�tvd�d�X��Ed�,��E}YpJs�%�!Y[�#�@ճ:a��b�JxЕ���o�ڦ�[���	t�׶;�3#� 0��:D��I#�:�p(��Ȍh�U�>'H��V� �zl�{:���V��3�O�V9���Ði�rǻ��Ź�0�-������s�j��Ħ�'̺���@����Sm̱8���+�Hxk��Υ�k�oX�obo-k#2��ẗ�)�
}��.�T�b��bw�Ŷf�[��Պ�Xh4�KS�d���5�"y�vv5 o��zk]D���qGs��P��{~lMD��@�`��9C�>��	��m5��$F׾Y���c(���A���=(��F1��U�5��
U�����~~K��g�1E�}�"
{����s�Z��q����
�҆�D�찱�FO�~9��=�\��i���K�ǌi���ڈ�^��]s�;�wy�=4���8����f�?�4�	�y	�	*HqR���p������`V�E�9jpI�be��[�,�������vF�����p���Vu#J�?̾S�R��8g���F�T�h&�:����e@�@}�>�C��6rq�.|, �?V�8�_'�Ĕ�C�ӀR+y�)��Ta��3����޿����R�]�i�CD+6 ����V</}:0�$������m4�TQ7�X�o����0~�òţ��Ċ��J�Ĕn4K=ݧ�a㜇t���Nh�o���C`�]Iy�G�t�)��n��@vf���� ^�ly3c-��n.�c�(>�]13f"��y�X�ǡRp�F�\bi[v�� .�z�"��nY�E&=E�h��â�j��+�������?g¾����:�1�W�r�����"g�
%��!ҥ��p��w��˹��.D�eC*	ۤ�P�Jk� �Dm�����=G�J�~���v].���9�����l�$&oD\|�ک+��'̫M�F�����ߕz��N"�ߖ	��4�Tn�zE}r��ab"�Ʋ�.-D7�N3%�8��R!�N��[��ՠ�Z���\�˖��f0�H��`�k��a̬�RB�=S��,{~�J��^��8_:@�ʅ���
��9*�@��_M�(��ćىl�0<v-��������7��`d{@�h��cj�n�W`m,�0\����1����Y�{��+���-b9�t7��J��%ˮ	R� �n�sN}��eKM�����g�6`|�(h[s��7w�sV1��>~�)QR��@�߰=�L�ՃѬo����Z ���ْqJi�IQ;��bxK�;��Z�F�IBT���?8R���򨈲,ݹ��w�]�����|y�=����̀��e㕲��?������9D�<L8v5�m���4���,�Cޡ�{�nmǄ�cȝG'$ܡ�uď���6�-�.]�!��lҤ���8�%�{@�挻�d�3R��⣻��@��m� �z�Wߡ:9���rnx5
[�����jXf�rl�+�V³��5��+���z�vuBN@��}�}�%�ےȃjkg��a�A���(�\�
�u�L��X�S��8R1w!�}���(/�E�p7λ�U��e�8����8O>���du������>�f�U0Zm#g��8�a^�N���������׮���(�0{tK�9 >.���bc큅�Yiق�DZT�*��b�u�Ը�;k�Y �Jݹ�rʘ��X1v.��O���Q0�
�,JB̮C�+����!�@�c�1�M9{�͎_v�3G�2�	B�m3Y��C�w�BH�xW�X�������ܸB[1�h�פ5O�u*���ZA�n��a��:ġ�\t\&F���#�<�g�fgɖN{<��dz?%�����<�7o�1L�f*ҪV�;��x��I�_�_����E����O�K���i��[=fJ�n74�c��^s]�b�Y�S!D#v��u��'���6���˩��G�"�8�@���	�5���aI����k9<_4�/)�,CT�o�ᄳ�㾖�mS�.���>�)2�.(�����[�/Je4ϔCN|�l}(;}����:F���G�k����>�,��5�3��l�nm �ɨ��;�"�.��V۽h����r�6��^�mݻ�l\?���}�����!�_F��LzOB*��[�^Z� ����\���ܜ��s\l�%D-ʪ%d?�R�O��O�{a�Tc9t�(�FN�ɻ���6��%F�`�A�T�)��m�����o���̬4�Un�	,�]��=ﲝKi��hE��W��d�l�w�y^��g�6Q�n�Ť��6���DG��ɥ@L][�cOAͻ�Wv=͙ퟌ�ha�m-��r��
���D�����>�Y��@��E����v�^x��,��GP���O	�|{�H�-vT�����?���"�?�Ըz�xHw���>��)��+�S���>�$��� >m�=W0���l��wT�8B؇��&��:�̓�-�m-�R�LN�+R�j���|JXq�ycg�z�����F7&�L)b_R��Cl��jF��9xJ���*{���
�JZV,�o'�ɰ8�cF��z�9��ݛ򑐲�� 2ᗤ��Mu�Ah��prG����C�:���5��Lj�7�9��[���w�n�P�P���O�W���ڗ�̨��'��p���2���^�����
�$�\���ïB��`��{{���O���Y�^�#0�R�:��$$J*��U�	����HB�H�����'@4�"��_�y��������Nlmj�h=KĬ�5!��o^�
��k~�ЭA��g"q-T�Bq��M��;�Nm����)�%�iLi\B��x
.>c��[�+c����Id����ً4��Pj^u�~��J�j��K�B�6�'x[���n�'`�O�$�`�:�������~r��<����V�G��'��-�ޜ^�a�P!}{	*���ˮϪz='�~_-��UA\�>�z�ƨ9'�'�q��W��V*c\�w���WL��g)͠SKF�U��Ĉ�N##Ŝ���_Q�Axq��w��@�8������J�'��î�	N��֐�~���售�u$$�MI����f���0�
܈��6�d��k��V�Ɔ��v%�Ө�<j�,iG�Е,��C���;�[�Eո�D���F��+�Px��k���z�I�Ei,0������<�*o��%D��?ߐ��zM�hz]�e݋l��X��]^8a�%yC�7 �Ӿ7����h��;_����� O>	�n�!s�/*�(19ᱽ�z��J,�S�����z��!�z�<�6�`�i[8V
��R��#ll�%���8�ѩ���d{��-\��������H�"��ߧ!'Cz�W�=ґ���f��}1i�TsWT��3M�:x�`�qg�Բ:w�j�R�r0��ӛ�L���6\2�&/4��f?J�� ��4�����*M(F+	�Zbs����1:��D��Ou����\�"��a���5�L$1V�PrR��*=>+J9��$�� 5}&B��C�Q�?���'ό���B�m"�iM���u\ұhh|f>ֶ_o��h
,��q���F��A,���]���_� �8��G�A���Hn�!�Q���Ie~��:Ő�Sz���=�S�TPo�+�Q?�g^)ʇ8�s�V�B&f���sQԎP�n��7����*X5�_��_�W-��@�N�'���|�+�7���
�I7���rO��n�v�~NA�B�c�>-���N�,�ьN�y?m�1�`�mh`m��	�+� ���G���A?Z"���*
7���_�(b;��a+����t���,�J'�yQ8Gm�J+�`}�肟�(;�>�Y$A��X�?��^���];�nSr� ���g�*,M�S���ze��9j����-#��I������҆!I��`i	�(F�B�D��Yj�p^��$�g��7���A��AA�0���m[5m~�ی"��`n��x�9J���t0$U�k�=�M_tɟ�ķ�F$U*�`g��H(�e���6v�^J*w�9C���"N7�F���[�}�B���c�_K���&Q�D\���U0�����(��mv�h�F���0��\& ����l�1CPO}�E�x��1�
�QBu�� ���a�e"����j�;��><
>dc_#���ދ!(R�G 2ߢ�u7a�x��VY`��nY�*1i��K7gc�nfнN _7�j8[����J}YM�0a�	��ā܍>�*���!\�hN$��)L	_���j�+]����#��R�@� �v`�E���qew�Y��#�-�Obʁ봫����&��d�6L�@H����8�z�f�K8R7��I�t��L�)��s��x����T��I7*x���?tlý,�y2�O-��:�_�S����(����C(Gp�p�s�g�7[G%�;+�{x���+��j�C��K�����;�
D�I�g�Gcu�*�?�cx�?�w .0*����%�I|p����&9s{�]	q}�D��ք��F[&$20��aLZs�R�na\Ok ML�ST�c�z�MsN/�tO}f �O�v5�ޮCMw��M���tጯ���=� ����q�oB�͸ $�_ͷ�#��	�ZmO�'\5���P
�����C@Nh�ԫ�i�ns��[KtN�O�D]��޿n�I����M���7Lk�6d��V��11�L_#����Ȼﲰ�U��<�3uS)Bntj� _��6��Jt��4&��s/j�hۀ_(b���f�Oy	����m���w�����,sd&��7��D��םI�	ţ���'LH�}P��R.JpB��uk?�C��D$?�ݔ�2��U_J�kbk��ü�b���e�O�E�� .����ل�wlxt�Dl$h5R`*�(t
��V:l Ɛ�4_h|���ÅZ6��̳?/�6D�>qO��D��D��J;��2T�<j{ggW#�E��qs�0�w�[�bܓV�iZsV���0�3��eLޏ@�=@����0?�Gk��=�ϸ"�-0,�X��-�[W ��6ն�yS>\��P��.w�'Z��e�W�����M��ތ�TP~H�����m��>ն_�����A]��U�������������E$�X]]G��2"\�hԞ��|*n%S.�0J3RW�2���EJK_��B�U%�}�t�z�Y�he��('�Ǿj�ԥz��h�AU=+�q���)����"-�l���>w*��;s����2�Ή�&U��Yj�P�e�>��e��ϓ��& ��h������F�mҪ������g�r�\�DW��z��wQ\`���s�P+�H������pr��weɁ/�����ʉ[nF|�}�|�+�����{z�A�� 5 0fWf\�l">	���G�w�>9|�դMW1��-\��xf�U���/M���yHl�vm���R�o4������L�����r�(����K�׽&��W_l�p�S�UY�UD%�8�a�NkQ�Q�Ӫ}�bk����F
�&��������*�xn$�_�=W�M��y�]CW�҆Ax����IcIN|��l2�gE���lpk���;kP��+�t�:*��@7�i7a!`>)��਎�q��?�M���',��蒎�Z��J��N�p*rޞ�1��P�]0{@���G�.L6��M�CW��(�)�����Yx^|s�+��0�Api�;�ǚ6$�P�)@ʺ+�u�g<���,�AٙV�*=6���%6�M] ٞ���	�M���v肋����Mb�U,�biva��>B�7X�����cS���ZQ�/�wA+k��p�-�oK��ȈkE����>��'h���;�4L�X��G� 1�yʈ�(�z������r�YҊ��ֵ�G��#�>�Z��l` ���C�$ܰ�y�jg��ߥpeRN��O���6Q
X&~�h���ŷ�3�:��uk�j���}�A��m�PO}�,�µ_�>Ҟ�A��
�a�-ͽ���g(T�p��@oE\�8^�}b�'^��1����h8��C��"A�.T'�����p?i���پ�4�r%4@ׯz4N�ܽD����y���8d9n��VWv1>~dBf"���WK9��RJG��:v[��-�X5 �(�v2�kr��Ϊ��h180�������^��f:�7#c�=x�*����	:��2���&B���I3�2�&�LB���/�J�ҿq9u�,<�M~�a��=����<Di�Ud|���(�fM����*�~p����k�i� ���
�hcx��٣7ަ8%��tk�q%Np���u����'N���Йyq ])��;�O&%��ѝ]���4���%���%��0��s�]���]K�Pksl��{g� j�ʒx����7��@ؾ��qř��l�h����0m R��q�Æ]����v=�����Ql��ކ����
�\p�p�Kn��i�M}�oڪ���!V�Z��� ���7�eA=x9o&�U���>�D�!6T�J�3�E��Q�����ޔ^��@k3u�N�p��a2�Z^Y:����ؚ3L���(����"+���u�^rJ��A����MQ��T�e�d��Ӳ�Y�Uu-]���WE�g��/dL�� r��C�:fT���q[j��1]����za�c����{���oJ:h@2lz��f�?3� ߶�6�����P����3�ː�W���AL0��S����]���8���@�8C�ds�Q�ز�+��Y������>~�!�s!Sp�d�f7M��I�ޢ��D�	�ΐ����Q5�q�X�8"q��C�~"e;q��� ~�����v��-�����E cʄlXT ��
��$ yl(r(g&b?����0l���~R[(޴�~{�Ɗ�P��ʢ�(� �x��gA�8}G���WkF)�~��;{Ȇ;����O�1�����4��(�
�����P�\R��=�8p̧�x����**8sX�ˊ�q��NRb8�q߸>��@�;̙�!+J�.�>�nrM��ǥ��7��޸S����_H|A��H�;Q����E��Ԣ8��һT�^���iH���5vև�XV%�v���Z�W�&�M�ԨC�t?�P�����%P���@���BIM�(��������ı�
"�,����N!�]�;���>�'��'���(1�j�mXw����B�����T�腞h
L����6Tcp�$a�7a=T�(2��!�R
�-V*'�N(����7��1�+���-ƫ�!�1�n�|٥�yHBڰ.��L\%������^�(lM����l�����{8P��Vu(�2���DxaK�Rj7���7�@Ch��8���W�UX��M�3T��3�M��IT��x����+�"d�1OVL1JN�:�3��͠`����%��3S:�	�`�N�'����~��؁9?�Q�(�]ۓW�VA��!�]|<`��t@�,�T�К�7R���d���9d���E�,����I�AO�:/����U��ui���n���[�SmbR8�f"����Q	\���fk���.�������V��i �$H�����R��u#�q��.���(�������>_#4X�O:g؛o@]|�����.���%b���
v�EHm�>A
,4$ �"�PqY2I�@En�?���l7��11oŧG�N���K��S�N��M�l ������Xb(���,0*�`臌2n��e�X�,Yp���4R���>����ubWf/̣�l�H���0ǯ�q��3���P�j���G�4���B��&�v���xW�^��(�M&[Mn؟��%o�����)!�Uw.%���H�c�f]��7�j��p�3kQ1Z m��8�`��!Z��hC(�E����p���rXI�p�8���~&��bӳ��� `�{���dT��\�@pxU��w֠��r;Q#$�;v&�y�@.���z��b<)��?��ԨG��d�k*R �2�{8k��P_k��$��?ƭͥU�������!6��(D�\�/{Zk�RS��&>3"�7� i��0�2O�,K�P�[$bQ;/�&Z%Bs�����[K�
�x�V�1�"LI�S�V'+�(�嘌������/��&�i�ǎy����	:ݚ����f\~i��i�R>�67b�4l0��Q-�_d��Y���=Z�(פֿTF���k���]�;?-��r�w9���Bn��;�c��h��T����-EX���P���U�Yi���Gi��k��`ڨD�I�)MV�gV�c�3ұF�f!	u둄��������9���?O��[O�Z̹���k<N�@���i�y�}���D����䘉wyv0v0 *���P�T�>���I�a������u.��\UŸiff.�C�5_^��О�Hg�N��9�E�M��� �
�zaۮ�o$��h����������A�֥��	�udڣ]����~s�w�i/�`P%h���yO��;ӹ[N�$W'��8��(ڢB��	�M�*Еe��lMҲr�[�{����F'� �â/3�~��r��ii<<��<��&&�¢l��~���T���q^	 �C�q��a3�D
����~y9�0!J��Di��k�"��7��89�5�)n���������s?��*B�R센5��8ꊝ����>_��h"з���+�Z��Ҡ��#���_L�I��Z�L*,m�(���l�v���3H�����L�7v��vSL($*���0�Z�����H��#+��R���E`����J�9��V
F~��9�2��Ծvb �A�a*!�Zbٞ��]��y��{B�&eB�?T���w0i�Hu}ʀHE#~���O��������
U@�#�	����ߡu�ɑn0OV���f�y�ןX��L�!�5�qsM�+A��N�N-����]�ڸ�P"���C�S�ep��hP��P]r�O�i�Ȥ#â�r��x��<]��h����ۏՁPa7י�&&���(ż6��;3[�]TPi�\�֒���s��t�I!���;҅��M���w�J�pp���6�f^u^��}��[�u?�&D~�U�S��m� ���g�,y�+�!�*�s9�*��2��a)ܵ��P�O���+�:Vh�2�d �����2N�>�	�}º�Wi�Ч�t�lm��F�)�ݮ]�>��,���\Si�Z��*[�	��/�TɆl�le.� �d�H�bS�k���T�%��5�N�d*�T??砲A�:t�jxUD9�IBޚ��5@�X�tf�lX0��/	��Kҹ�	�u��d?m;ߑ�5��F�BNymY�����cb}
�BHt�|���7K(�R�z�Wןt6������=��Go�-��bE�'��W�ZRv�Է��kM����o��A"$(�5�i��Xonp>`�9���KF���㋘�,��2t5=��ν7�SiP�0gI����z{[��HŃ:������ud\���5�=��{}=�渝Cp
i��T΃*"|�j0�FO�;7����J�l���2�A��<���?�r-���g�O�S�nu~��o���P&�b����"��Y͌K��!�-:�r�]%��#md#\
�((�<񓆟�$��nrg(�{ *g�(���fd��ɮ+�sX�vRK����Y�(��H�v�s-+���F�I�i�TR��A5���8��վf�ߢ;�nT�l��H{�������&��8���D3��qYY�Y�������#�"M��u��I{WJ�M;NH�ؿ���S�	<�tG(��3���e�kĲb�GKk��R�h�30�MH�^�>3x�/ىs'�
\{~��S���������Ӧ�? ���K6� �xN��a�œ���ɕ?PuNm���zS�w�N����� ^��O�H��8K3�
����u�hO�6�z�=�"3�y��SO�Q�1R����X��0�����ZI�Ѓ�cIK��L�z�����ԡM��?���e��-A��O��Nrw�91�k�H<��	4XS��|7)ӛT��H|D�8�bM�l3(�;w8�		���fn�n��H��*|M9O;弬<��b���	��U�U��IVZ7��X��G��18 ��>xG�>E���`�]��vא=���8�n�=�յx���ْ�8!��b�TK� �h�:�t+��e��cA{r�$�Ws�Xǜg�0//��0Nݣ� �K�+̪'jTDw!���(�j�p��1$䣮��QJ �)���������D#��뚱ȵD��rl<��N5|+��#0s�W��[�W�^��к#d����p�S�L��6M.�L�p@\/�"����KDA0��x�:DI����o������W��1Vs�ͮ����x���tHQHf-:���d����w��P`PJ`���7�v�	�u��]�R�5�<>�N��y�>;p���f2L���	�)阆�τ�I�:��d���d��
�c��P��7�/Y>��5��ֿ+��6�8=��"/J� 3�=w�P埖�I�?��j(���>�����;L�H�v!��ga���@�Sw����5�C�0�k@u���@�if;s���@k�rU(2�$�Og���1�f=ٟ*��ike�:����8Ls�a:�x�0҂�k�J��;
���e�%�U��є�i�X�G0��P$]����cČט��i#��rw8	�;��?�ӵC��;��@�]۸��l8(�g���h��]��|�o��m�w故���'�) 9�
{@k�]@��D����>�B/�ZΔ�K=t��_��˂�B�N����`���� �xƪ~��f^����'��x(+}�TP�yZ��\��l~�4�`�6^w���K�ci�,w/QDգG�u;�X�/���C�&qwx�<��Cn�~%N`;ph.��e�I�͌�RF�/K��R�¡_/��"��
�iˏƍӈn�;�F��>?'�)J&��M���+�#�I͹�!>j��yX�7����o�O�0�F]�½?�w5/�j�.8�e�E�2<#��]�⥁b*�,'Za����<�~!�k���{�1��I����jF�>I�{��OK�W��h�S�p�-
�I��v��Z%jF�BE��!�P��闵��h��U�)j��ew�A���9I��3���B]n�t��4�N��Q�_�JPo�)�S����;)!k�L���Q��� ������h�m���q~m;��¾v�Z������j�3趏�:����b	�~/i9�@x�>}�X�á
����]t~�s�m{V�.Q��|������'6�^�^@Pq�*1h���St��x�8k���^R�I���U�K��_����������ާF�8�4���l�4�R����]f�H��~{V V>�~��ѡ���X7�	�mUNk�[��hhj�28��*~�ߡS���I��X�9%6-��>������E:P��B��d�r�X
�)X�-����j�Y2!�]��=!�����WJ��U�!���"4q�<�H*�t!4���ס�Hf�w��۽\���(�@��#T8lO�U���E}�p��[�q����J��z�4s�7|�&�[*��;�"��J�"��Y($�2jekڛt�3�i�����I�?K:v/��X��C�n<C�sS<��8��i'�;���R�_~U�zɩI��8(�<���[4�@��3e@wZ)�Y�)��X�I�wN����z�"�S{9x��E
��C�~!h�Y�u�2z�(�9W�-���|W�R� ����D�����r�K����� =j�xo�VN�یt?�K����A��C��q��upj5  �����Gh�;fq�^0u�h�|n��a�/*lJk6Z"m*�j�� �7����j�����y�����^�@�o� 
oX�N{�Na7" �:@�i�{4y���)̧pmaMx*X� X �'$2���cP�[�GX��77_-ç|�U����=��ŖӢ��H�Q���`�~R1����#���b���T��;o��&�,S��ն��ߩP�M�_KCJ���C[��$��;c ߰{�{*
h�J~�W��N��"����Nk� 
�l�$�В�k�'��M�P;M��w�����0�6S��6�*)��l��7���>��s�dG>�i,������~X��_sB�P��k�/�h\f��6���ϳ���
Кv��>D�핢�U���,���i�ul{�|�5L\h��Ζz4>�E� ���6��F�!>X���� �"g��Q�|/C�G���}}URz�m#���_E��W֪�  ��/zA���g�+!��p�r����Ih� �[7h��0�Нp?��6���8��k���<�������o�y���:E� ��)]���a4 -�|<���<�{�l���Ge��c'��b�E�[]iG����Y����D"� :,������RH_��
�=C;=q��=pe���7���&��7y�J"�TM��r��21֋�S�~+����Ꝅ��F���s�E46�H�ĩ�bһ}h��BKe�W^���X2�B�P�V��O}�"���<��0L�xI࢖���eX���l��M�W��旞K�>'j���D�|TC%I�tC�JE�ly�. ^��Lk�6��+�M��*��-��3�H���6֋m�t9_9z��5<�3�����鶖JOD�9��$؄S3�Ď�7}�3E9�f���vF�=������ٯ{�چ�´ƃU�R/0�v{��O�K������ܳ�c�My������E���+L��6�͒��u�ɑo]�u�f|;}%�۞��wPH���t}_����&e7�%��cu�U�Tg0]�RR yF��~{K���=��!��O�L��4!ҭ3����rJ!����y~�e�&����<��3ps�8�}��\@	���X2���=e�����"g%hw�Ŏ��$�*�2z榿��]�Ƽ.s߃ɦEx�+��R�.a�aܾ��"0(lY��|�)�,�#����.|�(�D�cG{W�b�j���n[(�{�섬U���x�W��J��)�k�%$/�{�/x���7(��9H{5�I�,����j#�͙:�^t+YG FQ�~��v=)���$#�}G�QA �*��p�A4�@����O7[0=�s'��Q���d�M���)҃��wI��q���{Gw[v0��{\��{�8/L^�m*K�����p"bCi�ɲ ߚ�儈���9�|�����X��ү7��I��PF��`e$x�n��8�Qd��Gn���\T�~	�g�H�!��<1e���;��`s��c�gȯ����X5K���:l�����ѠǓ�=Ҷ�`8b�NM ���J������"�6�w�M�Q���a�f)����lN2�.�wJ���l�����F�d�;�����cJ7����J���P�s�1�JH�Oȡq������FG=���^Mr����r��)Y38�����>&Mh�;Zv"�M��7f ���`�>��؟�����~_Do�+�E�]dݼy%.A4�1� ��iO �ݫX��kK&�r�{1�J-��*!KĦ�&��s�U�,MΉ@r�/�w���D�~���L��?�"]%}M�Lÿ?��	�5���yr��S���`yaZ�b�N-��J�^�#7����W����>�daxi��2�H�[V�iw�Ru�����uI�|����AMI�R��k�����%eJHA󵞮�E0VZ#���� �o�:�F3�$(�K���Gg�MpR$�RLc|����Џ�6*$�;�0�LH�����4���E!~^�x��1UjH���+��\=}��rYj^���^�Y�oU�o"ǳe�f�9ڞe�c��8I�$�a����\z��$=�ޗ#�,�Bf����mZ.q��JW�b���~h��Ԝ��қj�EWvP��O���_��D�"�/,�����������Gߨ��n_RH�+��������)�}�`n<h�C�CQ��k67���,��C-	�#��A�BC�3uFBb�˨�Ē�X-�?EYhiM����Ǜ��ӓ�@��"�[�:���Lt�b%�I�]tN�����	j�BskYT�DIi��E��&n)���T�W���.o�,������s�;_��o�;��$�|��%���χo*�uu�<"����(�>��m?]��u� ����S7�7�G���D?�s0��5��*ZH�G�Ωd���e��@*�jGؒ^4;���uFs�hS��:�!�q�W	��X����DX?��뙮ry{T��=Zi���u}�|���m��&jY�}c����yba�&������R�Q}�ghp%�2C��,CB���!T�c�n���"�C�
�D��gb��U��S�	�����W�Q����޾�W���ݺuoP���|���{]l�w�@B��s�wjFG�a�U�s�g��L�� ��#�wN ����i^�(�u_���ז�J�1�cg��U���5�V�?��5M8i=�N)Vȼx�����wRm70��y�yB#=�h�gLGG�����7i���#|p�n�L��I�E�L)������PP�󛼶�8J�V�ѻ��T���a����`���I�E#�Y�g�z�~H�(i�_�S�iB��6dz/M�����B�fK�����ms����MZ��$�č�w3i�����0���,�@Ɉ�M A�W�3�IE����x���)��6�΃шIܷ'&"pl�Yt��B���Lcc+��6#��M�:�����5����6��@��F�I�O�%�M�"��d�rO���eҧA��u�Qrp��Gr�l�ҹז�\���G5�HV��qa�(�~���<���Ş�b28��s}�㆖���i1uQ�v���+�suG��|~��͵��!�����A�sE0!��e����n7� \�3�
�o���ߚg�13vAV*�^������@�ă4�Ҩ�+�kU��ٔ& �<��d$HЮ�[�a���D�:ȲƬ�36�cLu��b�ަ��I��h/"��rUd�%L�����%���j��a��b�M^�G:M�Xʻ�B��bΰ�5�g��c�@�;:.&������K�-w���b��o�z�wSpܫ�Ra��aǭ���:q=�B;]�Hjؤ��F�?���(��|21�Ζ��y։�N��N
�i
�����Kw�Ȋ�NTX�>+�'X� ��D|�k�ɏ��	j_���VvqWq���A�����I�͜TPPm.afpx����č�e�F��ے]I�ϕD�$vJ1��q�
&�UD��/7��*9^�o#�A��D9:���E���ċ��'���$�8��cI�2Y\�_F1�������kx5C�V��"cdW��<�&�1�!O]i^�3}��8����l�:<͖��4�����w��З�޾G���L�����U��b=�ݵX����4�� oc���U�'n�L�I�;m�΍��>�ŉ�ʵ�5w@"#6z��d�������g��5�^W�j&j��eu�=,uA��	P��i���r!��<�r��w�xGk#��4?�l���]p�f���	>(P��R�Lc�Whe�E�������>8j9���]���Ļt�t;���pRTBaT�c�)���)�;�$I���M�-�����@�p�a�-Ĵ݊�uL~$���V�~��������X�	�V�SU�h�^�{4�p�J��4�~\\`1r�/���:��A"�K΍��D
�N���KfA��U��o��'qu窄��,v! iI9t���ᗛm�7x���~�7��
����8�e�����Zסb$G��(�w�~�~�+�y��xm]f^�����q-*�W&zkgI��NT-�Ok�f�U?���{UQ�*���_r%�����κ�e&�k+A���~_��d@�kq���<�e�kgݧY�u)� ���1^��l�>�qIkϓЭc����b��I!V.9��}^݁x�S]��w��)��Q�}vͪQGD'b��0��l�	�  P]7�v����R#K;�#�i `��#�ZRIڸ�޺:���ϓ��7^_H|�ɞ=VMk��d�}$k6���(T[{@���(\9-"�{V�Vl��i�ا�ofL�߬��"Y~�;�T�z󁡊A{FD��ٝI��j��3+!y�4f���
AB�>��&ݴ'7�<�Y����1�<� D�Z�Q)sJ�L��f�'�#T�X0���J�Z��h�����7��oxԆ�z޶���y�!E\Y��֩��0a���[3�i�Ϭ��iWڗ|O��p�/�������޲�V�Oui%��?��9܍p�3x�����t�A#na˸�8��*�ug3��I�KA�5��A����Sτr2���94pI�:ծ��S�!-7ϳ)\���ek��K���N9�yw�&�j2����	��=wh�#+�]͚�+�>5���/*a܎���f~� �.`��G�F����6�jOPnSNK�w*|u<U����*����7��W'��Fs��욄�1���RЃ�����	�{��#0�a��^ʵ4�^�v��/�{d��y��PN3������2dۘ�/��'o��iW#]e�oIh�l���r�I�c�$��]}_�Xk����T������#䌵y}ӓQǻ4����k�k��p;9j]P�v��Zn��7��V)� @G��[1��7�k�{� ��S��\	��zַÁKc W������RzXw����OF_$@�3���]�����u䋭:lq�ГS@��7�ٞ���U�g}^�φ\\�$p�$��?|�R� %Kva��q~ɥ7�{�0pE����P�g%Z$6rnz�ި�sڣB�h��Y��[�z�АʑȎ����M��`�����b��Q��f���ieZ"��m�i0�e����"�{�$+�;\�3w���6��:�z�(��5�^H�����ŮˑN�����k��Ƥ5��#ݒ<�M��G�@`��l�fk|��m��M٫vԕG5�_��_!��I\,�-�#����R��Qb��dCrXf̘:fSS��g{F�����*ȓ�}""��4�!�y�B�_(;�.e��b�DV��M�t��O;_�_�S�i`W�8B`#g�7�Y'r�ˎ���ׅ�jI�?���v��T�t�g����B�l�����PX��Iw{s6b�ߪ�^m���%Z��a����S���L����l��#��ƫ���*��_���Z�y�N�/��m���X��J�Y�\r�C�+oP��8���p*^�W�
��!��,
��}�B�@�cr�̮q~���x���'<��@0�J����M�L&��@6�<,��;@ӵո�l�#����,���U^>���'�M�~�-��y�[��/<����S����U�V	1=-�l���=��nm��&�bҏ�U�����jC�e��x���'O��hֻ�6huh;�h2RJ�}`�3���"���ąa]��E�GjVy6�P5P����J�;�w>�l�r��p*�H��2��:X���EQ-��,ѷH����,�R�`,��̛���yF)��8��n,�S~�py�hx�M4���.̺aϬ�D����/f�x�s��J}�Fv��@��fX+B���}�����,nbI�B:p3#X���<��k X�(�	�o�ʶu����~�
~(;ꩁ���,-�|�{}HЫlт�_4��#'�#�M��������L./�����:�r���Bb��-,�#�DV�L=(����́C�tf�*��l��>W璙��m
O2~|�,�o������O9X��~��z��q�p����-�f�&p|�����o�m$u��T/��~�]�S	�������Rg��%]f�
��)*X>]��f�U�{���햷;�j� Х�B��t��L>�w��L�{��ۙyY���`Zm'�z����ZT��b��һƆ2y�ys*
��HS�+�M�.!qn��
����OLXAk[\��eU�~�X�v�?ZA��� �z7�v��y�B�£NsΥ��O^ {�+�w0��=ܱJ�n�.~�b'AY �ui� �j���jF�g��)�qy||�I�BpMN��H�����pZ��}�Y�ș��ĝ^Ym���
5�O�eBj�� �?�HIl^ �6�ͱ玨p��nbt�f���S}��]���C�'4�/ȹ7�Q~��cF�A�bo��%��i���t4H,�A:B�싔@�S�-~$]��惌<����n�Q��]m�9�������}��kBB�o��ksSy5�.���;ҝ��nɕWf
Q˵���A�8g���U+uF<>����t]m�%��wd�^es$���Ykߓ�;�\&���yg5N�`f�-d����ނ�'㙺If�ۭ騼��_�&f�	�a@3�q��T�������b���ց�3&1`s�����P��6l����4S����R��"�ϋ2�VD�4L�?���Tg�R�äT8�q���?%#���ǟ��4�J�LKgL1�I���y+(3OWX%e�����%��#�k�e�ᆈ�Y%_-+�i�����q6?��s15��n��h�q1�����Oa^�,��%���+e;a��.�q�(bR+9�7�r[�qZ�wa|F�5�q�gs�0��\��G���|��n�����u��|H��ZGg�/�`�MD᛹�v5�!o��%���E I�&����K�Y�]Ƶ	)-֟������� �.�����ǔ�h\�sw�a9���1��t������؉A�������J��2���� a{��8��
����cN���X�G����{N�S`���t�����Roj����=դ���s�e}T8�m��j�8�I�.]�*,N`Hjo?��Unwd�j�-���]��Ҝ��K@Vl���-�/E�c_"v����	h�w�\'�^��y3Ln!�m��?&�fkru�;�`Y8@ �0X6��Å)��g�D�������;�`��A�ޏq���	���j�||��C����ᜀpa��9Ճ%eD5���(���,4���n��y��V�pT �7<'�Dm��oP��Lz�9��b]�q����:�G㔩�����'��)�㧂�<1|g�ȋQ���4>��c� �����nsF���`؆��[⯀Fk���sז�����p���,���)�E?�a�W��X��y����7ﰌ>��f8.�¾q����0�M�t�|9���W��S��w^�1�'ᣯ�o�l��a�gիe��r����e�u%w��@12��҃��[��}1�=�{ޖs9Y���귅��%�S�;�8�?��).S��
^���}��CM��^�EB����7�
_���Y�Km�d?�!L����+/�	���$�$G[�� �N�+�+���Y��Tϕ�[�B�K�U2q�\�]H:K��~sV��U}�����_6b:�[ۦ�	-�Oqh���S�Ag�ֽY��q�x��5@��:ha<j��E�V���o�.�1&�
���XBy?�65�8�y ���$�1�`Dr�ĎM�o�>��N���7��/�;�
��ow3��Z�ݪ)I2���w�Nݖ'ԯ�$�,��J�j�����د;LKE�~�����u) I0��B����ۑ�5���X�;J�V�ў�U��A��zN	��ά+�$%\U��-����@�2��~!м�N/��M9=��@O���+l3:�����SFn��yο�����)���z��h2X4�`*V��(䍊@��b����L�5G]�l�[x�M���MWI���o��sh�d���A���p��&V4�B(�J�Bq��H�ܸ��� �wf&�L���� ���i��8T�n�Qw��T}i���QV��3Ы}���>���kc��>�}_��/&`�?�������{t�A��y��BY#[����O;w�F��t�cl��kT�u|r%�u�QT�(� 8۫���h
)i�|�0(nG9J����5	�#�)��rpSR��
ߏ����2�]�ƾF�A �ț�/� L��YJ.�uB����Qڒ��6�&�f�y<}`X��B�MO��dV<`1˝�����S��'^�\� 0噈�.���N[M)=�l_�zd!@������#JM�E���Ag�֟i$^��'��w��������	б/����_ޅ���ZHY���Ȣ����I�{��wd�y��+p|���[�4	2�*��(:3����8�)�I;�5`���֜M�L���K��q�\�����IS��р�pa��1FQDՄ�WPH�&��,���5�b�"��CxQ�8h�T�A��t�C����
��3��u�	J!�s�.���Pϖ�E�X@�D��d����?S��NJʗYJ���'�����|;��Gb� ʗr��W�'�û�������.�|�Y��䲨r��TA5��[���A ީ:�a�:�*��K��-��Ne�^�8N��A� ]��м��_�y;D+��l16�̱.��c!v�J�Nq�=w͕�5YQBD�ֈi��G�kR�q�f�O������;�Nܐ�}K���N&� �؉\~I��Y�(\	*;yG����n׃�D���qrs�����Bݍm: oG�ݍ��a&-����z3�m:���+�2���$J����n�"�C�>��.�r�e�Hf�
y�q���dĢ������\݉�MPT�?��ɠ�.`%:��&�����GeU�Mƅ;��n�4Ft(S֯7Oo�Z]0��^�#��HqpXF�e��,�5Q����$���r�������˚ꖯ�s�7����4[�"tXe�"L�}룅�58_��P���7+��2u�8E��@��)��U�	�,��W�7VA��@�Y��8�#�����3y��i���z����5zc �Ӹy=�U�/�˳K�t$�Tk@�RQ�w�X��il��e:;D�n[����c�d�H�O	fʯ�"��r��Xa���b���dj�H�*���P���f}��j�2��q�>�:��?8\A�3���>�D���۪r��}3�����?i#E�ѳ)r��rf�^h�DNx�v�� 4۸Ҽs��	]�v�@םh��~l�?�v��
~��|ӷD-�E�ȬJ}?�#��z�uzS��ۂ���G��x�:{�9Co�G���Jx�XR��_2�� 4��d�'�s��V�S%�S~��*ϻ�q��Cn�k�A@��Du���u[u_n�4MLW�)|q�O�4���3r��H����[���rLa����������<���� ��5��6�e�o�������T�$;�ԍ�k�l��F�t�}�G@-k3y��.��s����Z�.��p	^���R��?���v]ĳ=q��'4���AO�ۭ�F�mg�d�:��a��F<J�FfFv'f]�<"�Q�HK�����ے�}�>4��/ �8?%����,��h�� �:�t�q�w6�Х��zNnX:`�q���X�&�MtZ���}ޜ4@.�ƻ��2��&f�_���F��¬>�d1Qam���]���מh���/i�vGDZ��m�$��<��? ֣�lK*�=���K5z���|���^�S�?o~���c�Ԑc����&�s	������/�W� q�����MË@�]�(*f����{y\��-j�<�� ��2as�5�Zw�r#���鄋M��F�mU�f�g�I���n|}��l��'�[~t\m�ٹ�	O�V�r�a�L۾H'/�m��J��w��dΐG>�[ЩF�/�_�w7��4��L� z��[��7)��J����O!WX� E��`��k�����<E~�'�/6#�9��q,�J�߱����3+v"��ާ��5���j��V�둏�jeBߝR�>�������$f��WN]��m�m��i���Ԏ� 2~�U�x��/UU�v�۫�k��?��A��ͮ[�͹���-h�p������V_\qbѷ+_h1�����z�H6�@����Qĵ��f~`P�(�?8C�s�q�(�=(qo*�A�/rn8
"BJ�JJ��vi_�&g�ٶ_sJ�u�.�kS-[�#�hN��!aR�[��oĄ�!iKy�S�	���,���?�ͤb�w �n��pbM�����{o������^>�aJ04l=e�iJ��ч�q'���_p1�J�$Sc�t7	tk�

$!���ʤ!��;����)�U4�lS�j>�Yw��C��૛���NA�,�$���ç��^H��	��0��qp�(I��.�_/��!�l����I9��ΎC�3��5%�?7����k�ž�ޠ���i�op�*"��b^7p�A�o�z�^�5�L�u�96s,&|2(�L=��}#z��EH{����_�_��Ծ5y_D��˄|�}s҇G/�x��̱�N@��o��\���t8R�3c�1����8��y�~ C���GIor,���-=��KB�]/��q����$��n�Z�ah;	����4�T!=��W��@ �T��X����[��X�8֍8?)ō��4��a����&] -���B��!b��O�Z/��Z�u��avR�u�\�X�y�>:���@�u�O����A�ul�&��BC��A`���G(n��v@��6L�Uδ�z�#�zP̝r!&�I��0��Ky���Ћ��E��\���kM7?e�����`�lFp�-���['��P:��^d��E��|�eH�g���l���~��_�����c���O4���ɏ�Q=Il�DL�9��?d۹'��AW��z{�����&00ͺ{h46����3�E���Ģ�\Sn>�ѕ��J�:2z/?4@&�����C�/(K��;!�h��L�4�Ubh��7?��ɿc�)+���
���rr���h���g�,�~�SM�B�R���r��2��=	Dώ	��Ni�\�����Qj�Zq~�����]�@#d���X�m"Π|r]��k[���È���AX�(g[1?�7�e7Q�m\\;*Эi
8Wr-G[΃%ͬ�	��9/�^���QՕwZ�W�>��W�%6��I�	(K(��G����n'{�!�"9ΜY[:��d��@^U~!�/v�9��v����A���A�%Z?�A���|�e�?��g݃�]� ���젶��ޱ;3�?adQ���d7 w-Vii��wK�W�' Z�_`�vo��s�ydX��{��۵-OeW�qf��J���>	�{-.TU�ϼ3k��� N�p���AH�k�WMz8,������g7���]aRQ���!����31Jё�ٯy�R��L�=���}=#Ws*�����V2����\��~4�,��S�`���ml�od.4|�,-�7�NV��X��2��.�E�%���=��
�E����3�w�.?ۊ>-�ѕ��z}���h�ux*<a"��z��n��Ɔ�1�*W��4�<-��_R�@�Cӱ�CN�5vO�"9!\�]U�o���b�8��@BE�M�0^Fi�m�\��3�����BS�>������uE
�����8@�.�h.��z�ލ�{%z���s�T��u�>*��~|�5��8]#���K��1����!/5����`�тH�uV@�:�Xu�j^�#��v;3&Z�Z�Q=�_�o�, ����LO`IŘ0Ie�&cR&����*�ԕ!k蕕ߓ�;^�[OP���S�Z5N J�`S4��x��}h�`[���5V��`/c^�	��A$�;="3۹O�J�'�P�kTbm�=��6�d���f_�%�]Oϙ�{�ᘖ-˒�f��$�
���l0������2QT���"��Z'˨��|-y3��C�s9�gɬ���:�5!���k�؅7>蚷��{eE�uH��s���6b���"T�K.�ҋC-�֯#[U������>邰f�IY��b���t߯�ч�`�pl���~�xE�$:ỉ�1�0��3?͚��%/����D���Ѹ����ݠ�+N���J"��x���RG��I9A-��7��$D[ZT�,,��]��\	h⌟��U�йʨg&v=��c ?:=��8혟����!�	���J)�Q��j&͡���|�{^��UDr��:�+���)���C����T�^� g}�$t��t~�9c4��M�b�]��m��oA&hE;�?� �6�f�?�5fk#?Z��?�����fd������R�G�����p�V�Wts�@�a�eD%9ZmQ,	��O������a����@bS,+���� 6���1�;W�~$+�>�{;���5/k%�{x�s����{�!7�f緷�*��ߤ�4�Y��FK�Gc�;A�$#@^ڇ4�J���|1v8D��'F?D&whO�y�~M�� �
� ���qw(��7X�L�~j��0\��5��Β���#Vs�j��b�F�Bȟ���Cd����A��/�X>ß�:Cae��m���n��qn�qA�1��0��-sw�n�-��Zz�o��f��5p0v��s,!M�)�X��'޽�l�i@*s��Q�nY��P�ئ�������	�����f����%ÑL�^�32�1P��k�E���?���i�-�wM�c_�Hs��RŝЇNѻ��͂@�K�S���Pwg�8���/љt*e�+&F����쬏�2�^�O�W��Z�UJHv������^/�|�H�-*���~��a����i��K��jjn��L��1?bB�hH��(��!�j9_~���^�`���b�~�:�狞�����%.��T��AV��n�9�;�>sX�
A,.���g��XH���r���w[�q��ɣ$��_4$^�2��md�-țZn���ڠ�2D����'E���bq\3�z�91?5�:��j��q/���Kh�<$�`L�!��uq�
��v�p��ٺs.����!b�:.O�ϰ��y�ɱm�4�E}v0�7'�qt�������n��q���8S� u1�;�|�~3b%�S������oJA֏����,��љ:�uh3%�e��&:~��z39��'.����mqnv�eh8�Wԝ=����A�B���rGc/��{v���2�huMئjP �S]k�e�-��{�yms~�g�`��Y'��ʜmbSG��Hrj�|��z�:��)X<������ �Rϓ�Z���G��o�A�W�Ǻ��V`�7�Q1��k�	�.g�X3Cd��D����9#1j�#���C{:,@!��Ep�P�2��k�P�I7�����؋�����In.2�e��!93[��+���
֥Ea�
�f3�����
����s��WU��S(�OtP���f��p:o<���l�rcA�á1������&yjNP]߈�:q�Ƚ�D�6$�LD��~����h�F�E�L)�ӛ�g�����$�B���]����w	[]�S���{�*���A�3���(�Q�<óZR~x�[2��dFdC?�y�C��Ƣ�[S�t��B+0�y
��R����z�;�1��lQ���eT�?鵋]㛜g�+��_E���[)⪄ 5Ux�}o*`�-c�7x�a���w�%{�4��F�S�wף'�ŁE�TrA�DJNh�.\�Y�*�s�W7��Z�:�>ig��Kh�|�5�o�,�ȕ(9}d���헛�!ņ�Rc[b�W ��*k���bh,��T����;��lIW���	t��Ǵj��6Y���pq���8<	Y�����T��!� ���Cz��Z?Xi"c�󧎰'� �5�2��̪2��ՠ���L�q�����[5@�wyj��]���?��K��ea�q)����s��-y
��7���9H�4��!�/x�@��[��7v�/{N��@#��X:��f���B�l��,�������9}-_�!�.�����#Ɏ����>�K*��Aw�`X1e��R����*[�����@�)O�a5�L3�ؗ �nLfO�OL�99���qY���X������<s����<2��RQ���`���Ә\�U���(/�[���qO�,~� Z �����Js� 4Sp�8��5�ʺ:7�Gm�$�+��6I���5~�2�+[�0`V��}���x�-��ɒ�x� ���R3$7��=������R(��,�$_�h���]�����������!aԉզ�л�ή$�-Q&NS,��"ne���AQT�iB�3�-�N���$%41�;pT��j�U*�IT�v�[�!�
�ǂ��Az1�v᫘�	"*�0ws_H��<cs�~���{�D�~�p�/7	�Xa�\�o��~G����d^�����@�)�l��'�u�]:
�8����+�U��7�\<r��m�s@�η��U0S�,6��oX5�f�-;�bP�0P�p�^9�ou"T �9*���9H�ĉ��^S�H�ע�o_ڶ�����l{�+ף�)[S��$�����?�ENxl�,��� X�R]�1ǋW��)�����TV��6���=�����¶Y�|�� �2��ʀC�jx�\������� z�dT���F��"UÑA͑�a9]�|�o3j@�#3�9�FH�BK�!D�CbL
?�
Ʒ�~*�s��� �	ph�Fo7�ؘ߂TQh�NZ#�s��y���[E���_>�+��Y(^@��Fȼꅎ$�&B</�BĀ	�2ꘟ��n!~��vM�B�Z
OV�����'q�o��:V- X�p�D�A���2�UDo��E�z�:�#�J�H6���mE@�� � ���7Daiԕ�cn���ME!�C:�_*���ӟv'c����� X5��(yo2n_sҧ,n5T��W�A�l����M=��=�͵E�n�,�Lg$��B�W�M�}HY���'�e��m�◉��̾�����,���*�o���� �% s�x,��mgbɵ'�7�{s�=L]�Anb���^2��0}d�����x��E�"�����5ę�$�/� n��j 4���x���7����
K��I����UG�PܵR��ܤ��|)��<z:)µ�K�����3fQ�ٿI�eܭ�ftŕ�zԮ��sB�[�e˙��!{��xX$8���a���:��/-]�K��N�6x㠘�M���Ē-l,1���	��\uQ���X�
���.OB�a=���]�.�����';7(�h]���O�a�lX%i�6��sIq-w͔[;�k9��?Y��u���Wj�B&�m0۞S�HW�#]�PIZ�f�5�`e1{����s����p`�X�j>�������j3��,��x����x�ز�a[ңb]�Ò����skH�:���K6��o���	W��r�dpP�Fa�#P�B٧!�]X�=ʓ~L��`V��b��@B4��O:s� �A���1l��:P셇ale;�>]2����QT97؏�{@ɬ{������?}Zu�	\	<��t}L�)�� l
����WgX�֡J�>[4i�)R;��w�T��z��"���E.ݒ3)���z�������`t�ZZ9+\&��m[��
��7Q�j��@��=9�kvl��.���3�6NQfw�"����G٪���!=�c{:�C�)�t���;�j�W *A�B�;�ښ��e6m��Վ������mpV@
��"�R+�dC;?���!�'i���O���M�Ԍ`r{�`P-�b��D[
�!ַ��8_�rn�����W��)V�J�S�M-��ĈL5t���^�9бO&J�Z��h��z^��~����)�Y~��^�1őX.�U��C�6=�v�-�!��v�b$�t
��B���s�k��[��W{-q|!���<��	/�P����҅[����u��Td�p�p%J0�A�C��`.��f���
K�^o�IZ�P�4@�@��#��.�wO�9s�m�a�玐r��V�@��I0x���ΡgA��|C���nG�&?�fx�c��.��爠Y�i�c�U��Ʀ���[�'��Uv=����y�zTg}�zK�X;�0�s)&=�jCC�,U1�a�|VYLy��V/P����֖�ss������q��˗�Ҁ�I�X�t��p�А���0�ё�,.��i/��@�	�X'��dLCm*D	�Z�{����8m��+V������{Pk;�;\�����5��-oc��\1��䐞~���Ŋ~�yr9�C�On�(�X$<��+�c�b����U��V���
�:��M;�+51m�{y�E��՟�3�b�HR�cܾ�Tֶ��VF#(J��OK($��?� ��a=��}���z��`y9nx����-٦j}T�J
Z(���*�9Q�n��1\�_mq���<n4�>:eՊF:GϠ��#%���S[Lyghf8�n# �c�.��m��>�閂�R��q �쀹c}F��;�dX�`j��n�K�(��X������ö�u�*׿Ĳ��x�=h�]�!m�e��*nVQ�<[���h���k�� 2A��3��۲rK�F{��? ���2�����-���'r�%j���- @g���b�N>������*��ޜ�ʇ:���OvJ,f�?<�BB:4~��_��c�-����3[��#!���H��ϑ9��%ٷ¸@4� �*�i4�O����g��}�����Ln��&R�,����6�����c[@-8�yT��:�3�6{��Pu���=�q�_��A���s%�l�كiZ-���}��^K��B�+�k�Ke(��}nf�V =o�]�!��eСP�J��'�oX���@ª�C�8P[�o���B��d��R��9����{�o����]�;qVٶ�6Cg��]e��>��Ԍ��J�8G�� �4K:?�n����H�y�������&N3"@��Ȧ۫����2�؝�r�9C�j�ѰI� |ד�(%��T������`��C�ģN5[�w�=2�Vg.�ʽ��,�ՙ�O
�eyC
?f���O�%��_�<R��U�(B��5���P��g����{U�o��ؾ�w�;��M;X
S"��O��\��� 
\�� �KH����BDu歩�.Qe1~�%��Ҿ��-9D�pm|c��Қ:NGi<q7Q�$��!�~۞72�/��.�V{�pP���6��s���-`KtcG�; G>���*�y=��tq\5q��~hW�
��8]�I��&X�U��Y8i��$����S��ױ�_��k6X����2���� ռz�&kb��.��u?mw�9[�@�N����N����HS�+CT[I/u�8}���ܡ�#i]�ݒt�!�UR9����ﭸh>ǿ�[������3F��� h��w�K����,�U~��{�G���~	��jG������dX�H��&�b�:6Y�t]�OUg_�0��Xn&��}����g���'�؁%B��9md��x���e��}i�����&��	����]�u���`)����I�无͚f��sEwɄ�Wf�fGL�e�/���`��y}�����^$jL��n�H�39B�,�
�d��{�����C��_I�G��jb`3=�uW;$DL�1i�t�B��/\u}v9�.5�|@r޳0��MiӆRK���"�b�4[�a��J�Lh�_�+�$1׷%M ��!�c����IL�J7�q��j�C�L����7��c�45�@6�#�ȆX`ɀmY&��?,�Cz!{2+;_��h� =��*���J�y�8�d)�s�<�`��z9t
�)c	�Y�>�(iZ�����U�����`>߷��� KV�B2��DU�!��Ss�Ʒ���!t���#�m٘�)��-����ҵ/GO���;M���)�ɕ�ϛ�EG�,�/���+d<I?��J -Cs>��m�%P�����>"����J8�N��ۻ�7rz���ͺn�X�=E�����]�tVT(� ڬ� �4@������@*���n�T@��s��C���߯ɜs���n�)�l���ݻ�8�uW�"�n���������q@�q撾��ѧz�Ł�����_i���`:h<;�\�\��z�P���?��[-�UJ��3.8��="��glP
�\I빿y�Z9�Y����#���Ɉ($Ǡ,7����E���xZN�WB=_���/Y�]7L�o��C4�KA3:�&osZ��ߡ��3?���69��.x�k���ʻlg%�F�^��1��8��zo���~]����M�
��Bfk87�1��I\���md#kH�����7^�#r��<{�lA<Y�GV��Ȳ�:x:�ĬOɣ�׮���Bnѝ��V̧��R�Ϛ�S]�c�J�'l�B2'�R���"^�2�(a�R�����:n6��4e�8/F��@�b�w�/�^���^�Kyh��m�`\D�/�^��%���M;�� D��s��2H8mf�WNA?4{�V��K9���2T��єL����5��x�W80Ds#_�A�Q�l3��vvfc
�k��ѐ�ts��,p�$�i�HԿ����؀ �8i|���E�aw�6+�꧄Z������3��\�Y��a��\��ڷ͖���ծC��,J}�7B����("��\@>t �C��*�.��^��XG�~�UM�ߦ���w/�Ia%�9��[�@`9- �mp��ꡳ[S��� >Ҕ�����F��]�����i�C�9�d�K�qq+�/2��P�Ne�(l
�&	��ϴP!G���Kk�l�Ȟ,���B�+O�#�p�.W&u��̕���EH&�@t:���@��<|4��A6*��c�78݈�!�4ǆ�v��
��X�ݷyWK�F@h�r,��*�U���B=��@
@�����Gm;b� ���K&�Z�7��T��_��%�s�گ��Jz_$�b(F���V84Q>G|����]��6eN�~I��g����m޳�*����q4�u�f��.ae�~��eL��%�05~#_h����aP����;��*�ۯ7<�����J\��>�"2geA���*}Vzٶ����:��A�O�� ��e�����Vá��E"T��*X��_b�6�L����$�.Q�-z���Ɂ
�U��_�Mx��J�O�':m,��ꁛ����!�,�W�7���j(F�<��x����U1��Q���DO�!<�;{�5V��&�,Q�Tt�Z+s�>�w�P�;�P!���Ɍ�E��'��]�����)�;M�X~�H�Yjƒ'e'(���݁T�=E�p!wkz��If������2-2�L���L�z੆II��"�v�w|,�}����m�(��Z_�h7����>�e7���[�IbJ"#=�nF�EPZ7_�Hn�?��Ǧ���SB ���|�ؗڜ@��� �' :W�5Ϭ��<$[k�?��uf���p%O�?}^W��u��>#J�w�d��H@���I�y��,I}n�@��q���8����b9@�_�Y�O*�js�m��X��,�OH�A�d��q��8g�C���D:��}B�E����h�Y+�d������������01g}�LG�G��.Gzs	�-럫A$(5>��.�R1�>�*۽�Z��Qw"S�ZuL��Z���s���
 ?�'�b`j�b�Ԣ��X7���!������{��_f��kU_��?BT~�W�-��� �����7K�h��7ڣ?X��i@�����+�6��;)`����N��7م_��6��H���8�`�]ɬ���C��DT�:S�UZ��x�y��&��k���҈��6Gx�<�-�F`V���DR��*��t��<A�Ȓ@���=RI���ո�������7�Q$"So�8�X��P����������J�"�|�\:��=�������45�[xZ��N�}E'�����qrʰ�e���gE!c�8��W�M~h�� ]�D��S������'ݨ���^z�s��[���|�� Lh�l&�H�W�IɞIWG_���#�/�]3©@Vr �O{  v�W�C<���u��[�3O[O�B�L��G�#��~P����]|A�&缘m-�8A����$����l;�d�:aVy�֬=��3�neo_���������������������;N�d��BW���VƯ�9�<ox�aWˬa#Ī�Fɝv6�����l<��Z5�8a3�x�)G8�ԣ'�� M4:)T	FK�$	S�%�s2��Q�����M��HT�<Ǫ�|�S�xԾ��˦&W�h��$���j�o2���A|����q�Ö�����g@3&�&��I��h���4����n@�(N�DF-�$��y�gb����GVY�Q�o�5�*��\L/�_����='�k[JFi�(�y���~��!Tm��A�&q�Hjt����t�A̮����o��QP'�b��#R�ɺ�z�[����{i�;C>uD�^�V�A����cki���O1���r�$@0���͆�Q0��!�I��*�;�q�^q.�`8&�>�w�,���_l�e����	ݶ�{��u�[]�s�-��-���<C���.��3���C�a�@��$"��ow7�FG�I+b����?�_Om�3v��=��-���Fl	��>�#�ç_����K��8�kNJ�mQra�y��7�Q��� I����-cG�K��tں�$8��1-oeX�{Ԭ7er#�F^�0���K'��9�)|��Ӻ"#�����Ɉ��5�t�e�����@��
������6l�n�������@��=�z�FC�V�0n��u�w�3��2������X�� �!zkĸ��S"O��$���!z����Ò����T�k
We@�2�ڪ��'���p���Z�a��(�r���wb!�2���J\�D��op��˚ތ ���H��}3\��cc�#��o�8��k~>�g�|�D�+a��_F��UPڕR~%c��w��a������q�׌�����[0<�p��P�-�6"��X����װ��j��`�pa�
/!}�ݚT���U�CO(�>�Ĵ���e��B�M;e��	h@��������60�0�WRe����p����*�����]���W�feB?���)1��|R�5���.Ӳt������̀܁���x�G�&)48a��d���tbSiJ#��5��L����>9 �mnW�߸6��c��ݱ�7�G��N��!�?�M0�t<��
�*ޡ��� �j�����F���zܮL,Ћ�B~�k���?fQ�9!�y���83ӐX+Zz+o:�\2?x���~)�`ۄ< nX���浄PF�D3|�4o��qS�;j!���$K_-c`��1y��dqR�^��PJ���K�y��d��p�c�pq�d�Q�)S^�V��9WX9��i�P��HA���[�ƑP
����N�#�K�	��C�Z:��,���st�7	��m����Og�{��[�,��LY2�hT�ȒٹY�m��i�H۹U>U,�������6�e�P��I[	�#فZ�N�I��h8.��4�k�l����{1b�u����z>Z�0;JИ�ť���6'DS��oW(7G JG��h8�� �z�V���6�ܚ�y V)N�9_E�r��mK��oxZQ(����E*������W��K*\I���b�"૯,��ı�K�|�x��]����/P�o8ZqH���BV���v#�P��h����"�9TT���`�����`-(P�AX��{$N�^���R�X\�B�x���P���1,�>Џa^�z�\����4p�p^A�d��*���L�wY̤�=s$�mvb��X���!{U'���?�Ӷ	ٕ���>!��;����:�h�W:�irힷ��kG���XR{�*�Ee��,C� ����~����5���ՂAc��bK�f��`TQ&�Y�h�}�1N/�9�2K��F��t�xHm��ݦbYLd
�k��wG�>��NԐ�+Q"a��h��HGl��}]����Z�1�T�ζ���{����
ƕ�:տʛ��iY������X�&�S��q�+�3غ�q|�u��c�Rq�sFg��������ն��ߩy��-R�lF ���eD�AK�hq���D��T%�g���Z�ũ��S�j��Ӝ=u�~i�œˉ1�~�,pP��5������ϱ�a�i�H���յ�2eDΧ<��IV�Lk*Q�{�0!y�ftIҲqG��YFf��ң6�t�K����)�U�	�k�UcQ��Ww ��{���8y�+��3Pޏ��¸k�Q���ч�n�$A�D7�Un�(ɗDq����C
���a�+f�o��P�|?0TJ�'^�yE3���\#��#���A��$e�U6H7Ah� !x�p"�Q:��l�j�d'(����*�|�Ag&���m�#��	=s���� �H��=�-���K`�Ӧ�ֳZ�*っ����O8U�~�BIH���P��8l�0 bN������F��H�τ}l���#*TW�a e��P��0��R�s�B�M�˥�p�v}mc�H�^�?q���s�a8  8�J�TQ�O9``ߝ^)k��zֱ4��@�	�br��Eo�/h���3����^�jmϲ���{�]|�w��W\��%a��������&E4e��ƇK�Ѧ��v�ᗦ��0ĝ����p8m���SF� �U2[�	�RI/_ו_�R87a�6f�@��v!(�{�8.@$G(+d���;����h�i��!�oY��z̵*r�ף�C4c�b-��ǣWt(�ms��dJ@a�x?�4<��^7��� !����@��'s�ݕI��
�Q���!�gy���ĭ�{u�.݃�R��+�q�gl�!T��V�-=��h`�j�f���b�$ʶ�
iS��ws���p�F��\d\�\�$�sV���
����Zy>�v�(�d�q�����(}�=lU�A+����)�e�JkJpsˣ�����c��1�n;�`����yD%�*��#ՇBr������)M��B[2�$i�JW!R;�Jp�,��U��Iۖ5w�ٵN�ז{�ؚ]H�5au���ҹ6����<{%�����|+ؘ��@l�P��WA�7�zǝGF�W�Ј�k?�͠��B1��,p�J�6�X��U���V���!���v9W�Ʒ��
+�	�ӫ��|�|b���R����D���Y�1�v��}��j�am��<���)����K�]��@O���_�)n���Uv_Xci�	jɢP(ѿ��n�n9��7�:�����g������W��9�!&����q9���W��8`�F�Y����04�ʢP7��pHlm[���9�&(\����v��R�UI�U��ɛ���Ee��xd�S��FW~��C�V�{7��S��U�
�'��"�r��8,�U ��Uj_y��I8�q(xM`��i(�O�y��0��;8NA\��[�QXWv'I|CvG�bU�M��PZL���=S�P>���;O�9�_�5��D��h|���#Xs��Ѐ��ݐ��e�Nv�ܶ
�ݰo�^��n�eX1@mے�q��8�'$��o`�y�1��;��V��j�0�Yޫ�~c�N��FJ h�k�����Y��W+;��/
K�u���J�*L�4��C9�1X�z�4����A���A��j3;��B�����1d���5z�=X�G�V���뀄\ۄN����j��s9m]o��'���bRM����ݵ(E�[D��H�>�*�ݼ���b�N�_��X�.���z70�a�����@�&2q��A޻�dX�N��K-F����q��3Ȅp�jK]�7�#k���m��ѵ�O8�zTa��%�P
�t<�"͵B4]O�E|2Ρs�/���qĸ��y�̧p�z�Q|�k*�5,
���;�l�PX����8:~��$po쫀M-}��	oU�>i�1�o����w�OE��L�4���WtT�30q��z,.Me�v��Q<U�L1e�Ċþ�Y�Ct�1G��G��q:2W�!�����U[�z�Tu�R�Kv1t�SjT�{�V��nAS�:�Ǔ���l<V�.ic�PC�".���!��S����]�D	��)i��q�}�I\���V�i�@�T����Fe�,΅$+nD�\d���(�����T�*muZ��XR�y�>��b�0�c�:+7+���^�ƣ��ZbR����iV7�.�Me'���ʖၻ�SIyi�[�kq!�1���WtÚo�����=��\Cx�����A��C�@�������N��l���ht>�_Y ��d�4��f��=��5#���P�#�B�˅>
�� -pH����;�uA���?v[�W�Q<�QK��U%���?oI@X`���B���,��B["���;\DM"J5]���=�L��:I+b��1	j&��v�"��Ƥ�����C�;�G�o��@ZJN�C� �0��O�������N�9Q�{��w�$�Kb`m�j��EG� �r��17���Â����떋�v|�-�{��x�3�W���l����U�!����K�f֘n!f���"Ŧ���F�'-B��O`ߓ�/��5wS�i:��C
/j=9c�i��_����H����a���5Hb�����?�.�2T ���zmB�ֻ��7��G~g�vm~/�x_Q��k���Z1�Zp)y��IؗD���
N1��q��l柷_��:H'V��5gWԚ 99,�_�j=�5�L_h��{N��	Gď�HȊ��uMڕR�"�f N�=C�U�A�A�wέ�Gso�4���X�O�d+�0	im��1��7���:���0i�A_���	�Ws�����ݱ�����[��6tell����+�) �m����T����Ȍ�w��*�:�J��w6/^�uD��P`H����kN]݄���|�T�*���h�3����z$�l�J�s������Z�IM*PH�p�fU�6RX�'�\v���`�Ŏ�_QLu��[d�<&ɇX ���=Nuy�{��K�/�����W��D��9���d�}��x��8�i���En��^��*�b����Gi���?�ڍ�h�����+$�'Z-�v���� ���=��uaU��)b�����L>�nR����`�0�6�te�&�?����Tc�|������ sݼeHΠ�
:I�]Q��hlq�y-7��U
ˣmrcl]�g5�Q�h��K�S� v��0c$���L��"���l1���z�R�zq�:$J�������BI��h4����4t.L-py�eu\�:>R�n�$�=Lz ���L<Ś]����vfm��ۅ��E�Ĝm�I4�Nz��ia���t�)7Q3L�|�c����g��+���<%���`?��8�����)���H�	�!���h�Sےk���a�$+}��Ӌլ�'��S/9��<��*3�y��'әOk�������O�]l��"�"4\8��o��W����|\������	�NB��w���]qV�<�q�����8Q�fr��`���>֒���|�VF���G8d<��w7���GN��a`���(� h@s��Q`��NnXIpP�0��	��2�_�������=�z�py-��.U ����}gS��M�
=n'	x�Z01��ﺟ"e��MB)��H ���I��֑�e����'��)�ϭ�]uz"z(�A�S�f�4�0؎��HA<U�Y�J�n�~J��R-W1�ba��3x���A���z�WG8��gD'�3 f�r��q�L\W�F�{��`���|k�R�}WFm��>���[�s
���i<�?�@�,�w�mw8��|8׍����}#g���b����|_��a( �0�G`F��CE��;N��Dt�k����������`w�/�+4b>˞���l�E�dF}���㽮�j~��!ɥDE\��qca>l7ǯ���v��u &�h���6-�\��Rd[J��:��F���f�� ����_A����G�]��O���݇gܔvԍ�E�^���}��'H��=��Q���n��(�:��Ps;5yc�Qͫ��x��Vԏ��hbeW��yv��[W�e���A7����Z�Y�l"[��Nn�C�Oe��H��M��|l�c�����ab>=�u��}�N����{jGێ"�[�]�`%�	�����I�'�w���.�m���%jq����M��aQZn#߂�e ����S�.W�Eԗ���mu�	Q,"jU:�7��3���L^�������� ���V�eYI�?q"���%�R~�|'�r�M����p����u#�������+"�T�XMO�?G��n��"k
f+�_���1b�-��\�	Z�����Kir�p��qk���4Y4�G̚b^�BaRޚ�l����H6�����[�� X����5��tj<�"n�U�D<�����u��P`Gؒ�J<%H<@�Ń�/B�Ɵ���HN��ChS�~f��
�BA+�׳��!�m�C���R�>+:������Y5�=sŷ�]CC4����`���&�#�p���pX��wA���^-K��;^cm�#�)����`e�DG:b�h.�XB&}^�����EF���:I��o9d�$ZEN7��P,+Bդx��k�Pw�H�;�2��5#����9kO�Ө���W��f�Ȟ��nĈ���^��k/h:z:�r��2� ���$>{c;��n�i�2����Y�G]Z��NDX�d����7�+�5moӉ.)�O���6;u=�V$��M���J��$�(��)�,�rJe�N�U+���ͱ�*���iҰ�T�ƟZG��C���]mU�T�]˱�� �0�u��O�ۍr�1�*�P����kA���Ɩ]b	�M0@mޠ����.��@��,P^��-}�,A�{�9�i��-K��ѣ�ڐ��*6��0\n' ���ǱSK�f���х�E�H`'���P���>_�Jg������8�|�!�T�!���}��"�v��Tق� [���	(/4��A�8�kI]"��gB$VB�Q�R9ͮ,Ú�o��nm��t��P���2_h�[��r}����J��1��7��Ev�{JS�B
���<b��F������#�v�RO[�
��@�k/>�R���bs��0���[a@�P�Y0�̈́�\�!=���ä��.���N?B��~��I
�ssl\�<0�������1
�2L1��r�A9���K9��M &S���3u47��=����?G�
���AI-S�{Y���yGB��Tk�pIv={�c�4}�צM��v�0�o�FS� �}���t�X�3�U�|SdFy4V<���c%{�ɾ.��m��A:�}s��ocl���zq�}'C���|<K��8@pA�-~���M�k���	@��,r��e^z�=���&�4MTH��T�_�É4�p��#�w�!ѷ�cR��=�4��Μ��/�������;�!~y:��;�Uϫ�%dҽ�gP�=i$�4j�$.�"b+��y#�J��Oy�[�j�t��
:�T��EQ��L^aP��9d{Vq��2��m�5~��q�xM��n>zp��S�<��6�	y'c�?��OE	�?���j��'��=6���G��K/y)�_����^�I�����q�?�mQ�x���B�~]�,�ĶD4����i�%����H�s�q7.�iH�ŦE5[�_�"���c����K�Vg�ϭ�ۃ�N�$����/`��'Ўc,.��0��y�_-�.�.8�Yڇ]� {VϘ�'�l��/�5�!�Ip��O�eJ�Ó���*��g�u |Bd��Xz��6 ��I98�vsD�2r ���c�ѰTRA�`lm^�����<ʡX�	�|�;m��3�v(�������"޾]}ӯ��N[��3>�}	æ� j�/��[hT bů�Fqn�+�~ej=:l��≛6kT+����G��:@G��Uj���l> _�B$���]4���4�h��q�Jly���=3|���3-���K�7��z�u�mS���E��ʏ�{@���Zh	+/
>�u�~��${ˑ`���K����u��-
@N`T�a��Y.��%E�U,&t��C�C(�л��X���nݿ+
rq�Ԭ|����~ܔC(Ě|�&�ݻD�P�H�4��xy��? �g?�[�A ���NmT��4IF�!�B�W�G�|,�-��vc1/X�\RQ���Ko9�o�+?*�W?�S׃E��[��◕�:|����"C#��"x�L�{%&��x�}1�!�J�;?f���s	��qb'�pi(��&�,��[']D��dȥc�S9�۵�r��t���"(��qJF\����Qp��b�n����٩�;Z9Ok���ijZ`�cY�~f"��zͪP��[��������jBT"���Y�M`ˢ+U�ZJ��d.Nq+�y.�j&�q��Kd���׋��Na��F_�{�L~����'C���K�v�̨��˩�c�S"����t�Bq,~�H�|qg�\C/���縐���K.�ɫ	+%2�/�YT�I������t����UM��dp|��e,tj[0�%�'_��u&% N�͟��և�P�*�]��{��Gײ����_X�vr���ɝœ�;Y�b���{�:Z�v\f^r���!8Ӈ�#&2{�U��A1�5���p�rS\�i���(i�1���]dM?c��l*'!}����URH��Y�e
@�SX�tª/u`���l$m�q׹��r����\dJ&Ӎ���HFa����U|&`򱦅�=┺	 ������JJ����Ung*ɚH�5`�2��'&B�tvﲮ=��{۷/8�h[��Q,�?{%�[Q`7ɻD���-PH�Y|�~����$W)>��{v/[�S���M�b�џ�^~�/P��ߕn����`Ꮩx��"R�u�
�	��/'�'n�eO���(	��s��(����E�I��>R� ��<Y��N>�֬����F�_u�{���]H��:�?jf�j0�]n$"4F^v��?m��Q�)f��	��&l���%��p8�����n�O�[�k�����!�'r%`L�	�l_/�C�s���-�r�ǁi�_�n�~"��XrA(�e���ɦ]`،g��]s�o�(�j�C@���qC'Lx'?1L����1z��8H�\�e%�A�1,/v�Ӧ2�=9L/r�29�P-vӾ��g�������3�����aAyC%:(��K�}kd0�|�nUq3���pC@��оIs)���]2�H:�
+�v���.i{Y��62&��Z������N��y��� �U`������?w}@w%��j�8ϵ�Ǥs��Q^��P�P9�6�WY��yM������$f��R����H�c떆S����xH�jv�HN�ɂ�y�k�*�
F�x 3{�5�]�������}��@��n4��Mx��UVWO7�?�1�Y{>�9��ӫ��ŭ�WF�!Q��X�k�ְ̂ݠ��;�M��� �S��Ҟ?������˵An\f���:��zA:�"��+
溾*H��ƚ<�36���L��M����w!�؄�tP�τ�p YЅ唆��B �;�b�M�%�e���2�A�w�p7yd
����TH]Z�q֕�chax����������P�R�j�Ɖ�u� �e�^� �+Q�l���.�����B�z:4���"��	9��Ԅ��'B��v���j��%RF�L+������!zF73�8U�]kB}g�M�b�5DVw�%�^d>�]��mc1�0ƚ���:��Ȓ�+���u�0f�2�h�g?XcA�p�W꺌�W~uLM�.l�t����+^̒G��^۬�����Pfb
ґ�F
n֑ �@%5�Uտ�lƉ>���-��������T?��`�Y������@ �Y_�({U�s�.n�+g�������ٱ�?xU���UBNA%���G˚>�RP�7�U8���	��������Efb2�c���\/��,�2+`��7��O5N{X
g�r�^�	�.��l����1�v��#n�sڡϥ2���%����6���6�m �W+�nC&�'W}�ho����H������Z"�?�`Meg�h�.����kY�'��k����1U%A����䱝�_M `��q����-�!�w��ֳ	8�P[�7'�� l"�b�������A?��OB﯍,WW�O;��_ۓ<`c��(4�i�|�
9r�Ι��h�L�����b����9� ���{��pg���@$5�β��d��h�sdF�bSڟx'iOp�f2�\f�����u��<J�[G�N�{2E&�1P���ɕ�$���bq�DWi&���:���I�բ�*G;@�wg�Ell!V�oj�لRH��Xz����\����{�s�`�����=
���s�����q�ގ��/�ǻ�[GE��Iᘍ:)̶*���\���p�TS�G�n��>%�V*
��M����w��E:�6H�Ʃ��}�݈�0z��w[��?�%��n�$���p�o��-��.ۊ�泾.��~��7���g3���Eթ���C���! ضYS�8^�_�&��ȈM�J���݇�լxB�>���J���1�δ�������-턓g4�j����c���fo�EHҨ�R���l�&���4���c�#��>�vBm�uħ�&<�t�c��y=O��m9����@�|T̿z���D�+i֍�?��!7��g����{��>�¯��ew#Q~�o���6���4�fޮV�%�����,g���t����xqΨikC����R#0���ǣ������*_�s��=*��u1ݣJ�g#`4`��C����r�� $��YV���1��v�����ģ�����h3�ﳼ1��&�����t�eï�9	�x��c6�nYlA�hiE��I�ĦaF,�!S,����F����Y*xߧL�0l�h"A�Iw�ɯ5Hpc�LQ�2�&r]ZQ�K�CD'o�{9�a�o�C��! �C�>�S��Pm8j��N�K�c�_�2��'�'�K)Hos`�mj�CYu�?�0��.B$@,�IS-.��o6��g��t�"���?זMr��\Hկ���׮���X�!��kv{���]��s�ƌ*�IV=/�� �:h���gY�rpZeO�t�T�7�0َ�ڮe��X���l��R3��/C�贝�^gQB�B���ZR�����BhEf�a�n�h ��$j;��nO���E��
��F��0���³�dp:a�����n�뗁�J�d�"��
R;P�\���@+�U�1�0S|���bd���[��U��x��̘A���N����7�m�F$�H&#�s���		�z�0��j�ת݇�kI
�� ��O wjH��.���"��.��7��\�0)�=�����F\똟U�/�
�ߩ1.��V�8����i�&��P_P>��Е 6�Ӕ��8�I:�RL>O&��H�%�[Gr��	�!�?A� �<��u�5Ar��b��s5�_��'G;���w����N�d�N3�V� c�x�3�C  ��{���f�dOe���XI8���X���	)̼�)h��+ɧ,�.Ѯ�K�x���%#��!�5��\�D��C������|��jx?rf�����A��ܙ*���k�ja���@f��:Y�C�'�ՕA�!�*�N�����o'���eA__���T��{�p�%������/}�<��U"���χ����y'eX���KTWK_T(�ߕ���0d�Bu=?T�U#~�0/\�Q7c�K)K�2�,��jݾ� d,[�<; KY�;z)"~����n�'Xۯ���SӤ)�%̴86"��L�� v�2	:��;�IR'v����Q$,��Pܗh	�2��uH��Y^3�3�G�^��>�r����I�@�uuWݕ����Bu�0Y\
I�<����2��x��v��V�!��PK7q��TY�Jrp��n��=g����g�X4oZ���ju�t|��q��c l�U$�D$�Z�(.H���8k����+`8ؾ��/^�6���Y���*#A�I�w�d/-�^ O��-_�J#z��*�.�,?ӑ#4�Pր�*!f:!�V�\}��F�&�e,6!D��&vlx�&q����gYN�Ż�����<t��ʗG{�c�J�9�P%@px��(�Dֺ�6���(��_�:+B�z��61w�&b��8c��Qp�,+��}��鬆�x����s�{�\�P_�3%��[ّn[������(8�D"�r��W� �ṭT=aN.���zy�5���w���a�:��y.�lQ1n�(/%�!D��u���v������@˅��>T&6��HA�.�{{,Y�r=o��j���/����?����O^[����@� a�D{N��,v��+�kT�X����@��&���� ��3��g`[�����0,�,k��@��������6�tJ�'��~�K_�1�R�f��x�l�����5AM�(��n5���3(c�Z�[�
 m:ak���u}��4xj���9(}S������	�D�=��1���곕礶�Wp~� j!�1D~D�\1��I��k"��L��P16�w��F��_oo�����e�r��RT* ���!Sp.���$�U}9w*��&���1��*x�{ٟ�
�X���cqi���N#���.����v��@P/I<|�'6�j��_M}�jrр-�m5b��|F?�	.�k�p��HH�_s}�FJ�D�����Ƅ��F��l�����&&����7��JK��L�=NS�)�]���W9�#�Dt9[��6i��I~���+e-�5\�|���X�\w��$:�����Ģ	���x����9����k��#7�1��[��N��n���D�ۡ^�#�rdϏZt2c��B�I��E��|���p	��M���pn�&�֤Nfi;��#�!գ���w�MV� )��G�T�m��s��UYC�2�νC1���=�2wF`L-a�%���-B�jYd˖#8#ԢJ�ݔ�Ǟ�P�)첣D�:�c�����:��ƌAk��V���5��z�p.w��5=I�_%Y�pH햴Ce]�TY���b��G!��M�����f�%�n���3\P�(l�6[˄��D#li���)[P�~cOkYK� �SuK1Ɩ��zG 3��v�i��WO�a��c���	�t:� �wA9���R�f#�����5�"�m��Ӄ~���T�Q�\"���z��;$�.q�=C�fc�Z���5�9gi.�����^��5�`:�U@���3?V���UV�aAD���ᨘ�ܗB�[z<#]�����sp�*g�7ݜ��d]������'G�w�w��9��������\2�=������h����0B����͗{��'��pu/�
�m�7���l��FFaA�e�g޾X�!��0r^M� �����'�_�"{
�T��z�oF�zb��ֺ0���hs
'�X�BY��a��nI�rfN(��<X���a�lSnx�jҷ�GU���LJ�����ގr:�9��3�TH���ΰ�6���e�f�F�e�O��눺���'����
}@�����9�j��9�lU�hQ��,�jYKt*G�M��.Br`ҁeH�΢�F	�D�;���$��rڻ�G��m�*�yR��4�*U��F��[E]����e�"�����w��rN.��.=� T�*
蹿��M��Յa �]Nr�J�skמ*G��AD	��n��,V��xW<��P��i��`�]��Èh�� ��g:�?1�0��Z��P��L&�0�|�1�l_��*xu�:����a�5Q} ���20�Y#�!����b�&��qJe(��'���9�0YhʨC��Σ��m^o�@���1V�	-�P1�2KduE-�F�����MĊA8U��"ٌ�.T2�8��+��}��7@m�Y�t�U�F��\��M�H�Q�c�ac�?uQp9�X��{T�a��<R>�X�v�
2ɨ�B0;^A�����D~Y<����h	���H���F-�h�b��c�[�Ҥu;	��W/����*~�䮪2E���
���af�x�%|{ل"I������;qӶ�S�L:?`���]��\���w&�V����̛��
�GW�e��c�8�}ٴjI6�.5�������.Jgb*�*��~9��ļ�N�>�C�Իɩ��zvl%���)��)��n�D�q������d|� �l�5��GX���e�8)+=��;<e��1�Z��5]�� (^�����T�{��"Y����/)���?ˍ���l������74���h�O���^��_��` $���f���mϋk�B`�� 3���ʘ1)ʇe]�i#ũ?L�0�}S�L��N�O�Z����E
�sD��a����eQ��#�t8�⁺�=k�k�y �4�5��ƿ����?��	��/k$#�[�Ⱥ��r����K�z�ð��t�����Z��R.˪~5�=ƌW��
�#"�0�����_z�j��]/�>i��}"�эiۺ��*T���<�u$`-	���a~Oe'3�S>�4HVZ�d��gYQ�H�͸7"������T�)$�튦�rx|�nÈ�^�����N�at�Ƨ"a�������k9*/+�lcs���3���s�����%E��3�S�F�#�c*��k��Y}rk`�X-G�IJԒH8,tD�b���t���&	��0 Q�&h�/tT���Z��)����M,a�;@� 8�,C[<�/� h�d���rKv��dVs�/�޺��:UЄ���Ǩ�;�䡭E��
 �9��H�����X�n3k:��*��P�[���џ۪��V?3�<A\�ĭ��9C�6L�D�۩���~{CX�摬�\���qk�x��:׬*�f|�F�������
�N|;) W^+���@���@+�k���q
����yӴ��c�l�P��!�vp� �{l�L�J�y�}X�b���:�#(u�X��2�BNIX��Sq	!�����d�z�z����;>(Y%�E��t1������[����n��+�p��gӢ{{�=W�nI�����J(�(�\�Hٸ�.��DK��EqF���k�
�*`��/F�,��]���=�o��0#}��3�cW*�*���6;�F�uw�ȓik�~6�fz<��k���v�/�n�D�ZOؼ��du�i�-0Q>�- �]
x[u6uz���.R��q������$\Fq�,�y�xz��=�Q����N���������1�]�oh�m�I��`��<xK����^��e�/���u��Am3e�w��`�!�Z���GV�:���`�jf�\<h�D����Ǘ�����`DFa7�̘�Z�yɮ��$e��� 4�Uĵ�S�B�w� s=��m1%_�|�qx��;�'"�[p��T�VK�J-��G�`F2۷�M]qE��� G�;z_��6t�.���1˫�.���z��)aD��t5:�41	tEtPDӋ[ԏ�ኰ��N
'����N�1�T����J��e�"ϛ�]A�|nϾ�����`�DLyL�'c��xɕ���8� Ɂ)��)��&n+�vpU!��&�Ϭ��?a��i�yS����H5ϱ�גe-��R�6l��u�p�cs{2��բA�򀻷�#b��,:r���L�p���Zk�@OT�j'+���������>Df���2�W~R
BB��2��Sf�'�Tح<]g��5}��W�&��H��������w`��9s��[*ɛ�o�K�dR[�9Ο~��Z�� :%#Ҹ�B1�X�4B��������f���J�c[erN-t���z��[�43�����lv�|!t��G���������Fa9+���#��2�����"�O-Z�ֆ��珦v�%tZ���C���X��ڵ���RI���j����l�ԽQ��g��{2�Z�7���M��� ���\/��rP�PfV� Rሧ2Պ���
�D
+u����������d�U,ax��Sy����ѝ-r����M��!�n،�XJ���+�M�ua��@�/k�T�� �ȇgT�#m��3�)�@���!�y�w��n�X��N0�F�!k̺}6���x�ؼԼ�N����~p���3pzิ(Ul�*��鰹U8��+g�qy"2��8"���������8k`���!���(|R�g�Վ���qj4.���'@=b����T�*e��V��K(��d��p(]�3��&34���](t���k.7���kþ$/�K$�pNAk�_�����y!���>�B�p4�|��-Xh�$ �=�C���U0��9�� "7�x4"/̦�#�^��g1�D�A��:N���;�V�ԛ}��>��u����Q,O�@�5Y�;*�]���ۙ���/��[N�f7� �:"3Ct�Ș�|+J����hW,�FU��џN���[Л���G�2w4��^� B։�a*���e���<��_��#����ѷ���&+V ���ǌq������[�'�C��E�E�r�6AWf|��a��y@�����xL��>�ix�r&�x>�[c JU���S��«x�.��Cm	@8�B�V(�-��ٍH��T��W�/q@�E �z��E��R�Ϝ�'$x�eĭɺ��z����a�L\��c��n��1���;m��r��{#���B-���is#9ӄ��N��4T+]�lZ��u$.`��P�P@R*��WΎl�p,l�l��$����e�2���U��@�i�R�9��+�@4��JV:Y	�8�`�
�)�.fFqn=w�%�}ET;��0p�ԩ�]d�rw�Hr��\�Rȓ2K{�{Q�H�AH��/�w���ͳ+m�u�pj_i�G�ƚ%�!��yj�$|EH�{IU�τܑ�-ψ��`����y@���7�IVGY��,nw~���zOU�{z]����!}�O���	p�oIR�	l��vx&����OW��f�-��oo���
6,1xB
�pQ��3�c�j�5�vŋO'e�����):LPV�fU�^���h�ߵ��S[�0�������ɖ���u�Pz=]����7��n�ql�p��8��2��p
1L�gd��O��A`��Ni.9e	�Y�
[�+���(L��������IkF,�*��w�h��Zl�
U�!*����ac��kJ=�^*#D��DG0�dR]���y1�v���2'T�fy��_~O����g���e���v֤cv2����!#�I��)�>�MON�K\e���\�+p;�Am&Ȉ���6�����f�x0�y�*V����R����T��B��4���<:�%[xy�⏯6�|p奱!� �s����<��#s6���2]�Ի{�Mz\�l5Q��6-��(N��8����{�Q�ggQˉ��R �ݠ�TQj��Lm�VK�̨ۜF��0�%�,Ưh#;bg����H��\4���=���Pm�I�T}	���Ze��v��J�d���,������Gc��I?n��#y�C.Yb#�L�Y�3�,J���v�P���:7��7��'ə4��^#�
�i^$����f�C��!����m+�7ü�����5n���$KbQ��,�"%����^�Ȓ��3��������j��Vٱg�^��!U�_�*� X�s{R�m�#f�e*���A�:S��7��«��T�i����LDGV�U#�d��{ëw%8[�w�@�1��W z_��[����vG�A��A �}�̊���(B$H��&�1v �j����̀:b�����f�`�H^ӫ�ӚĖ��pQR3d1���s�]��sr�"���[!
*J�����Q L�<����hr8p����Kx��O`�8�1;g��Q�E��n,��B1Ÿ@պ����l�KB)&��؂;��J�é��1��x���yL��z����O�^Q��.z�������nad���3�/�I�>���T�����[}�]�h�6�"{���w>��;��<@X��%u�k��*�|~W���gU�[�����H�n���>\>4Y�_8c8P����16�d�_����1�D	K�d���LOdҘ��y���������WފXVV�L�UP��k���2�'������с�4�>rUxɛ�W��ԋ�4�86jÓ�)F@�K�M6��h�I��p�U�'�[%��\�ط U%!��X����t��:��D���%bކ��9�H3z	R�r�Ҷ��F]EΔ����Z�bɰ���L���a�YW��.u��ю룯r�mc+\�>WP���P�e�w��6DLr�>��Rco�Ac�|^*[�4���ł�N�����iUS�ϟ݊+��ɮ>���9^�"/���������� uA��y�[øJ�X�>FUG��/���eU��|u��f0p�C�^R���2��L=�_L�NځIӳKf�f�B	�˵���%���as�΂߿�ZL�[�%`B���$F�7��<k5���45�s���>��)��dF�"��kxb5�&�
[w��y!E[O��	����%vC��bg�f⎽٤<l�|q�5�q*�Sg)����=\�k�#Pe���Y�*c`a�)�'~�D΂��'Ӵ��$���Տ�,�����$a4�p�uAO�SX�vX�uM�&�h�Ĩ�����9���AKmŦ��1�8���Y�4�������6b4m�.�����X��X��0���Ľj����SC_ϸ�>;�ϔ�)������_aB EO���tN��8��������E"i�v���Q�/O�8p�0�q!B�N)J�jF�5��aҁ5�r9M�j
���p!�yj���F�,���h�y�p���!a)��ׂ�i�.H�R�;��1jqRLj	xi�ms=�����+Rh���D�BO<(ХV��c�p�e��`�׳�5~�%&�"v��6Z�VMҸ�<?��=���6;"J�@ 5��u��qJ��w�������m'�|��p�cL#�Żp�m�q)��֜���CE����T��)^�x�=*�����S�95)�����ڂ{w}L}�~X�L�l�Y{1��P�B�r�m���:��<2*��ql��j�m��N�����<����E�jL���/;A`�X�;����&s�ux��2���d����؄��� ~G�%a��{����x�摘��L��K��&���"�J�ºĀ�xX�$���ٵke�Ft��<�����9_�=!%�k�����V(�,/S�;����hl Qi���=YܮE��-�����݆����*W%��C�P��7n&Ys�(�xr䠝̇jxW�+�E,P�gBcx
M+�h�Cɔ9f���S����|�<m<T�9=1-� ���Y ���k�`�dL�(��Y�����.W��}���y��L��WL�u&;���+�>|�IUlN���e�������UO�h�ztԠ���#���,�VK,Mc���-[������\����`��dY%�%��aϛy���<a|5�O���M��Ա���F�)*�?G�[o�z;a��<�:�;����I\�j��z9�n&&�{E��b�0s<�IEۻ�'bg&gu���O3J�͢���@����t훫�F�o�szҘ@+ǐGZ�ng��1|�*$Q��,5}��¨��U���_��A�EAo���o-�8`����Gp�1�'}Rg%��B�؄�r"���6�#��)���r8�tt3�Rb�8�ĉ���V�ܛQ�Ȟ���>�����O�f\����~�����.���|�R�R�N�ٔp�4.t�y�sȡ�C�QX���9aa�[�$S���-��l>o����3�����a�&�$�&j��)�����N���I+��Մɇ�����`(��NK.D&	�o��}f���3�z
����;�=ȟ��֤1���z B8�9E���������X��x�+�'��c�kn�ѵ�8 ��B��;Q40�tY<nsSG1|ygz��C\��f�r��g��Fq������t��w�t�s~~�p+����\�y�Tr~��U�tYH��rۨ���.��'D��Xޙ	�&N�T��m�Z�We���]]>�w�� �=k����E�_L_��y�e3����x@�~ �3���� ��A��06_A��u�:�F����z�L�r���A��

�]��Dx��.�^�v^�rE��.��+�o�{�j��u޲隒uEx�>�oW���O(��
�,u>v���WtbG��P8�(�j2l:�Mj�ub�����t�4i��D�}���<�n%_��"/�K�<k��y
{ 挵1��K�Uf�<�ʎ����fv0CK'~Lm_�0��d
�ZQ�ub��$xR�i.��a��S��س ���r!�~�pc�����ۖA��}�(��
mJ����ܢ�����(���
��4%�}�ΗsJ��0ԫ�\�$6��?>���;4u���ΐ�ё�V���}�a�h:
zy��Io�߻<U�����L;�R����o��P�,^?�o����ל�J6���� o�F���u�����>��*������F0�M�	X��,bfTěC��c8_�
�r��&���Q��3DVYhQd�-���䴉�m�wGEғ�����-ؠ��?�3���~h MT"��Q<]�Bf~ w/��_jl䒾�r�!t��\���\�`�����
��ua��x�����߂-^�D5oP0���Z��2h�p4ĩ��u,�l.}��u�n.z�x+w4�_@ʑ�6,��y�Q�tS{����i��hT������w|���c��J�w��lS�w��eN�G�z�K��|g����k����[���۔��Jl�f�o�˳��Ջ�@J�@��س�	rY9)E��El��d���%��1����-G����54�����znȌhs���t�'Rv@H��p���KOt3�)H�W����Ʀ�6[nHg;���T��x���\!>��x*j�����3�� �S7�Ή6wK�������@ �Ξ��s^������r�:�)������%��[��#�f�x������=G���!�c����{�OZkD�1,�Bӛ�6 eq�=0�'-RR*�cq��(@G�m�.��c���q2�,�x8�O'������4j�v	a³-/@��SH�Uk�����4/5��wa�˼E����Χ�lX�ncE���rWNR+�I6z�S��G&㧎V:M�Eo64N5i��y'��*f��߫J�O+��.��n��wR�('�E�{ /�~E��!�qY&Uo�QO$��/*kvVx��_A[s��=`&w�I������q`S~�d�pI�SF�R�1z��磗J��.Y����}D�U�K��R�q�՚����Z�;ѹ�.�S�B�R���S<�a6Q~p�O�&�i�D��+�<�l8۹c��!��d��cO�tMP��+�d#o��ؙ�rA������+Qi�)����Z;�XZd��A�ۭ]@D%[�=$[��ll�Pb��`IQ�"S��2��pnv
�9���04�A,�Tac;�q�Jl;��Ý�eN	�dg�:�~�-�n\�;@W1�afufv�8������'�?U{��M��|�ޫ�/��"�m�`����?:0�s5'�קS�ܠ�XVkGWL�ܥ�G� h��.�	�	�gC�����fck}�r�^�>8�6�,�a��iNȼ�+{!�Ԫ�q
b�8J.X��	m��&߄>�w5�k���\0�R��UX�_dd�"���馑�ϊ�[���{)�pp�g{�H���4u�w�8ëb;��|۲�s�Yg��~����t��T}�D������ԂĊ�}����T(��WR���8\9�����,�7D1����ϗn���$�<��?5��5�ݶ|��F�xu�QbW�S�*?ςiD����/"�	��3ef���R��)g|��l��Utn�f~2ОBz^��o�~u��O5ӏ�+��奤����!!�+���Up�&��Ɲi�n�ƾ�b�^��4��H5<%uX�o���šD��K��_�Z_�y�(s�O{!��,��{gTVc�^J�1�f�;hB�:����	����G1h0R#T04���/~����#e��|A:�,�T]���3Q�v�K�Vo�n��FL�3��*%o\M~8�Z�k�~��E<+���=�e-kp��o髮�ylw���a5��8��D�ˀ.И�*4E�7)�P�&�-C��w_l�������U� HУnK�:Wr2ph1��^׽R-D�YpW�b� B��G�o�qo�����S�UG�v�z-���f	SBg�H^���4�LM;t�9`�
9�}h-�\� .plw�4F��U�,x��Q�Z6�"*�&�t� n��[|53����̧#���V�A3WdՈ]�a-��a�������1���Zdt��J�
 r-_\%Li}�P������5�Զoa>��� � 6k��4�׋��a��~��6c��s�q>6gV��/Ź� ���1�F~��8��g����8���W�l*���2^�2ǳM����>-4�
')��j���rQ\�t�X	c��Uh�1��£���t,��<|����6k�D�R{"��fT�8s�ې��8'��Oޱ�Fr�I0�۵J�-dG�+9��"��w�#��+����,G4>�4F8�-�@n[���˭�+~��^g���K��H̟����/v���Kڛ?���i��� :��񰦹p��<����T7�ts3d	b;��"�u =ލ��[Z��? �XwY�L��}�!a�=��IR��i\�Hr �ڻ?�J�R��P�A�h�t�ݥ��q%��o5��G��H�:�a�� �j` Ǹp�ƛ�=�C]e�����uG&�\�Ol'ƍ'=������Q?��:�cv�ndwA9=[1�O���'�ol4iM'�3A���5������q�B۹_;̐hz���������ƼO�e�r�f��,�)������i�$-Ş�ឺˊM��N����ڤ�f�Ft���l7f��;������z��_�9���)���/��`�R�@L��V�N)�ҳ*��)�����Oc���?���u��G xc;�B��P���
k�W�u�5�-R	e�|�h*�)�*�'���V �VQi����<yf�?s⟕�ybq��p��]6M�u�KʶJx����Y2�-e=�1Z�4�j�3�{�l����s+*�Qn�
��"��a�dN�0�	�zAF�Zc��BGZ燎w>�#�w��O�N\/�5��Ot���x���h۶f�+��A 1J�>�Lh�Z#{2��T�Rx]��il�t��Q�v��`���;5�\���;�Ӂ��Z���e�݋ؘ$�G����˞@�3�u���E��}%�Dצ:��,��Z�ؕ-�M�+��,7�%�����,i�в���s�oC���t��ev��sE�����f9'����Zx�'��	���;���<a����*¬��f�����n\�%� �5�Y8]A+�c>��kH�<���6(Ӵc^��'�����fKb�0,{�(�V���!x��o�q�Z�f(:�Q��;?�/ߠ���_}�ŀ���:�� �g�s���4�^w����5U���f�BL�а�����4�>�e{���x��������w�������:�A�)�:EK��̆���3TwM5����_�܀%�k��K�cI^�=v-�0#k�!'�:Q��QK�l�}5��/�ʘ��,�pt��c�
�Rփ�g�m>�r�r�:�iCz&�;�����[��x�u�3��؊�!:eƗa�Ң�3Q(�ő��?Z'�1떪M})�1P��9��~���\R7�����#xn�V�+�H��.���2c��Y��q�!�1j����.����L��_ġxR�Έ,]ot���������iɦ��#�����^�[.��	#(V��NT/i�p؂�����ݾ] >�}S�Oo�A꽸����e�lO!��FP�z���`��͈l쓰>����z�O��>�3�������̶�@�1�$ս��JegE��Yʼ��\	���,I/ι��Ψl��Ӑ�/�ߙO&�x�u�0QkD���t����Oe��-)2=$�7Ddn�����&z�����u:��-Ի���dP�`�u�q���p��[�+P�1��P�%�B�|�ݥo�wj��G.�3{Z�.G!-���?�8�}x����[p�+W���͛�ʪ!�>�b��4��iCs��}
.e�+���!5 ��0��a�noM�ں��G�GH<��w���`ύ�c,h�Yw���=�X�K�� }£�/ٰw��!�OT����"�1a���q貀�SleSN�?�(�XA�n4�#b�ذ%m����!�_fvՆ��pLж��+���>��6�?�L=��g�ށmJ�:�nd����m,I�P��y�<�3�HL�!
��|x֝JcN	�\�@�"ځ���~�\�r:'[�8��g�]��;2����<H�<�c$��=��u��,�o+�E��]`L�4,@�ݽM���t�	�$���
y��+�.��1�K���lf�"k�h.��������"ֲ)���V_;I��/~l���X���xʪ�=|����Ĝi����o[�)������n�#����e��18�{�ِ�P�<����̩˰�R��m�w�9"(�S��
����ؗ�
#�H0V�5d��aҷi�0Y�8/�$�.14�����L���$h�G�Ut�EO�QE����dB�ʙW��^ؘ�'0x�=:q���2��J�,�����Ƚ��������Q�����M�	Jy�g!N�6�H�}!�A.H> �@+td�
��.�M���/�v�xiJa߀�5��A�N��R��<7�w��S]��,t�*\/$��1��3���4��&�+n�ȋӥh@��7��y�V�R�`U�&�0����rY���K9hh^q� �|Fej(�r��x��*��Z�9u�r��y�LB����9��\4+�@	��i���;>�?2�����EO�C�lӲs��gA��z�ᯙ	��M<����6�MJ�v��ٳ�9]}��(�J�؍�KFV
��.~�:
R���=��r�{,����1�(����:��3_���ZM��ܘ��._I·���͞��wJ��V�S����U_�`F������_S=s3n(K�<��Y�:̒i��񋙗�Dig�DM���-�����U���ll�c]0��u�m��[���0fMƀ(P��7�p-KrTщEk&��ۦ��r>7�Qd*�R��Eg)���c��
�����2�\Y��(�x<���Sy�~�Eb��:֡�����
v�����������&y3[�d"W�����w���);��a�ȸO��昆m�z�Ta��vZJ�z�	�� r)B߹��-R}h,��Sn�߀l,�"R�x�9�$����~S?����=rW���ފ�DPs/��I��hf+N$O��$�� �C�֨H[�M7�-P��Q�N���΁�(�uuv�X�O�S� W����t̘Gn��/�^�#�kp%LkV��V�k�97���R���������B˚��/&O6~���8�TIq�%���f�"���QH)]"�1��h�g>}z�\5t,�%�Ϣ�>^�`���L���˺�%���L��x�
|L(�V?�� 5�9��];)�c������)�������&�r���j.U=T�g"/Ԍ����;�����5{ɇ�����&�*S+�Ҋ5�j�"\��n�>gT�,Gi�����]�d.jVL�zF��-�55wF�q�µd%��J��{	�1`y*�5g�c�α�П|�c�$�fU4ڡ�ؑ��^��������=I�Ά�uh02h�W���XC_�e� e���-�a f ���DE�����m���q��k0ڶN�v�Q��(�pl0@�K���j3�˨�eW���j����%�D�� n��B���n\��.C�S���Kǉ��S������|x#���y�%C<z�P��Q�OVG�Y� �/���T"��eW e�MOͺ�3Q��׀E�m���a6s܃,^(ָ=��ME�C��A�� �����o[��Yk1+���L������8C�8�i�u������Hod�t0i$?��Q�_��
kF��p^Y�Z4�:���#��1Q����� ���u+���}f;2Xz�5H�G��x*��j5�wg�U�GW@��a<�	e��Vτ$hp[�U% �YV�+rt�e�_�Ez�O�K(˘�tuN�q�j����Xx�1کF?�M�Ҫ���0KB�Թ�/���"|8��<>�W�X�s����Z�d�Z�,j��s2ҁ�&�~��0UH-�V�f�^ͱN$�'��C2��$�����
ET/��p��H�~m����mX�b��Rh���@ET3�.!zʕ�jY\�i�r��Vqe& l��
 D�|$��5Gb��/�΁�>B>"p�x	�vH � �7���!Ի^�>�s�O�ܲ����:V���#yD���6I^��@(M3	�q��n��X8�S����J�`F�uU���ˊ�2�LF%VA�y�o����|��=�(���G;�����B�$�ރ��X]ouO�8E�X8���q-xM����w��)vcB(�d�0��:��4)�>7����<� �>_J���Gݥ�39��<�W<.1#�����&�x���i3������i��$�f�w��avU��|����v���χ�0�3qg��X'ީ���>�9��B<x����{�m��fpX��a�V&�<&T�A�.ZL�&<����U��ܔ�K��#�1��D�Z&�S}�E��Z�-A�Ń���:�_����>xK��X�k/?|N>P�;*)���H��w;�^��	!]C/hҾ��v�F3EL�݌u��bڱG0CK�%�Ii��)���su�9h���/z����Y��]&�ʴ}V�Z��!����E<ւ ��HC� ��fG�������lt{��"��|Ӫw��#�Y�d�^�/�1���S���;&OB��|&�u٬���*�GŨ��u\�W����*Ʊm�{~�����|kr0�n.t_�0 K:ا��Kڀ{�m:4�����[��En��h܋R�bP~Z�[��ѐeg�"�Rq��Il���Ml�@��|�vM���+I��C��Q�cϚ�u9��H��m��*����Xj��ѶI]���S!>�r:ɫn79�ˈ�G��K0�Da��$��%/ģ�9Z���*1ƚƘΠz�X�dO!|4���\�5�U{Q��Q�w��O�LX�!�������xL���\[�̠]�'5�I4�rkB�e��/t��}��T���2jpu{�E������f_�<>)��U��o����f�y����\�߰y-v;�7�j���|�p��e(.�o��2Ņ�����\�6+�K����@ᇝB���%�B�Х�
�ҁ}m�[ЁZ�����X�N}A@3��n���Sn�Ӣ)�`�`d'���QЅ�8���`���[C�O�r#�Wo۸1�M<V^L�ֵ�té�ie3Koo�z�!��N���PO�F�1�d44~
��}��3d�S�Z�W9g��!?�^����o���I�A"wD��e����ߝ��v�E7Ѧv�V��y,�̞��5��&�7~BG_)b�x`�*I�D���>b�Bj�D�#e��͡�Kp"��@a�
ȔD��1��q,�%�!<.;n_V1�����\LU�����j�Ma�d�S|%�±���u��dLcGV��^�s���mp�mO%PNn�A/���ӉI�����M�*y���f���B�U��_X�f���Hi��Y=N� ��`�l}�C�o#�)�v�E��I��N��4@�e/�I�ϼP��:�m.��^֓�e�^4䌯��
�B��܃�ȣ]y�Sr���j0@�F��K<Y��n�)��=Yۍ\��>w�}����*e�w��D ��T������[�cqWi��8� �$9|��T"�W�$�0�'���W��)�sW��X���%�d	+e�^TM��>hݛ���m��w����Y��afZ�K�J7|�2una�ʓ�>��� ɯ�t��ѱ��C�g=�c�_;�q�R�(q�bc��">6�	G�@�� ߥWA_+�͔�Tl=�s�>�
�8-�g�� M��awH,�;
�u��T$��鑪�8�.��϶��M�x�4�����Z%��Y��p�.��fV�ĺ��l&Rs �G�Q�_"�8rw�B��H���N���hP�ۨ}#�����5�#F��4�mه�ik�ġ�$�K���8®�*�ԾJ7W��pi\:������4�����B�ߍ׌�K�z%��}�Af�S��!|5���5f�hT��հ}�P�hA�:�=;�B�
�1z`gB���4#E"l��8�V.{Ĥ!զ�����������XK�u�q���~�����kA헩�GX�&u)�D�����ט:O_�D�T��c��Н��S�mJ�K	�[���˪��8��z*NЅm�?�aJgo�i=0���$+
�����/L���{�P)�~_�p,f.�/�p�҆	VҚ)fB��%�U���V��oz�3�f�t0+SY)�t�@0�Z���P!���Sڈ(�p�!� sN��]��Q��.}�X��q�q���� �*��i}-?hñf���A16�e�c���]�؝�\ah���	�
���j�:[�z���XPa�[9q��}w���M&�&�v7�:cj���&�-y���,}�=����
�����#C��|������yr5~3P��Q�6�Ӟ�{4��S��jL�/1�A
K$\h33Iu�14V1���B#�s���1�9٤|Q�gB�kB�Cr�YZa�DL�(�Sd����u�h�S"xG]i�?y4+Z@��NÐ+��!X�Yc˷����R{���1���/�t�_k�.�wv�eC36vw?������-���W�+��߻�v)L������*��5��i�pzʑ͙�s��7!|h�r�J���
OL?	G������xg�G��+zb�#T ��`���ͷ�!����g��2��	_l,�S7pH;�1����5P�S69K�*���Ηy�qU-2S]�_��h������e�DL�Z����޻�2	��aʝ�҉����y�}�?t2��8� ���"�{�Z>#� ��O�&ƛ�3��]�o�^�o��:!�|�%ֺ�K7��0,ɍ~��8�8$�͙�b���
��'���Wá�A�^��C��sފ�jn�d8]p����^EW�>�-r-'b�byt�ol���#^�F�q��N'r�{�<������2�yp90�H���*���ў_[c�9.)>���.�ݖu%��w�Rl}�菴�*���sW��U�4w��B�1��i��ӅH����$����r*�n����Hϱ[��0��H\,�>�Ck��aȜ�ˠ��	'[&E�h%�d���7��!{ӓ�'K@o)�0#t�$�08tњ�<V��	��p��?�r���BGi���O�!�	�P��+_�p��4m��Y'�O-��qn���%��M ��'0[[�6�M�p��9	�B���tӂy�]��	^��k&ҡ�Mf�0@k�����֮u�I7����8�P#;���l��uqPĆ@��yV"�eY�l��(�h7��m�_xl�*'kd�T�G6��VQ���,��Sݕ"�<�Y�
a3e��Mes�_�voU"e:b�6��Д���+�ȋ`�5���^&�P_���-A`�]U6�����&\�}�-fW�R`�B�T� $3�n���DhE(|nc\�ɮ��/�:wP�t,�tד���.��sC�%P̀�C�~��1A���%'P�c`�l��ؐ��X���E-$\�T��<���
D�ea������nr�ۼ!���^���(u ���� �����ҫ��������H7�OM�
Nw�h�~�햎p�]?��V�v��g`��g�&��N��ٵ�M����Y�p|�z~�1hq��,}W�`�Uߧ��j�1��')t_]0��t2a-���U�GK[�=��ﻆ�X��)�;'��f��<�D�z���G�;�wS9I��1���؂�*�#��ow� �x�}K2y�@�(x��.b;?o���Ľ�Z�|j���I�(.����N�lk1�� \�KoS��9$�$�'$�ܡ��a��R�`���J�N�㊷�/k(.x��y�����H]c^f����Tw���������z�!<η �Ԕ�˧�j�V˙C�*l��RcRZE?�@t4f`z��x	�p~�~:=��7�]^�d`gr�_��y�EG�VJ��	�zF���W���߻�&��F���q��:�軭1�6�{x3�Zy��V��jৃ�ӆeS���=�z��i�G�DO���7�!P��v�1���Y�3Q")lb޾�d������,�w4���:�ۚA��V�y�ps1n7�@���L��r?C�� ?=�$X?쫆o`��ū�&ߏxؔA[��Hh�q@���,���-&w_yݩN֚�}Ky�j�O�A }!$r=~(���
�<�y��D\2C%-`��<Mrw��J|�RT�e������� �(M�!q2�!����Jv1�y�d������(�_�������Ur������1�]��>X�E��eh��f[:�<�6�*D�,b8֝��[���_%�M��~�����g
���-��p8�G�䪱z�Ӿr�&GP��k�}�kݠ�II=n&��d�/�u�̳f�I�h� ���j�A
�[��
q�iF��c<˚�;�������x��]v\�3R{s����d4�hЛ�g��E{�}X�۲�b��:�m&�����
ch���j�锇�."oVk��؅V�#i��!K_��JfB�͒�}#�*��1'�pZ��(m��~�i� �j�O�M0a��>����񄯑L}��g�'W�j��U�˪hs�`pj�[X�u���������!&f�F�V�ƙ�v��.��\ �s�o%��	��V3���)�6`+�%�,��גL�Χ� 2�kU���`�9�؜������&���[�z�;�����Ҭ��#Ų���V�Ae>ď(�S�Z��u+8w�+V=dO�ؘ�ޚ����'zU`m�!wiB��!?��Z�O<��⋒q#���Ӫ��l�(�a
�g-��kV�96���E.�����v�*���=rW0�\͍��j�8eg��<���7�v�q�����y?�Z�p	����2�1Gx��[�Q�+X��������ꁔ&�e%�#�����WDplB�5�A�	�T��*��tR?i�@�rџF��k�+�0�0Zʔ�WC���1���F"dn�b���3O:ll�xW�b����#�*����|��%�:ͣ>��uj�eh�icn��2W���Qp�Y�X��L6?rD�|Ŵ��SN9�a(��K��XM/@j��x�|�5���4{ғ6t��
�EN��+|O��΢�PR�Wt�yP�
0����co��FVi�Z�`U��1/��������)�=�
�	:��z�C^�W�±�<ET%݈?��������V�Z<�쓋:\�{[]�e���d$��̳ wl���{P�]l('��|KF��&�@+5��L플l߭���hM�_b[.�=O��,>�#�ͷ5�P�9oɿr�}�-ug�O�iS!�e�Ye����,�
��l��ԥ��0W�=��1�f=���~~'|@ՠ��|�񕃗�4^�^��1�rM�z��I�+��M����Z�h�Q+�L{#��UdNC�3��E�'�2�����N]|��K�y5�=%���(�qo��*�Q�����p�Ar�6��G�y�1C��[�R� Q��N�S1��IӛqX�%���R�����K�O�q��a�-s��_�X]Ћd��9����h��t�˫����"�f��/bJ�8�A2���$+�K�%��	V�?xZW�?Bɛ�j�I��7:2�@�!��V.���s%�� kme��)<E0��I`��?HsE��߭;�F������F���_��?o�'��?�iu�,�CBJ�����2:-V�H'}uSF��EZI}kȊrz[	߲���p!^�kC��f��d���SAc�C��#��ʩ��u���t>�&�>
��"�"c�Z�6�O�Kn���w�*H���t�9Oˍ�	��jd���r�]�X��r1|�����28!za��B�g�p� ���S*�~ԗM���e&�u4���4����c_`v���p
�y�}x�!L���k���8e�������k�r�׭ajf��M§��m�r�ǿ��mz�O`҂Q��s�������{aG��Td��[aȴ��%����94�!��F�GlcmBb�=�%�'���yAq�2�z������^i�u���]��T���=?.W!_sfa�	/X�uu�	K��[�p���\A��}h��n���Kf�DHq)�*�2��>���t �}������󑡽N�?2����s���`�-�X1��T_ ny|�����kZ���>������idPb��,�R��|Y����|��_�A^���F�uf��M_@F��6� 2����/؅��<T�R-�*�.Q�#ؤH��	]�7����Z=[���?�ۊ�𼡄�f�<�����V�f�n�9�oc���.o���(�)H�'9�
�g�=1
w[�.�Q�Z.�@�w�>�-&�%W������?uP����kǯ�wxW7R-<�af��f´���1����q�0^e"���1�w�P&6a�Ә䃝aМ�O����M%�i9�p�����2����P*�J����908Q\DM*�F��9R�2d6��إ���:/�:h���l_GK��}`B��9t�5���2��J"{H�{�e����hOH�o�n�y��ARcAF�����:�wҩ��: I��a���oaQ].�cTf�,�	!���mG�I���<Ro������&�b_S6&h�!�������8O����3Ԣ��ieb|�p 6���2U|�0pv7	��y0�|
� 81QD.�آJ��,eH����o�bD���Q®��#� 5��2'��D�����
�v�`c���[\����_�
^2w>j8�2h	Va8�y�܌�R#i!�N��N�pr�Eg��[3���ƫI�I�;����@h�-����0�57m���u-{րkiJ�!��ۗ�]�3�Y���]���2�=���SEC�ҭ�	�q��;��?����rG�9��Ya�+�B�k}۰[�(���ǳ��<O)<D�n�n�.���y�S��k�e��j?�;~O:'�<i[���k���r�xl@l���K����O9	k�W宪}'�gr�D�ƨ�y�=�|���O��e��/�V��������c;̄�붶i�?D�Q�!�?y���W��j�_u�]��%},����&0߂m�[T�ȫ*mO��(�Da�n�m����<q-���I)�#v,pu\��;��kÖ��t�z%F��L��ǥ�Y�C	KfW��2�q�r�#6n�t�ubK+0�.��1Zh���V�p �k|��f���,��"�̝��7	��'��ٚ��z�3��V�`G���9u���w+�������X�4�1V3�.7΃C�R�����T/w�6S��_US�%xQ-3G�7��X�&����6o�A���~w���L[�N?5�Sp~���{�ɐ�ҡ�f`I�7V)3�Ü�2���^��랠}�C�|��ǲ7��&�X�j���L�?�:����,��C��dM���)F�l��_�1DJ�$��7�<��R����-��$�{�bg�DX��*w���8t���~	�@�7��V��ur�Y̝��ٜї�'>^he�ކ"���q�7[kT��w°�����OT'L�p��ͽ�m��dj^AR�O�ч�Q孛��;���Gw��x՟�V9	�
^���`^��2K�C��L��34`�0����`���a�9pU=^�Qݱu�:���;��s�u��@��x���N���Q@��K���sn�IBظ?�^L�^��Aa>0K����75 E7�xy*�|^[C(6�<��$�A�B��Mՠ��a�ZۊIB�ßM>���[��pr�1%̢����.-�0ֲ����xs����L��6@�l��k��~�Y�h�]��Z=��g�됔ϹgV��-�3_�ص.�H���xM��K�^���U�3�zQ�U7�C���#�m.U�S1r��\b��Ϊ(�)�W������B����A�ex�]���1�����(�=9ah�T?�C�ecD��^�!D�;�$��h�St8�#��К�d{^c�:�6�����[�`!
C�Sv�`���C�L����`-��ܦ��A��8=�����2:5b
8l��:���Ī�z�W��� *���n���Ќ��p�HŚ�w��.j���P���̀ ̀�P_C�[��rmz ���Y�(�J~k�B�8x	i���b�l�I�|�]~'��9m��J��-E�2M<"��B�hH,�<�t��^����$t���?�¾��K)Yg셖�kI�dA<����W��6�j Ʋ�y�AE�%;��M4���=���(�9�N�c��R�8��N����4�T��$(+!�ÐO�ϰ@�O��0%�o��_���t���.��.X��}��f�R�~�N;uM7��d$(�`P���X��,ǍU�h%�ݫ����m�U&̯�-�:��:��#��1%�w!��y4I�*� M/D�`��j���
��*������s��58�]5>�e����V�ה����j���ϡ�����!��/�'�<�Xzn�ߘ�Td9^��p�'�Z��y�NέD��)�f�I=_���[~������h��t{���jJ�`�:(����%b�x�2���W���� ����˦x�@�'�<<����'�W��n�����D�}[�قs����G ��aJ���U/�#B�
�K8:�߫�\���K��`��u�����uYQW�@���ӃGZ����Ik�i⠾]���$�׀�(���8�,Ou�9S���8�'P� c�p��������� !xc�o�?��q�!@��*M�F����؛�|)��X�Cˇs�A(R�iX<F\V�����Z��,��N�,�򋓲�dQ��d)1K����ݛ�d�`I��tp"�?��h$m�NAڽnZ߸"�l�7�� ��H���m�Qi�	���c��� �#�KoKZk�̢֬Q��kW�]��C��MMI�зP��簡������8&�S���x�0TG����Y:��~
hG;��Y��_�0z��:����$����
�<%��t!�}p և�#Jw���j�4���-�Oӧ�_U�|��-3����W%��b���_' �A,�����iR�^r{���H��|����N�S�j�f	G9E�� �D�$����(���tֵ���}h%6��#S�˩)0����!'�\AM��J��fY����2��݁sӼ�_B>�v��F9��`&J��� ��q����;�$������	�SVS�	�0�)�=���"�[�x�1��
b��'�Õ��kA�z�� ����*����K<2����J�P���+�pN6u�q
���!�i&�4ư�u�Z�!g�[�7��T]Q�yxE��Pw'�S�h�@hss��i�I5�Z��E#�&E��c��Hߏ� s2+���������9%�c�A��Veg���*1VV�sQw$/�U>��¥JY��Տ��9rs3����4Cq7�F?���7�­�B`#XXg?^�W�T5��&)Dt_o� .�>lI)�j�݊�ƓJ��B�[�-�yԎ����Z�� ���N��� "�@*�9�`{����>^���)��kC�5d�jB���KH��P��x~g��B@_�`I8���P=�C��Yf���
�\�|
�v�lD3�Y#�ʊPg���,h�e՗H�ׯק�̦Z��](-E���7Ut̉l]�ρϋK��A>�Յ�����Ur�LiJɘbE��d��C�+6C�n�>��|!DG��#�^󩐫t�I���3-1��@�E7�r��)�$z;�)(��d�k��Kسͷ"^eԆ��L�S�y�L
�	s+�~~my��4���tUNq�7d��c�^���Cy�U�2B��^T���{�˟a����yW#[�7�v��P�4E���
^M`o5�-@� ��pw{���r��T�>'���9_U� #+�XT���O2���@3������j���%'k�����A"x��K[s{��V���/����Mr���<D8�,B��
xc�;���P�c=j����Aw8�k�ý��!		MU�Q1�Sw/ߤ�E�by~�R����Q>=��`C�'��R�dдn��gK��WZ�u ����\�i�����C'xD	A8l�Z3�N7�����^�dny~���k?"�!�4���p<��f����)����� ���*��pF����G���2P۝z�6���4-�ʗo��\��0�|Q�����y�bǰN?�ʅ��N*����y�P��G��$���\0%C���PJ����am���rů��n���d�+��g){l�Y�%���=G�.���*��a�rgcW�qE�r|��ڇEx���g��Z��3��?SF���z��H��K 嵁ժ�<�z(��]��J�?Ǡ:��7U8�%�ě	�i� �5;�
����!+�'�P�q'�o %y�(b9���E@��Hk���i8�,pI"oV�y�o�"̓.�4�4��{{;��Ҏ�[�<N_Iց�K���}P6���abX�@D��F�C9r���j��PVv*�٨�/��tlt���#w &u�C�ca�Ν�{�'����g��/��5-�!��X� �h�N�N{�Y�&$Z�䔔�[2�-F`�ߥ^�����d��^������v��:	vr*}�Yn�P k�C���3��G��S�k��e�ep�p�@�%�h���=��<�,5k-���
T��
k��E��.h+��B��;�h�q�K��4W+���C�l�}���g� TV �Y#���إO0�k�:灵f�I��إ�W��.3��(����Ӡz�+]^VޮV�F^!���\ػK_J�W{C��m'!8�o�23�j�E��,��|͝	}��m�C��^S�ey������A ���z��������.gF͍2�qZ���AH*�i�G<�`;�R@lec���(J@@c|�
�0����?\��m}V	ؒ�AJ/02����	s�b�Y���]��<"�"��х"���Zˮ��AH��@lSæ��㬙_�JS[n�g�I����@}���p�/UI	mM��]&@����  �n���&��EH# &-* z�%ƺ���-����;Hn�#|��8e5�ᗸA����h[		�P�>�B u��g|O��wW �[t��sQ�Hӆkcy��l�$ ������*�� _��G�5���š�6�912T]��i�C�b�9���U���]E��|�7[L���YcvP���Ms����m�(���[�mR��p'G�8���̛�(	�1?v�&��:˺}�J�q�ή��а�S�%��ӹ��^�A�C���*1 đ�_J��"��HuA�k��,��� p�M��G5���I���h,�q�H7ɼn�ZWp�8Ȇ\ ��l�oI�D��J��D�/����\����,,@\��2���?��T�@�_��C��|8���]Q#�D����x (i�s�d�'�ы E]l��λD�Em]����V���[�\%�pV%���d�_� �u�wo2GXq4o��zNrp�H`��*�;�+M �e���q�$
�Yr�P��C���;��tAt���2�h�8`It���#4�?���~�kٸ�{����2@�>S0l���F�=�c]n�'�����{���m�����Zf�|��.�G`�L*�������7-���"d3�K����D�6,ʺ�(;�4�~��9����1%��c��y�vDl�l�bP����A��^A�D���0�,�yu=H{�_��R����M$�^E����ih٭{G�Jͮχ��V��6��Yz���%��ڳ�s/�M��z���h͙gb���!�U%�"	G�=�ꤩ���+���������ht���EZ"�L�<p���z+�4 �~P29Xg��yL3�L��TЎ��S1�/���<��C�C��7���FB�Ր�a��C���s�q���~k��J����Ex��]mʀ(���c����m�����}&d�'j$9VDq�� ��z��2D�W��ZߥL-����Z�� �$�{�,������.�)�#���I5W��ߩYۧ-�5�Ϥ�k3b�-�ڹ�8�Y(��gsp�mj�	�тb���]LN�o�|^g|ѳ�2
E:�2P��=q�+H���O�o�Uw�(��<��]]W�ͮ�T�p߿�����AKþI7��V��U\��R��Xȗ��z4�X8i����꾲�Y� S����h��!NK�:�&��ͮm]m/�f#��ݸVq7��~�r3���Hd�wA�&���9�Z�߸��%/��N���Y���������,��B�M	�?.�Oz*��F%�5-�9^�a'D/���"�Լϔ*8�^�����\��"#�CU���j>V��|��g�?�9S:�Ej�Zs� ��B�4�)�o`�?���E6u�p�n*�]���7h2����"D2�)>�{��t6@������p|�&�o�3�\^�+�^�A�=v)j��ث��K�
s܊ڮ�b4�#[��,ᳰv!���HLPv��{��HcI}�N��KO��}_�eG��,�0 ���PzO�FV�P��v�@�h�8	I�f�Y6��;U�
�������{v;�\��K�9OG�]�u�Xѩl1�z.������+��px6��mgT&��N<<�7={j⬅��|���В?�Ao���7�'��ԩ�獲��W�o��7g�9B6�e�%�n��J
-ȓ�#�S�l�t���IO��=�;���3Ȩ(S`w]��9���3;-�6�=$e֨yHߐ�8
!�#&�94�e4��5 ��ܨw���:��SA;�?�/��a�?7W�pV��ا�f�.I��s�Y��L:([�\3��$�^1��{��t����ߕC�;8Y���R+� �Yܿ}a�4��IRM7��)%��+�N���΁���I�@���X�A��4_��xz�,�u�S3陌��'eq�C�YOv�G�ƿ��E�?�C-�p�C�&����ĜX�8�3��v��E㸎���4����B-�KI�����s�R���S�YO���ٸL�f� �V�ܴ\��Ã)��ܪ�r�qx�Q�5����/2�����C��/\-��]NW2�g
V������.����S����`H�����0^At]P4��J�r�e�9Q��O�G���R5�dN�4-���C�o0�22h�;T�J&��'�(�Ҫ�IE�<�("T�p��OB5��uJ��%�*���/y��`Ñ������2R,�e�*�s�ۢ�X6i�f��a�6�5%���nׁ	��z,�l�� -rG���'�[���'E�k�?�B�=A��C�Gd��H��	�Y���02&f��B��ڲ���o���Y'�B����;Ѐ��K��1G0G�:,>*���d����L���$^k{�+�C_F!D������i/�Ca'�߲b!;>p��m�M9��y��*�kg\�	H �P,5L���C�&�����O���
��"	ٻ�~(�+��9I��)Ӌ�Ƃ�l��H�0�?�B�[q^ G\v�����ۍ)p�_4���,!W�/�7��[�=��*>Ŏ�w4����L��ܫ#�۠T�m���sPe0U["�7��7|-5�4=�j��l��{�z�����f���`v�,L�z�ց�\����.I�$��1q���t�B�0���|���
&�<��C1GL|�/L����\�I�
)A������=۸`?ˉU��A4{x}W�r/z~���B[�Y���B�b����l�y�БJͥ����o]t�"��\��  ���C�G!o2m����W�n]AnhD�v�ӹ�-��z]L7� ���)��]�F�A}rEpu�6��K�4�uB���UP�Z�&���������qG�zb�����Fd~np$t8�G�S8���ל�D`q�h�f�]b���$Y1^^A�D�g����kUŜ2���ژ1�bE3�Z"
~��>]C�iE�H-�ډ����i]qBƦ>�z�T�ӹmk�����K+�������:	��r���v�=��e0N<;�U����Y��@J�%@`��H��;�ہ�6��y� �_w��I�a��gC`�$�`��+� �`3��ޓͽ>�vADˋ�ׯ:�Y������ T��I�y�@��e1U��v��g�N��+�>��I�G�i�!�� �w�����k'#�pa���h����۫�B��/�DN�OOMOCfpq� �@t]~Ŝ���_��*e;����z�A~���ld�+��+����_��F|�.��)��f�]u��Q�ɗy��� �������t#�"3�o���e�9s�ĉ��VZh��{��q�_��'�>c�]a��7�^�T�����K����\�*�I*ۋ�Kx#���2�5
]S��nF�څ��� W L�1�=AG�*I���\T��[�&_kF1B=q��\��4!
-6eG^��jv��,�\���D�fFjL1NԵH@2K�����[nYћ�~$�C�߃�,�q<�����K�]�ؤ�Gz60�D�N!��i�``\�Cj��ZY�%'\J��U�.�o�D;슟��%�i���7SLP�z!�[��sl��Wj��� <S^��w�0D@��s�$W|-s4��>�3��ڏ�l!�[_26ʕ��mю��z�22	�P�jMW6��Z�`N�l��-�FK+�J���m��,|BdF�%��Qb4�!�
�g��ތ���� �0��퍣Zk��lZL陑����"dQ v��
�� ENY�nB[ �ڕS�z_�����ݓ���SSY3J�Y��Q��aF��"=��an�5�V�@��ǈ�1��a*Q��������r�/8�mJ<�"	�z�G�h-�� �[�wQIA�wq�?�X7�33z�'>1����l6g683LM�	��TM=�z+*<������D�{$��nҎ�ɮ졋Ou�Q���c(�ceҫyU}HO<
o���<�?hH|,f�S3�����;Wp��j�P�~C�o�`�F��ڄ��m������������v��ֳ�
���6fUxu�ݷ�g.o��z�������xXZ��������K��F�M�4&��k��`Ҹr{�{UL�����7�Om���~�����M�Z n?�^%Dwv�q�Y���+���Q̽8V�[$Jpr�ܒ�"���1���᭜|d$$ͯ�T@��{�b�ԛ.��N��sj�~�j(֜�!\[M�H�߇`u�k�bs��Vik�/�_�M�����v���0�q�k���X�d��,[r�\��p>%(bƘM@�����;�;}��[��E(��-pe0'�/|��k�n-'?��9,<��0�uP��s�-���f���I1[���d��~ׅ����C������:�,`G���5�[	`����qX`^�{���W�z�UbA5y+���~W�u�ǉ+Q����e��/��g�� ]a��'3��N5�FVě`�U�	h��P�*��lji�uJ�r���0|x{җ�O`:g��CW8Y"Z�c6���S`���j,3vo��N���c���JR����S�%n���_1���5��о��6|}7�>��Y��Dq�gP�����W�f�Ya�6D�+����v6��$�U��hYC��%�-q{f`M��0�����b���e5�wenH�_O={�����pș��w�J�J,���aE�)]��FO0a�:�c�#ٝ� �9�7��q�h��ɗ�%ScH|s��h�GWȧt7��`V�N��^���[v0s��ݗ)o����d
��,e<����ʴ'��9U�Xo���)>B��w���K�+Vj2��`κ���A���6kHN�#4��#�\���S�,�R�b��-��
��b�׺����7�?�nA����H%Cd��PAD822�~�� �-ך#�*K�]��3lѸ�ob�� `�O(	*�F(�����NS��I]�3��A�6/~o+��
۞P�y���:�������M�PO��g�=��Re4g��ċ�&�-[3�����3d���*���(��z��>��޿�U)��O(n�gqtHv�jd�KN����G��o�����1`4s������G�����퍎[��B��p߁���!�L��w�Q��Fm�i��Ч���
0⍢������=�{���6���6\V��>)v�"u8���<����_/�����[:��ǽ��)W���?�n}M�G���y@�inKX#���(��A��q-Jx' }��|䈡~����NM<�/��e"�/�ƐQ�0	�rF	)K�MqA`� ��B���'B��C+���Aq�Y&�yM�N����&5PL��$p�!��
^���i��0ꀸ�y���8�*$1�:;H rU&mX��1�h Q_!���z�����&����]�b4��;�x�jo^��q�#YyӂI*Ό'�0�N���k�K��BD�������{���A.�)s�/��<�aڗ&+�ԔJ�iP��D��0�7@��J�Xܥ��T�$��������3�YjdhsҺ����=�n/��*�X��C�&f�W`�Ό%J�!�e��>���5�����P�wYH������`��"�ʉ�8"�lŊlibmn���FBꍎ��^�����QH+�dW�P�����U�f-Z�/:.Q�$s1^�����ѳ$�/}N����GHQ������z�Iژ 9�.r8!8�d��I ���S<
����9��N~(�V��
�P'Q��n�+�Rw�.K�����w������H��}�;�+{p\@���%�
Ч�0�yv88�θ���܄c9�z�=�٢�U����'ZD��LCq�TV�H �ދ�"���T�
�/�τ� ^�/� i���][*��
�Ƕ
71)��$H"�!Z�����>0U�E30<�0�ψKns�<�y�53�Jw�p'��ɬ��I��8r��W�[/BW�9��W�Z*u�]�>WO���o���N��b�����k�����N��\W��.���"W�n�M)�̼1����C�
J�r5��h�OWl��P_�\Vy �lN"��W�`���i��:%�.2�oO�mV(JPٜ3���s�҈;f�v :I/���n�|���B� ��\�jx[L���s��Y҈U����=�s�m�L�hO�̈��TԌa&o@���իz2���P��d�e`��ȑ	�4@���`d�6~�M�����f�����H$"��M�$p�
�p@lJ��V�1�Ι��J��;s$�X�bE�ۅ>#�9C�[��ʖ�z��'��y;�e�z�D�Msښ���������@��# "�aVԯ�j�*
u*a�\�����Si)��J!�Ŀצ{����x��c0�b�٠魑?���ܦ�N�q?�V���@�A�}N4�H.�v˲��{y�Y�R��y���S2oē"L�z��D��n�k���d}�m���d�h���:�����rH	�^/�R��+�蔂zH!t��,���v��~��dkb���֩����yW�0=��>3t;�Wꁤ�$�����X�[��W��9�/Bzb�J)Y㼉��%WCR�����ȱƜ�R+a6VK)����b�~R���AT����Ԣ�-8e�M�y�aW����
W����6�/�Ŗ�3I���8���
����!��{�=z�����6'F�<�x���+E�ї���ü]�8xI�X��Lulo	�'�#\`�>�u���^f"!v���h֡�,�� �������=�o��%�F!�$J�p��t[^ n���0H��厂��شm���Ň�����kh#�l�	qbqf<@;tq�p�����p�{2~�2D��2�3���4 ���������@��L��X]k���y��.����F������
�"w*�����*�3$��g���Z G$|��>�<s���z�᫖���{me^��A�x_�����)�������L�b������e�W����\��z~<�K9ր7��vk��'?*�S��8q���xɸ�j�6�s�{ MV�k��4�L�i��G�6�љ�r
�z��p��l8;�YgjH�]�y���W�(8s�^c�!�c/�n��=uT�(�sP"3�
�.���[cȦ�N���:��<Ú��Xd�~kD��h
��WR�2�\��$�e-ýYZT֩��Iv�/�f��Q�;S�X�=pa�;!���SAW�E����x�	�je��X&хd6;�'���)G��Y�)��D�6����S�1�!����ӕ�v�x����'+��+D��M�%�m���`[�H���:��� O	8�fNO)�m'�xv1��Cx���6�����y�܂V�7K�,�Ci��Mo��[��j��dD,x~O���5#2�O����N�CڒT?��3˃�4ZR'`<��R�"�6���xQNY����#@�k��	nV�tn�=V�h#t]0�`��R࿄)ʵ9geI|T�^`�~�^�ƲͰ.�m ���z�iA�aTK��`��4�J?&���ᶨ25 J��v�א>M�YS&VS��k��gy"�c�sI�_�TC6
�����^���OC$��6��e�-��cKK �X�דW�z�pEQ��4QY{�>DP���N�z��`�6����]�`oـ#	��[ciL����O�<i�(?���c'�����`�]��Pa�ф$"��c����3��u⽩���ڳ^-���Ⴕ�J��hRv����g�L��)
�O�x���h��V���W��3�;�v��`1�1r��������An�g��#��mvQ�8���U��#Jg�Hh m!��0+� �H0	V���y���+U5��W+O�h�L.ᨐ ����uQ"��!#�1�@����aB���+ ��e�h~��GT��{I*ba���'�n�������U9Zꠖ;0�bJd�W}�r�)���P�y�����N��P�E�L
���Kq[����&�"IE4��_��� ^N�o�F���d<�ޥ�Ҍ?ಟB!h�K�CBf=�P�]�ڟO�{�i�w�Lk���5i����{�>{4h��7��t�]ӓ�w�Q�����L]�����i
�fzR!�ҟ�8��� 	|�=!�L_M5!Ά.N6M&!%
S;�0��o��MѨw�� �!2�&~SLŢ,��n|��rh��_��[��XW�|��.��$#��tX}~�v;GqХ�c\l�	�N��x���^���1\��2�.r��y1�O���Qv�s�q��&1��Ƒ��0>;��؞��������y��k�ݖ����.u�q��y]��� �����-��+�*��j����4���{���ZG]$�ߜ2����D��z��n��!3��3s�����������S�<L5�^!e��kbr��0��z���!k\�.8�[�����R���9����+8���ɢ���9u�!��W8bG��C�u6�('!�9W*S��u�񓺗>���F9�<+}���\+����V'c�g4���T�i�8?��Ny:Vsf{<�K�����(L�~60���&�4�!�k�w�>�ň���'wQ��	��J�Ґ�RE��4hq�383�1U�q~|��k烒Z2&&�I�O,1�G
�`̢,E-84�Lɉ^�ε�5E��p�\����閆_WOҵ�r�����1N��C�eP�H�W�'��Bg#��މ!O��˛sM��_W jvh�霩��ض��y�2�ޒ��P0)74����ͮS�d>��E��/���5'�jY�1�6oh�nN�¯�8S��i3�����x�
3�˓�\��=Ӂ]͆,��|�+=3y
�T0T���ޅ��Qb�����E����C�Q�l������s������4<A\i`��� &����v��c���'�'�1�3����?��{�MR�A�l��!���G��q��zHy�L�|�?58M>Kf5�)�8�j3��{�*���IE���<"b�s��ɱ�uvA��\)"��r7!O���ij��xE�㝵ek��R_{��i��?�g��B$�����YG�	xx��ԣ-M�DW��Ɠ�����%��������݉�Wؾ�Jp�g�Fu��vq��F%���x��T�%���J�䅟�r��˦�'h�=�sɐ���M�&�kgT������II�������T�
P�3 yM������o�:�'��j��'�I�x�-H� �[�E����PLFT���[�?�s��=��v��7��*8J��8k�Б
t����F�T�K@��ʌ���	]Y����/|�Ʒ���B`se�B[�&�^��K�A-�y<��m��J������<�6z��}�%�#˃3I-4EO��E�>fL\侾.�J�A¸����)�C_�w
�7n�Lˣ�U��1Y�=��Q�}c'��.�̞�'5w)���0:ֈ���.�2vۮho/��<&� y)�P��G9}{�8��\�QB��Bon�?yd�$U�����\�B���\^+f8��z�t������n�k�C�c�b1�+�6LhX	�\@�,d�a���[�,c�<[���y���ᣵ�{�rnQ���	�
,�zV2�h��5����V1
�9���p�/���s%~�6z;1�C�ʝ&ښ���?��{T�eb���2�O����r���bA���4�~�?�	��i��t�6�Ca��R��7}��R���X��e�ᚥ]̘Gq�i���(2�yw�PC��	�Ѷ�!�	��K�5�\n��֝ ֒�@�	��DM���{k�B�4H�D�{X)�}q�ĕ���l�腀��Z��fpY ���CJX�<�#.�:c7s�3��4ނ���+<X��p +�P��!
�3�dbڰʁ�����d����%p�+k������ ����E06q�9T��$�:F!��]7鳲��-�]+Y�H�@����a�	9�_2�S��:��/aez(�i��b;�DR��>uLI��E`F@{�ƪ���:��`���D�m���e��Z�͎��A��­��A�C�;lhԂ�<��샐��1Ѭ?��7�9�If'dG�A}[�o�����'*R���B�
F35���6og�Ui������c�2ܺ�̣R����FzFpX��p��-aŨ���Ԉ3
���@����7���6ju]Ъ5隙gc⹪M�t0�Gԡ��k���'CuW$��;
���sMR��[/��助j��^a���2��Lj��=E����am�M�!'o�]��8j�L�"ߥ�d��� -x�)1'J��q�KZB$q��> ��C�^a%¼ ������7�4<XU�)��A�\�W`؉�����S�8��< ��Q(�2��o�s+	�ѕ)�5���֝�,^"�C/gj?���|"����.��6�+!��`�Sw�Lu�jn+Q�y����q��-�%I����~f�����vk�6\�w�v���N���=<��8��cs ��j�#���K�Dφ�6�V�GD�H1*����R�p|�����:����ɪ��uM8���g�J�gx0�p�����ؼ���2���ժ��V;4#�OHcN/�T��W�ps���0nqЋ>į��5�0��%�7ֽ��C�M����9l�g���p0,g�����mZ~vz���ު���k8�Kb �d��i~K�`P�#�h|��J��LJ�f4�j�E	Q�B >�М��wBߜܖe4l�Tnt��8�ӾX��:�{ݱU+G%�M��*��h=�`-Ż�P��]d�R�����)f;@��nU�.�'���A�6�^8�S[]k�R��K��k��]�,-	�	h���SBUܓmA��>����I�g*	-(�5z���|���������<ĥg�vƵ �>Уo�2g�fO����g�}
�J���<9z�J'v@U��h��:>9H��qd�k э]ol�M1el�O���p�雴Njm9�4��Y�����(��x5�q.����|r"�1yD�,�M����W�;�������[��2 �7�_�GfF��x���_Z)$΅������t��9�ϊ��:#[Q�p�㸋'���!|� h�p���0�"�� 	�~�& �uR�@�3ZD!�p�gY���}�-��j�5��7u��`!8�j?�RϷ���V��X��Mr����H�Sj ��T��%hT��aW@��Ts���W(<�FƢ�0��FV�Ѣ�=�bА�+�&�H�%����=��u&L��rϏLoWl]V���H1~�I
K�,I�4kbZ�N�9�?����x�UG`t�b
�� Z�� ��H�����2��싼�$�-Ov��|Iݳ�����z`���1�mz&��1p"�,/n��4�A�1Qn|�?���N��R�;e���ũЭ qn�L����k�ȯ���T
���W#::KW;؛��21rBG����3����Q���N�ʅ6���J�鶤@�0���"o��l3����,��]F�Wu�j �PtU�b��Hr�d����ֈz��� =�+�z�>�{W�Y�@�S�f�B�r߬�=�@^g}c�8�G�B�) om�O)K�8`���Ug�nb���p)�G+���JV���9��<����
����~d�t� 3��HU�vfw�gs��Vt+��6K��$���~^�&��\���㊩��o�z��&���I�c(Ǡ+� �1�=S'+��`�4�Vd��~.#W�����D�R�����v��շ�������*�]6j\1/ɂ���V�E�a�3�W}�$�JbQ�
�e�yϾ3���R`_�-�yU�c�g���:T��-�8E��a�jf���8�:vc���{�ELO��9GR�//�����1��Q�����sp��.o�|�A�̒�畃!�a�!Uy�C$�}��أ�C�fC�6��|Na�	Sr�k�����Ό#�N���d<��@�kl1UՎ4����F��j�o%�=��4�=�q;O�mr���o�M��^��V�e�!�c�3�:�K3킫����@e��8^��s�T���f�uXc��H�[m���RW�}}��45j��>�EF�܃��a�]����]x���ߺ!C����K�.֛�AV�˴s廖ӃB���+�	���ᄏ犘3�6���-�}�h�Sv��.��7�_�<CZ= `��w|㟴�ޭ�h%l����v��� N"����ڮ
��R�K�������+�aa���k�y�1���FK~������#�4#�KW�к27#g�iQ3xhI�L.��ӟ)kX���>ٹ�x}��V��$�e��]А�Y��F���v���ٹ���p9��Ҡ�͟���<
�⒭���s�ثp/���S���Ճ�0\ �]�tǰ�Hf��'[��M�6<���=����֬4F�=�a1Cu�M���r�8(#/��!0���	-n��)��3����Q�h����� =�!�m��*W�%prD�T�<�;U7m�����������' ����D΀:gk�`8k��^�a!%B����F9��B�`:o�H�l���)�8k���KݜxH��sVY��b\4u�;���<�ٍY�zB�TמI�,v��-��3�A�j��n*3��fċU ��9�^5�#�����f�σ�.��V6�2�����l����v2��nɝ����'����g��j���{��c$�Z��r*�q'�XN�tp�0�:p��b(��<Zc ��˵n-�G�[_�No�9I�ܔs��)��E�>0�K��cݓ�T@G(�}N�0��khA�ҭ���i�4���%� >�
h�R"=��x�����Q?@)N�&�I6~i����B"�=Y��R�����&����j�JZR���wKb`۠�-M/S���ߤ�,���"$潕��$u����Ĝ�L�tޓz�M����������@��W����"�|��� gkCJP�ިF�T���m����~U��Ϧ)��m��)*�@���?���!ne�q�8�4��Z8x�7;^9wL�@,������޳߰iV%rp�rvT|i4'�)������R��2�Ù�O�xy4Q�ұ��@A�3��+(�u�(eC.&�q1�qS_@n�8/1��Q�G"?)��saa,Q��H��Wԗ�۾��)�������2��Ffp�����5�x�Vȍ.T	�ј�2����Y�N� �$�����*/�5p\q��$�W$�w�]����)d?q�)LP#�[p���z���٘��9�e\�d�1dj�uY=�r��qY1HA��-���+������B�u&���Y;��2�{�=��r#���D�"h�4�*B�)Å����N�h��=� >���	۱�v�l���z>u����-3A�|G%E�Vb�&�v#�c˗-��G�bCb������4���շ
8aD��	��j�����'�lt
���u���!�$��x�9)
�N�����?�����v�ƽ�a�+P�iVL�6�y8�Հ��c�>_t3ʯ��Do��hO,!n�6j�aW�J�>��6�o�~�H ������|�v�3io^��s���5���̳H��%�a5?wOAĆ�+>?�p����΅M��g�����4WE�xưzyLk6� 0�u�M���d��b����*��`���m�j՛k`��1�	[r1X���ٍ��H�o�dW�8t���N���.���W:��W#�T��۫;3j��i	� �I>}sT�Aֿ�?�[���P®6�P)r7����T2:�}Ճ>+	��
��iN}�J������t'�Œ/��VPAT���%�Sm^lI^���8� 	�ߍ܁e����T� r�y��.�]��M;�C2�F��Q(�K���o����g�*��5]R�r�[���p����Ա-l6��8�'w�)�I(-�*��������bC��>{-��f�Uon���D�����5S0��mǰ��0�㤗A�M�Ӟ-����κ-����pީ��Ȋ��P�e����3��1�6`y ��Մ�G(�*�kt���μ���>���V-�N�I!��OQ(>~�N� �M��J�`�Za�	u��|�U�ק��20���!��G%c�H%2k�2ĵ��q�DG�ApV���筐@��e��&���K���M�KJ5�|f}�Z&<u����بwsO�9@u�������g�lt	�Gv��_9(��B��fٮ�t�gN���E��U�2��%��Kf���u��
l�sz�P��p��)3e�ѽ��[�`�}$3���C�6�?jХdD'�f��.	]I��G�|�ׄ9{��9���^�@/��ɕ���/kib0���㤵)�'o���I�v��q�ƅ2@A�y�?��R���9����h߃��wME�*�}�� 7�����h*^�\�!A)������f�OO���В������<����Q2��?~����~
V���B����a��.��L�	^�"m��c��d�#t�ؼXTގG��	��~6@��s��i�ç�>D�f9P��hxLW����M2fM�>� `j�ٗ�մ� ��|y��x1�Plޙ�U��Ŵ�m�=�hy�:�"�j����d t
�XU���fZ�R-p8SxuV(���X�F��h�_�~�l�2~Į�s@s��lB�)��n|�W�`���"��y�a��0:��t����d%��fR�Ndn��U5��m��� H+T�1"���_��n���x\#���cjg|a��v���$�z#xu�d:�v�#;5�)<�<)�Y�҂`�p,JT��eD�8��u��Ynb�7�k�ʛ���4#̾˯�Q�<�����h����)4چp����.�Ez���ף|�D�@�������9=��7$=�'��Qf�"9�Q�f7����˵w�_�2�{혪���/Zo:s�0��D�F����Gl/�4�%�!2�4�P���Q�G�k\ Gwi+����ZZ ͈�2���d��
���s��+�SJ��覫�7��uu֛��'��T!��g�=S_r:Z[��>��X0���+����[���g��*�O	��H���A��9�GfQK��SQD _u��u:9I��Ӥk� �k��My�z�p֥籣�O��(�R���Gw���妍 �8�:����٦��|��Q���#n�P�� �c�yƿ"��&C*
����H���l�9���G[@^CE�%H�+�P��<N1�-�1"�`/(�܆M=e��vۖ�+���{�{�Ʃ��P�8@��l��y���;E?/�ڷz��]
����.m���(��I)X��-HC��-�G!"����)�d�O"���F�_S��c���Ɓ�z���)������ۢ������c�[*VNR�f_�16���������0O�|��+��|��J*�uKa�s7C�(�M�T9�tADGB��w(�Qj�}�* 5W��36�٨(�_Z]��֭��\��'y�ҩ)A �a�qVl���o
2o�f"u�f^r���֜��.f:����3Y'�	-~Gb2�#S�c��颬�j��As(�&�|���Pxb��W|-�0e�9�<��I}��jM�Wp,j��e�d)<�A)bZw_cP~�����T��.5(� ���J�_\嚵
T��)҈�hu�IaoAB��V��؏���V��=ͳۀ
�����%�'��%����=�H�:�����:��U_�J~�_��<%��	݌��0ǡ�F��ݷ�H������HF�q�2p#C���T��K�])O{nzwi5%�匕�߈4%�*���ea��9���+ܳ�f�Z����]�����VQo"��[ѽ�Հ\�Z� �%�\���m�.�B�����jj8��?x��,����E�F&��ĕ�Kk���j�L�~�X��g  j���;��b��t�b��c�����H�d=V(��
�{�8���u!�D�>����}v���qsM������ӳ�d�4Ǌ��Z#k@��-6���Z1BкI"Ƥ3�a���ˣ�^>��^������t&���}��񝯀�y� ,�:���ޞ2��v�G�o�h��/�y�����%�=�������D+쩁�?KciWF��w6�w�2ý��a�N&��H�Z�}�
��7��t^��n����f�Y+��b¡����1D��U�N����%�Ȍ�X�l"�ƱQd�v4�b;;��H��CQ���?xU��TW� ��bP�^�ҩ��+�p���Ƞ�x�lЙ��>�,�E&�A�4�7��-�zo�H4#�A>z��7o 9�m~�sJ��8A��.�����qnw|��҅��T�I`�y��`-���_��=Pe]�2��k1�Ujv�*N���4]�i�����e��np
h�B6��1d�{m�ۃ5���k
�o𨝃\�y�ힲ�M�M��k!�Jb�Vk��<���l�øb9�W��y< i��OK�Z���jQv1yxP�k��P��q @�2��l�R�V�'d�������/b�A	qS�����0d��x�N�O��4�&�$�0�NoW�:�V�����SȮ�q�_��m�4*V��0��2���ji��G�]
���T��ވج�L�_�ZKt*9&TR4I��#�o�����}�Z�e�I��*T2,�D�>څ��o��#$�o��?@��U��zW�ٷ����Qy�ox1�0���<��&/j��g��'ĝ���^Ɲ�y��J���{X/��Wa⇲ȭ���[݉@c�G�}�������u<�N�����e�x-�n���R�1��cU@z��wu' i��Y^s��Y�T����>���D��ny�/+n/S�5gʚi�������l�#+u��������t��x�vF g�DG�|��Qz]v���vV3�%W�ɒU�s�L#��h|�b�ye=;9�i��d��2$�ς����3	\�F���XiM��RK7g�y?)�mw�n �$g.�ќD �R��!.�^!A ��)�C׽���Kds����@\Β��dI/}�ƵO-���D\rCSl���iĈ���T'���N�}a48�4/T.u���f"�:�7q0[�,�z�d=�A˙����H�A�'z)�Lq��$ ��A��(�Hؐ�Cz�ѽfZ���a2a���F�j��?\�55n��3���@=�,n24*��3�{��_�8��Y�pP�{\�x]�ٌ?�2b���6hw7l �a�$����d�s+X�FQK	�RU�-��x��Q�s����B����k�j?���r��
P4�}�FeR�*�D!��#�2U� �5��jL��몢�=O��{"���,>Zf�i�@�Kct!;T�<y{��),~P���ҝ�+��kQ|����(������k(g�4��=�@��_���(�-��H�j� ��ٷ%Y�`�(,KĀ�U���J�冺��0���%2�����3�lE��|h�y�A�> �ב��t�J�5�Ev���fDr��)9��\pO�링���4?<�(��#uswz�K%�[�!�tPZM$x�r�ڭӬ�}�w��5�ȏ���ԃ���jE�#����k���ӻ���'���!v�K3�i������rJ��lDn�=c�9`H���|�%�7�n1W��� >��
6 0y
�����y�$i����]n�����v�Q�i�z�{�I4�-fz1�(�uN�Y���΅%
���땰����[E�hEp	l�q���wP=���vvO��Xt�Ot*�klZx����~� �^�\ h3��[3�]r=vq�a�Пs�A�K�:��-pt#�T�:����2�����'N�.N�vQ�ǹ�A%������'L�=�����8Q^��d�QG����a/�@	��ǐ)	H�xN�+�DR�&�@�3�'a����(�0@M�6� C��\\�W�[�v2�� 3�t������Ɋ�w3|��ݽ�Ieg�u���+mz�EH8������������U��h�~�=9w���U$��ƒ����J��z\Ǯ��U����ѡTd&Ȼ:�zFˡ%,o�P�>U��Z���c�K�C�#��!L���&ǀ��3K��ۘ�|�kY�u�j����9B.���FaV2��?�@�>E�,���v�E=4�B�8�́��u1`U�E�جa%��)v=9���̒�����)�!4��L�yj��»gb��,�����������ᑙ��Vn���������"�p����c�0�Y�+w�\�RK�q�,���Is}W�Vqؿ����"l���弨{c{I��Ɛ��	�?�D�aY��������
��O㏁cR��"hT��$H�_����N�Z���1���������y� ��U!V�J�
�8ޱ]�Z���Tc��h��%%g��b �5��ˮ��Μt/V�i��1-���R �^JzY5/Iz�[-�}(������ s$�nn�@_�����:N��7��S��\��ѧG\:6G�l�S�':!X
ds%�H]��:�ʛ��>ų��S�����dSU�ͷ+�9L�����w�$���<���(�(���6+��Nx���6�-7��E^��}L��/b�i��5���[�	��Kc$��3y@E+�OOd��b�Ӑ�6��i��z�ԵA��L�-̅��V��:�f	�y�8~�e�O�`��X�=�F�Oh�1ySxO�|��|М4����
������۱��Ƅ
~��V���/�q�ة�g3�ci���/�Z�n�3+4�R����Th�&}|�c*p���K:3����e�2U�fXֈ[Q��ʉ��땧l�$m�v�[0���)�����o�(��Q�S�sc=�F��[�q(�~���x{Z�4�8���X�����,`9����Ji�˦�/w�l�''R-����*�#���[���b~I(Q�v"�}
��AڏmN�����ύ#��Y�R<��%�%��o���^���RN�CON�Ca�;����;����f�GTZ�N�4 ��p5`{�`��b+��[ �kW(�3�'mX�0���ncS�bԮ)�(t��I6������R.;��( ��il��hʥ����u�U�?�Q
@,���*����O��(��g��v�c�ކ�J䬧b_T�*�Y
�aWWG8�p?���Z"��ʱ��L����hI��1z0a��y����u7�s%N=�Ef����QD?�u�*�z���)��\<���{P?f3���daIPbYJ,��Q����qэ	�"^o�SU=V7K�;�]"�4����o�a�%4�f���0A�MQ�GR�XUtc"7ż�o�{������3��Vs+�<ky���a��&ůd�2o�~*������.@�"�J�L�#D)�J6-�Y�p�Q:��Q�:����IU��H��f� `�|R_Tͫ<������Z������
5���������R��K��/&��{yr��x��A�����p �T6�G$/a�S�k:�h+5ط3W���x��o�#��FV�b����(�]E�U���#�[��Ң�h�7�O��CC����2�wg�h������7y
����%	�͂�HDQ,}��2�(�\�Db�M48;��:�p�or=��@)�?~	�c�&�)[��ՙ�4ӗ��«�����_V:+�*��F]4��<���s���E�bT�7�8�!<�P�l
�Dn5������^u,{���38�S�'_';h����*�Ux�tM���DT��l�ۀ Ʈ6ib�&��ZDU���QA1=Icg���y%&�o*�FF�{R.��\m+����pfr�I&��l�MK�hؽw��e֑���K������g7���K�KJi�R���o�$����|k&m9OOD���ө�bϻ��J�4��%>K�v����8b�{�e��=�13GL�$�T��?>*2�	��T�S��[������ A?Kz��-�ǲ:-�4R����s�	��|����Jw���p1ܷ3�[T���d8���#`'����2�Yl�j�a�{��Ы�Ma��:�?�E�n���!�x�{���3ъ�Ũv�k� 器�>h[ڻSOd�)`�F~{��r����&�¾QK�U~���Ln��q"� q=�F�L������������U��,8�!��o\3�c?1߫���q�4�`t|?���r��TJ}���N�s-��6�(�� �e:g��'�J]U�⎭3"����'�3��O��_�<�zK�0,��U;�I��u-��è:g8��zp'{&
_����1i�%^;�DZʍko��Y&��?{�ڮ'�����:HR䂌
�d��?��G'���6�L���7L}�l��<3��h�`�y�Ҟ��	��͜��i�]KB�t�|�d���E���k�����c-���E]�~gO�A�e�FXT�S��_K�ۑ5�*f�rଠaX:�e� h�E��2Y(&��k{.磞3��&��S�����V'�N�j���9�z�Wq��jW�=	�(��ET�?��ʟx�	�����^�|d8t�o �RR���"V)!����9�M��Z0 S�����T	J�����c�uC#��d�8_�lY⸡Ӟ�k3�J��cA��02��3{E���	uu����Y��v�H����1��%�P�����(�}ڐ�I��$���X
�����(V/�`i�#��D#��o�G�Û<螺��])�̤�^�5���:3�XnL{ο�}ۅ/>!��u�����Gda�@�	wϷ��~0�E\�0�(lԔ�0��A}�)K��<�S�
�Cm�+� Iֆ��	���J��FG�8#v��/@8NCٿS-�.���d�ȈZ�4ѱ5ؾ���������"t��4]7�&f[�����p��埰A���ޣ�S;�O��D�}n��yAK`�b�(�f9���k���>C��kg���Iv�c����*�r��$hrj_�z�tf�_��� g�a���-�X��@��
)��ťk����G6�����Y��6���R>���� ��>p�Q�t��5^5�`��d�|�����CN���?�x �w�\�o3E��z�6R���g"�7����ݭ��\��9���Zg���pz�`�)
u���#�.ī�լ(̵�1>E/���`%��G�\�;@�N��A�@����vl����J`x���C^v��%_x��(�%ʪ���,F��P���0ah��cx�mی7(�ƃ�w #G2E�lG^fwY$�u�j3uK� jXJDB�˪Z�gA�-wŦ�p�fWin��B>Ŋ�������-1�q/����^bʆ��V�}y���}����e�J)�-نK��w���J������H74��w�������)x�P�"/l�~=�R��w!��3������[�uTl�/ I�R��S�쇄f%���"0@M�D��w@\w�Ջ���س3h$�^f�@��, ��ͭ3�݊d8Ռ��X�J[Y�ˉ�fa�iT���g���*�y���)������s!�AD<�����#\B�������1��[LN�cK��T��܇?��Q3Π�e/%U����o6b��ߝe�
���}�1��A�=��`%��ZBY+�.|������@�S���O � 4���3���<G��zN;U�'Q�eqڠ���H^�,,8���5�#�g�Y�Q��懷k�D����Y{��؈����ڬ�����ϧT8�T�e3$F&sÊ�*6u�IK�`1X��&�r�t�U6��*@V��U�E7s�>S)�MEꬃKj:��"��<��1��c�_qxQ��p�@g����n��;VD텰y���($�L��*gO��/�,�S�;תA�����~��g��8���/�xU��"����V�����-�{���36RԘo�iv�����j{hc]��c p����Ц�>����h$ %q�ofAai���sUN$Rl�	�!�6��|����F*f����8��1w�������G�,�jh>���=/iE��Z��\R|���gxwǡ	�A
���<3��,�G�й��ˑA�?-�+=�%�2oJ a�������L!������W":-]�����x�f����ew#�y��o��_��A�ssw�F�CL�Ȗv�p��k��F��lm���
����fK ��]���4��WVKmo߿�ջX�^������}�Ѩ������0��e��O�WQ�R��v��:ky��J�)<&�4���DȔ��Y�c���8�n�Ӭ:~n)H�©�i+�6 m��9:�(E�\rG�����c�΁8���� ��_Q0p@N�+��F��\dL˽O���Q|� �O�I�l�0|�m��)��͵o������U��g5r����X��&������:�����\��Z'�l�`1Ƹ�o���a�{g��G��%�K��RB��ۄ�٬;j0�8Ta�Ӓ�`R+Q/��1�k�x����N5C����
��\��2��a�^� �uNp^��˞_���V��l�� $Rd���Ъjq��9W���a�����[ي^0�X�#:��۹1�T�G����dH�9��E6�yW���ۥ}s\�Y/ƹݫ\,��oḿ���)��=�G��qjw�V�.Gį�Hv��KI�����}��T�%Rl��C����E�H�W�����9O���f@%d���Ee�M�g�&�4��t_��ϯ:���r�����f8�X/����0/�؆g�Ee�e����{9ǈ˟������7u����	|l�>uIt!g;�U�z�p�Ă�!�(�R��;2�:�ie@~�Q�Y�'�*�����]Җ�7�M��`z�7�]�|�5$�A����E��en�3uA�'3���c;A��ƙ�ɛ:�z�u*��ڭ���)M�/��o޳�YLiΈ����9�B�:���/�����Mp�^��$��O��)�4� ��e��e�_f�O}`XF�Ӕ�ɹ��j۞�{����;��e�y_��僑�l��p��j ��l�� �ȏ��
0C��ѱ����UwF۝N��_!`�K6U��:���~ۿH��T����W�xv�,�dl5���L�� )N&4��:�]���#�pߊ�;����4�+�:<�k�u�B�2�k0�Aq�L�\S��|�y����,���7Nyғ��<��M�([W���ޤ��c�8{�J����m$�2�y��+���Mo�R'���?�� @ٝ���L�B�	�e9
�t�ajU�(Jĕ��"���8r/�r�i^3Ax������+�}dO��f���V�y�:�mqaE�)3��;U�:�H)����HK
Q�V�>���� :l=�\�b�!��J�AF���� ���f]9��-����M�r3�H9FAթ����q�_GPx�3V�u�ۖl#37�:=�P=���]����B��Q]:��Q/�ׁ��{�=Hk\p�>/R	�/��Ȣ�<v�����n�"N��%!�)��eʿQ.v�m�u��/��,�M�j��r�"P~�:e�޸|�)�}'���E�q\�?@��8����FX�7.t�������+Zp�ȍ�N_�h��G�d�i5�#]���b�Q�~���T���v�"$C���W�mY�_,�ka]f��X���#\�G����,���I��rj��9E�����-���u+b?�b˒E�$�Um`��Ti�ND7�qlݺ���ÅOO�J��\/-f0:�]�hg<ޙa-��4��.)��E$z%m ;]�������E�s,u��7�+�j�+����d˂Ȅ�� <{mz���_%#��ЦCA���E(d��	2)�=�� �1#�Q�#=�6Em�U����ǿ���G�/or!�ϹV�L�8D+�8�D��s���>D"����'��})�ќ��:�H�3eAү��~��]��z4HO}P_��U�@W������@�.����w�]�σ���{��򵦄��ٳ�K��L�#��[���4�eH���Ծ�:p��[�4\s����d{�;���Q�Ao|��`N���h�O���/��Es��$ҭ�Rn�OI���c��R��(�e� {~����+�d�y�<���i@�^jɀ�T�~�G�\� �C��=����b^��^��c�iZ��'<@�R�������yT�FYFw�$d���� �?�q��SF�Iר���	K������H�^�e	�ڋ:V:�`*�_���؃tQ:�^H�G%s@�Z�ǹ����MD�;��ȝb��MMv�2�ݭ�s�H�i޼'������"H���yy�T�>-���B
��#�;���V5��#Gp�Q�ë��˯x��@���ڍ���v�]���e Ѻ��b�����+q�G�i��k�}���ƻ]-�T |}�	d�=�r$�&���U�U4�)����xl��!��ො\+JΑMNn�E�P�l��`R -��GP�,8�h�&�
��,�� %�Vy"*�h���� o�+Ŧ�h%��Y�m�$rCNKh5x����&���g����?�T�D�hP���6ў�@�.���h�F��j:���P�^c�?W`U���nش�x(�L'�C?u\��595��N��3����	�;��l�<��j�Sit\���\LS���B�c��J�H��R�i�����r�FMg�нf |�b�6jm8��͓�YB ��O�>*$2��%���,�7t?���RJ�9�K�Oo5� ���P�Sx/a����:Gm�% ��S��y��#j�в��ܞ�u��c)�aU2%ћ��8�k��1��Y�I={̆Le�H��eW��<Q0�ΰ�/n�:>�D:}�bϽ��`����E����(< ����%\šH�oٕ3єBQ�؏��ů��]}pwE��`�v���-�tN�Q������,Wn�9�e������t��:h��\��x�ʼG�[@�~a<�5��Q'�wn�"I�U�O���6�V�T�r����Ũ,��n.���6[������6+e�|�Cs� 4��!Zv.�Q�]�a%_,{v?�������І�3̅ǡ#���\Ϊ�*a�Vl�)KވJ�J+�G
���V]AE��Y��'��)�w���I�#Ro/�Z��LhL��EW`S��R=<E= ��4�P� ��n`��;%���@�rQ;�����yt����bb�W���Q� �hk`�c4}��3�bQn��2oۯ��z����(f��M��`��g�{|XO��5�"y��,o��>�/ �~Β����LK*q�Ւ>{��3���o[M���!���ޙI�����S�w��0����]1���Aɰ�e̫���l�r�os��.Ĵ]��Z& �z,������T^T�^�z��z�TTZ��Ѝ�=�"$-F�`p�iւgxT��&m~�%�a��탑�Cg��>W	(фSM��V�����AQ��r_-���?�E3#K�
ãP���ㄥo��,�^�Nki�9��1e�a�g'Ϭ���ys)�\ƑK�b��H6�.���R��w����+�m_�L3�1ٳY�/��Vn��O���W|��0S�e�.��~>��p��Z�+kk[�k{�PZ1������w1���-�U;=��-�bt�,��;4f!jz��3 �Y��ݬyl	���Fq�����P|&�����/���8�I��.�SRA{��<���&I�Y�q�=�cꟷz����V.�-�I����F�M���i8����fĉ��Rt��f{<� _Q�6o�n+d��,�8��j��A�~�	�z=�+������6{9�6���;����	�tY#H^]j�#mc�섪3�5��0į4M���g3���(~;�0Kv��v�9��Bu�Ok��@v���:��=n�`�U73�|�Ђ����_#=�Y4��ÉC�(`>QjH�B"\���Hv����ʜ� 
�҇Cw�B�8�.����� *RH�j�����H5����g(��~�����X~�=�r��4��sٱ�w��j��VI�8���UZ�J�FJ�G�lr`�#�Ȯ����|�a����Y;b"�z`6��v�\�®��ѫ�ȅm
�T���}����&A?-���GU�fq`-�4[P\�XT���{o��tb��J��D��rT�yQ[�k�~�$�z���i��܈� �w��@�b+�QZ����ֶFx=��Bq���J*�n
�ik��z��(skw��&�Ϧ쵻oҥ�G.�	j���������+b��=��/��<�s�^Ǚ����lP4�I4��<9�,����Cՠ(pdJr�EK�2z�#O�`�����z�>���zL\`|'��W�<��۹�ktX���[���-�mb�&a�>���L)stٔ$�z�q�����ISɸ�����N���tX����=����~��!�
Xͼ�C݋ky�r��<��dL�k�+�����Ce5�&1u�g5\X�5����{�_p�"�91�o�н����<Au�͒*Z�^NX�/e���yҒ�©MJ/�K�e�)��Q�
	���j#E�I½���yOl[��{{��������%�����M�{�w�=��3�^�v����*���vr��=�d��s�x&�"v.WG9HfJp���Ź�H*�G��d����wg�Ja�����K�S�_Z���>[,T7��"{j�c���>�($r���NO�ư��	��a9�(^4����}C�xv���>ɰ=�GKt͕h��� �W+������g���!Z�6_�` 7���{ �h�Y���:��%|%���,���]x�_y¬��@�1�OR��S��[�ŏ�;�cj�9>�uTZ0������[�ؽ��vB�Ө�5Օ/Q女�\��R�[s�/ۜ��V���e�3{�N+Q�\�a�٦�H*�H0�֫���z�V9~��Jղ�9v�m�H�fT
-k2P��ULz�[��Uy��ZY�����P�G��"o�%=�(��c����1�VB��A[Vi������Ss�-�E�O�`�2]S[F���r'r����A1�!�4���II�T������5I�zZ��*�Tz��o ���.�u�e0�d����uc���ؠ����?pX�X�ㆱ����멄�0q��#���.k�H�
[ܩ@Y޷%���l�Ц�A���Q��J���A�" �\H2Eͳ	q�r�]��{R����N����Tޒ�,�6�
v�������V(�I
�뭲Xv3��	�i�V���r��q���m��}����XD[w��b��)��[[I7�^kB=�x==nwB��Pm�ؾ�scw�Y�m3�*��l�*�F�m�0���QG�J�P�
�V-�P��4�}y]j=F�/��XA<SZ�ȳ�>Xq!�/DiYq�r�)g�,E��t���@��_#w�)Z T �~I���F�Ք,�g�RO\�=IO)�=K>m��@8���� s�+�-��UE��l��4f���}r�W�v�̡�2�xҔ�%���8z2g�B)P���bx7�[D{�T���/�����7�+��>�u��i��U��Rք�ni|o�;E0��2��u�����pD/��@�h�HƗׄ�u��5	�QoB�K���E:�p�B�C�rV�UB��bn���؛J��	��������D��#|ȋ~#U_�4 #�s͝y��U�R�=�i��z����Q7,����b?
� �����/
��[B
)�˥nx#0e�Ņ@w�����G�iҥNal��E��]՛v�x������^+^2�Rʮ��+���z���ljobm]_�G�֖�ɧǬg�CY��7=6�ծ��J�t�^��ߜl�@L	��(BZ_�;�v�g��X������ѵ�K�}��$����H�ra�M%}��#U{uR�=��u�>�&I���h�����ӷ���?`��k���yT;�Ӄ�Y�`��v���2mC�qį�_���?1�$VO?�N�!�����!�� a/ٌ��j��(b���m����'k���/9�������g)�1�~4�)X�
�<z;�'i^��L��P7ƾ��Hw>T�ַ�O�L������7��V_s���Z6��Ԓ��k#�l�-46X����|J/`7@�Q*�w%�����*�zZi�[�>���j!�EE�?����,ɑ�˸�T�T�����˒�a��Q榲�?kB%0�u��]&��QS ��A��O@��@G�l���+ۜ�+�-iB!�/Y�%�,�}|���5ɘb���A��� RS�*@�@㈛(��c{�1ԣmʱ+�~δ�J;}(�^B���C��n$B�����q��Ҫ�_ =�X,�sx�1oZ9�C��J�ʢ�����t{����:�����fdt	�V��M��)^��T<D0m�+�f0'؞2Ǝ�J�xj�o��㍵��/>tݑn61�,����|NW�q��+��T��/�����mb�]�u�h��m��&:׎��S�,`Q\K�m�:͜{�8Y�6yҨ�� �����6X���:��3e��s�A�K�f���~��u-p"�CVB�{�wr�#�{j�v�����e�(���lS��rtoVK|s٧��J���t�U��'i�&F5X�F�x��e��Pb�x��}qAp�=�Aa�?A^0���3f���~0q(y�0SŦɳF�L[����a��ՁhB��zз�au>^���B$J�NR8�ZU�)�}��I��Ջn��M�;TJH�:�[cw�a�c��ogDҁ���.�^�k(�&�\�.��S6tw��E�c���@�����ڝ1$����b��~i��P����\W�F>�sLZ�~�����!*6�Q,�E>�iȗ��H����n0�%�]��ݫP����,��$�Jb��iO�isp��f?o�����P%z;WK��a� �f&��cOnA�s*O	�S��'Z}Z�ȫ��\~�.��oW:מ�xP����<�l� �e�,=�n)���2-zϹ6��.��&׽H�=�Ef�^ιzw8c�J}e�ל��x!����
���z'�#�]�+�6Z-�5�b�K���e#�D(=*�h@�\�mј��]�Y�=���R!%�Oύ�s\Ӭ�݇�uwVN����]I�s��5<ޛ�,�hW2��0�e��*ڤM`����5��/d��E��Q���F�ot� k�;�vu�'��ƞжx�Jv�R�Z+��_ܽ�OMI�R}1"�ui�W�7ʒu����pm�٥!�W�-���M�p�wx��Yd�>��I��ea�K9��!�}���f_X|o��L��J��Gt�XsC`���yU��XzH�~�\�ӆ�h�J�i�\Ks��}`�G>�7�-�<���N��e��
�nG��]�%x!�:M!no��Z���%�d�?���j��pc# qG�ҹ��<�l��A��B+�YU/��/���R��4�.��kњ3k��(�^J�6���L�,%joX�n�KF���e�g��V�2U�n�p�����L��q@&p9j���U�2dK"�Xt;zQZ��!����zj�U2�Z��t\\����ߵ�:.`(uZ����籊;K�Ow�������7�,���]?o̒N��ܴ[��ls�hɎ����9z2d�K����o >A������:-�!��нؖ_��O"ɼ@�%?&��6����	>Du��6��dS�1r�i�d&#��Z~�\b"��챷,Nz��1�KOyZ<a1�؈��m�wK���o�ss��-� �;��?�.�.���MJw��"���9����I��$���@Mֳ�y��5O��^&��F�����:M�z�ԯiEc�vG���"<����20�m�Yz�5����5qBu��!����K	�Sxa�p�c��Ce�#B
@��E���i?rk�F,p������0ߺ) mi��	`��[vӭ��v5�-+�xM+ܽ�J�|+�*y{!�ӥhq!s��o-���.S��yc`�*����s�7���I�|���A����%�չ��!&&������K�*��>IS&B�8��5`�J1j��@O<��~w����O{yXЂ����U�PUr�:���wy-��Ǝ�3�"b* sݦ�a�r���_�(3�<�|��	��k�U~m���֝��u�\���ۻ��1�+��/j�������[�%�Ujm��O�
\f�T�
��9�tN��b�\fqd�2���qt��ld[}�v�hLHţ��9E.�=��
�8��_��*h��*���7����^ �!�C�^,�������O��r�mC��#�L&���b�c�Ճ]8EOH s�-K3/1�$����滰�*F}l��z����<�z�3>e�+&t�i6_���h��4y�Ů͒����ؘ�)U�$,*�A4��rs�DMΑi�a(�q��JO���s!ೖ�Q(�;Mq��`��$�_H8�^a��׭E��%�#~��'�%��ΕR����@^����r���.1��w �y8F�I
�mb�Pк��f?#�؟�lTnN�ڹ�-K��6�ND�8I�-��3v��.8t���g�p�7����൳�,TG%5[��R��J�N�oT�7[TTy�1�?����%I��y���& 3m���%d0T�i�=�#���zO'Ĩ��uU|F����rYu�ޞ+�:a(���x�3�S�43�S$�/5+6��P�K��� ����cO���"P@�^X
)�6�_���Y�Tc�&
���r	Ú�G҅��1�}�bI튆�kn��M��P�~	�c�/��la}��ʛ�tű����hi_����>�ȗCjc�ޮy���,Kf���������K�v�~�=Ȯ���m�E��]iO��
�Μ�?��]��|Z��z��9$}�2�(᧿�.ڷxH��s�L�V����	��Aw�@׏�'3�"�^�����^��3�~kה�j@��Q �v@+�L�^�V��T%�,j����4��9.��,,q�\Vmb0xU���V5�L
-�;&Z;�Q֡�8
��D=䅉D���f��ۮ^�Y[#�3A��&ª��[-����M�	D9a	����5`�0v$�04Z����0lF��KX�oN��輪OL��i�pQ�v-#��3 ef�]����Ld�#h꺬{B��R���U_/@�B���4��Ի;[��$�פ_{���ٯ͐آ}�2���K����t��h�Ĭw��]c����8S��U�E����-k�n�{Bc#�1�o7@�ͅ1F\��Y�����9��:�5΍�«���:逜��w�em�_�h%����� 踣�_C���0zϚ4��v11b��σfOV��V7�P�Y��IJ�_�� U�w�wwx��!����\S�?�Xu;�0}R+F�w?�͙�kK�79��H��Qp?:ò|{�u��i����+͚B�M���p�m��
By�߽k��[m���F�j�o�\�8��89���SCk�� �֖Lvv�|;���ȕP�OG4H��7ߪD��H�Df�+]�.��v�6M��ɘ̧$�/���ɴ�l�4�2��1��[����"�X�,oa|J"��rG�pk�<]�����˭��d�Μ��j2>*��n�G��4���,G��sWz�ƉY'�}l�En�Kl��QelD���>J0g|�\20zR�q���b����oI�Xw�Ǯ�v�qvhYg����N*pHI!C`F#�sMh�b�D����5&WF����,�jsy�G뼘Q\�=�,����=��Y�S0��Y1%��հ���)v�m�f)2�:F��,���,�@�Ky��e>�d�Wu���@P��E8����HF�&�����B�.S�S���ϋ'$e���ú5R r)J���9�KY~3�	�a��A����˅��H�r%Zu���PIFD�~��L
O룬vS�Ww���m�gsiV�P92#�ӓ{ắL��`b��˓���<t���]������$��M�,��l��J��p�8' u�ޟ�I-g	B^�&���&̖i.8E4h�a�MPK��X>{} y�˲���nVB-�K�TD
�צf�~���g�����@�Y9�̅���c>���jj�n��<f���a�`�S���*�:�,U��٠� dY	��Y%[�y\��❐ �GraȀ���J�����_йJ�ʄ���f�h�ޜ�L�5�H����;�����=�� ��T�����^ӟ�M��[l��T �i+a3�gt�f��n������x$�Q�C5x�!����U-u@�6�t~Ck�t���϶?u�s��բL}u�ó ~6� �������_�Gpu����oH�e-�'����kfؕ���^��ǯ �O�E3���O{�#I����Bv�5�wy����(=�\�[���)�N�hp��3{������f:��Ҭ{���%5�t�a��E�st���9i���Ch�0�z��NU���;V�n��*�(0�7#d�� �V��U�cR0�c�i��])(j�.���Ha��z�6���K�����+�'Iڗu�~��e��wɨ������m���j?��\x���D��V������ꛉv#�=���z�P�Q�������F����wmY����2'�g��g���ݖ	� UùY�c��۵���^P���]�ֺ?`R 6�L/@̞��x�®˧�^f�YwkU��F���Q���ͫ�+^V��e[K�wݥ�+q���DjA�k�˷�=���[�M�~@2��/Bt#Ӗt�PڛS���^�nȤm'����o̙��_�-*��T��<9�:"L�r�l�|=�U:d�p�XX/�r���c�wR��\���os�rؼN�=ϵn�����vG	��(�[�d�~�ᘣ�|�S�h�g�f(�Φ5G��ed�~U�^�~��Ψ�&���$bØ��؟��!<�
c�Z��U*�FA�3Z�z%�>��)#�0,�*���%�E\Bb�Z��wh�R�oD媊���h����ࢼ�'g��v��d+H�(+�&䑍��SP0%`V�g?�����Jp�畋0�m�L��E��_���:�ET�s�h*�2��a.D�⊘; %Xj�wo���z֫��ǒ�|_j���wZZC�?Kx������(�y9�4~ݏ%_WA6�p�!W�G���C���U����3?���a>ͦ<Ϋ���{鿹��T}��s[؟���y ����J�y��2VGX
�F�8�ˆ��'$Dbm�pY�	����My*컔E³��?^��%j	��	s|7U7�C.�T���u�P�%X��*�;��^�xﻀ�h'(p'eҜN����k�u���V鬥XѬ�7�p'�3=�,L��Zɦ.=������HӯʐDE��L��>��ih�>o2��N��A��������
��ۻ�H����������C���}�S�$"��@���P�"sx�o�Yp�y@����Ų����;6����`c��i�:�B+�N>�Z�
��d���A?��h�\B'+�+��y����N�o�y����7g5y�d��]լ�)��7�cX+��G�fw�@!>eHDE�>���
���e.6�g�V�
[����j��o7��=f��r�*!��l��'Ǒ����\B�n2Ozv?mq�Rv�{����0EDn��"�[##X�?���1�/Y#P��L�4c�rS�B������� �ǿH��2�F�M/�t[�6�W�HDz����{$�v�iq�`{�]�q	!+��C�x�R� ^���_�C
Uk���(�����D� '��C�������Ω�~Uh����:���։61;��Og/BVA����:L��̟�����S�#�R��쁅�;���24�7�n��g�r?�g�s;kKu>�����c�f�Ե�}�gڙ�`Mcu����Z��~�L8��#��P�әٺ������a�n��a݈B��Ive���v���]W~ݟ�m����|�Up� 	�mJ��� ���T��6o��	�����͇��[؀��P�
���W dS�����"����1����g��E S��G��c��m���Cj�G�w��v������D�z��$����OG=a	���ߜ�5���T�|`������u��0�m@�_ţu����jg ��  �Pw�~��9#S &��<`xFc��Z�)�n�_���#�F
g�/TvB�ǰ����S��/��KQ'�:t��4���L�Dp��_�[��(,4����&�'ՑV޶&ۏ��+�H�=���+Cޛ���tC���<��"���q�i��ǥ ����D4���>�y/�3")�Huiw�0��[��\^�Y.ӐC\����B��{�������r�+����|�K�D����W��O�&j�G{d�,'Ry�]���J~l*����IUW�#!�vFJq$�S"����ڳ�������۽�� �|8Wʍ��9h��m�p^*�µŌeҜ�9R�f�}Th̅B	\s>b(�
$��^��	����P��4:?��C�?D#������cK��S��xWͼN+.]��>�f�w����o/�Ms!�F=�b�b��=��F��8��Y>�<1�b�JE ���DO���dz�.���UB(z�6��*�$���Ͱ�ˁ=9���SS<讛Ⱥ[v�FiwLgc@��B�u�<��� �P�i��鏦�7"!0���$p����	�mL�
����Kd�X�M9��a&>��Oq���kxx�f��_`�/c_�0DH��ņ�x�V�C�G.n�/+�Kns���^#�A������lz����y���_�<�ݞCN]|��X_�&��h����m"�yI�Т�s����o\�)^n�ag-�Z�������#�M0��e�}�@���v׊Ч7a��:B�ab@ѐH.�1�?3յ�����Q���^H�n�߸�s0{�Fih�uB��R��ߌ<�
.TjR$]e/<�A���珜����4�5�H�!&��+π�R=�lޕ,�F �b�E*)���"F�TϹj���V��k4����	��X��f -��JN��X��J��틾?���NW�d�Y�.�-"Te���qK�G�����MFr�-��{�����w̺g�:b�V�vO �ZCf�-Q�>׮C^>]��Y���i����M��P�Y �@�{�Y�u��~�d��� >�	�"������9��h��w�=�Hsk)��� ��Z ����?�g"�8~ВG�2�I`���Ű���aIt�q��̄�K�j�)h
����.qn&��A��I-�4�������4�Z%�t\��ᜤ%��Wߦe<B���Ad�}�s�~0X�dL���o* ��pO��S,�xR�\��RQ�@���Pk�ݘ�)-��$_��만:Z�s5!�8Ѝ�?y�:�*��UyU��O9���&�ݑ�̻�^�2w8�0'����D��1��F��[�M�Il۽���R�K��G}YgJ'ԏ�(��g����ߙ��Jm���0w
�D6bo��Y �!�s,�:cF��P�D�Ĩ�LC�T搛�5�����?��x*��c�#F�76���]'<(�f�V�t#���2�9�jv;�x��v����ɤĢ��ou��1b2P�q����x�Ou0SIv#9����[AT�+}>1��w�룟�1i�����_q3.�?���� *��W��k	Yl������8q�k�s�J{���=�c�����t�&9�܄��ZvO-Z���I�V%ށS�~�y�Y@�r��g]O�c68ď9N��igtkӿ�l�i^��t��C��<�"�0š��<@鴲W��E�Zd�*L{��U`�Uut�P�T!�� �aG�5�U-5Od��þ�m��X\@��&9~i�������hqD����)��W�!���,���B/&��(��Z'���p_��z��RSX.�T��TN��*��Z���z�:j\_�2`G�tK7��
���t�
^��'o��0��ID�]Nm�D������� �N�����e#��k?�8쀄�ۇ���L{6��7.�nߊ	F�3:�ԁS��@���b���G]�Z�lk���m�>o�;5A�\���Q�;/(���'�[���uYkr�'BU��W�̊Wl�@|N�<�n/��o�z�u�Uwke�&�8~�ߐ�͞�t�cB��:�coV��H��7��� �u>�zQ���O�a��㬈2�3�\_m).�������eq��y͝���&���;Pl�A�n�������?�e~~���a��-��9C���5j���ԉ����5:$8�f��̓<�1sG����tZ�c�Ž��F�
�����/5�5�`۾l��%����#��a�����۳j:/B����R6	G��΂��[㝶�L�qQ?d�5l�
~H/�sz��9��'����u�dAދ��,���~�v�Kn�M��|��}	�2b����iW���Qm&.�۸����^�r���Y�,��
|7"�p��2�^�}���j�F+q�~�����U��#l��6dZ}~˶�J�>;?3��D��h
����H��ը�e/�l�$����q�xH���F{�L�� �����b�&�vYe���ͨ�;�e
�^O��F��jy��U@{27��kW��v�^0�{ۙ�z���`�Z���1#ҵP���~��C�[qՑ�lB��i��
89˳�X5��@7V7-{��g��,b�?fp#�����.���=�q�U����/K�����ة���%���fC3�E�\MC�Q���e��Rz�Kj�ŰjdR8��Y���
��fH��O�}�S�r"�QMI�1��h�����ߔ��i���<�}gۇ�o�H���m���&�����)�@�ⸯ���v�E����2�|\
�M��ܮ�;�k��}�8��7���%�۩�����.\VMQ<���`o��0��N
g2���'n���.��At�F>d� KF�hA�=+�!ˑ��ip��֬}���M)��:�;23����C��=���ۙf��{��6i�k��M�{��՜
����.�7h��?�lu9H��,�fO3q�V�t�r���QX�F�5�B��H�u���R�D����W�7|�S�+?����惜�Jz���Q���6�r����}�>��I�@_6��F��7:;�
��˃R#�����ދ�3� l<�4�+]�(j|�j�O9��r9���]{���9�砤C��6�Y��S	��X�j��)��SA�>�c�,F�F)�X$�5_Φ���Ġ���x��o��Y�ff��`�����@�UM���y�6��TV�w|c	/to�p�+�t�]�r�����-�Y���7�aL��+D�ٖ��S�|>J�g�|��3�>A�H��k� X�]-}jHB�\ڃ����^�����F�M��D�lw�^r�\�Ac\$j������G����Xo���n�o�+�e��RS:<���V���y%+��$�D�l&���K1���݈ ��
�n��r>x׫@�`�C,q՞o��Mo�3 �9#��1e���O+K_Γ�a�}��~x!!?F��/F�_�X�����ݺ�8N�=S��&o��k��`�?!�Tؗ	)��L��	S�^m���i�X4.b�f�� u��eB�z����0��	�	��V7�˗��0��
L�@��ɗ�*GU��:��3���a��֫��C����gI�
�&/�xMU�:<?��\��k��6��1�͂��͉s�oѠ�o�͒0�M�)L��-l�s��3-]�D�����kE�>?�'{�i�8����CH*t*�� ����Ȭ��jM*�K�r�v��dXJ���	k5���^-R���Պ�~�W(�[�����А@󘦣��%��M�|�Q�ˆuL��ܚ-
�*J5&��;E�$^����&s����'�s�Hd�R��=-e�R������=���[_���yb�;;�y�#�-R���乓]�("F_R\��L�aj���ӂ�����E�0:nL��LP��}��xѲ2VR�@+<�����l���5���ܬ�5ڙ�%�'C�-��p&QV�F�@�4��S��:.3���S�4���9`��aS&Af"�m��/�%�&��F$˿���W�u)��(�g.Q�LE�XC��L~��ù%�9H�..hF��/|��ls��7��ɷ��gf����,�Z��=���\LU^�u�@���9*O>�`d�t�V6���:Y(a����&s��(��ˮO�\&��|���I��W��O@��M����Ub�/"��gD��Ӧk�S�w�B�Qw
}�1Ѿ��#u�[��Ru����⏖&qb�������L�]fl�Y�}��3��U�t!��4������#�7o��V��#�߰�=��%/u%����� QH�ݐĎ
R�}_�
A�o���k��7��g&(4�/��w���Lu騛N����q��&s�	�����qL �Z���?��l���^��2Y#�E+q�/-?x�r�W8ΠD1��rϴ�ӬX��*is��t�ݿ�ߛ���bPhZk�Jj7�⃣|W�Dn|$���ɾc���*#�d��k
k�QN6�w�o�~�#<H/�I��E���k�B�N��r��Z�ߠ�K�:�����{|��th��� �P$<��nvs������ߨ[���� �a�����V�h3uC2�4�]�z��m;��ůX.�b�"Ehf���w�������M-�����s�A�9J�_TM�V���ϧo��>Q�{~�'d�<G,۟�`E���5
��񕞸���M �B�����!�ihȂ���z�.���G�6���\���ղ�Q��C�(��5��К6�	/:��T�0|�&����8�4�I���Jb;��+-w�ç��MɲR��*��X�:��~L��)��h��KT��+C��fXl6�xmE8�:%ˣ0P��@i��{OD�Ҝ��W�\�u��I����[�,�8�
���<�8p.�+���.+Fc�������[���V��݆�����?��_etۚԾG��E�H�eb1��ŧ�ӄ��m:SrDF�� e�W��� �XƔ�۠�Ye<��A����\�£���?F����ui$炚L��@�&"ۙ2��)ޡ�z�vՍ�Hzl:�F��_-��ΑS���@�7a��[hR�]��Tl���/�����~XotBqk���;[OЇzU��w�K�l_�r��x��G!�6��<�wGr���<]�*�I��Α��?��P�5��P��ѫ8z�>����H�0���mEi
^�dVG�ޢ!l�g�/}���8�faB�l&��9T�v}�0�a��紸�)Ø��0ص��iB�}EgTh�xHd���,�J�4��W8|*�zuO3G�r�����=��2q����1Z�}Q#TSu�&��m��C�f��`T������1��t��Q4�=��$/	{�n2�e3$ގ�r�;�l�#F�\�J��S���?P������5~H���Eo�8E�9lf�A98�2?�>+�U[}�*�^E` 崉<��-Y���#�����i�W���� *3�k@�%�/�xf��0�?;���L&�cd�{��Ў�1{1_�8^ϒ[�#~��@�[k_{�\5*���p>c�BEI��F���\��,�sޒVVp�}��E��3WN����Z����g�s����)  x����\ ς9����(�}�x�;ᩪXsp�tB�MѰd ���A��5i5����d�x∸}�sH4�Qpm�BNc��)����6k�T`�A>�Cd:0��'��5G��!�zB�	O��U�4����FS�~�&%������X�G���4���y��0�۽����]@A!҆���g"���dFq���; ��bޣNUa�Efp-��R�6�D!��������=���mb��o!���(b8k+�D{���r1;�(4@,+!�Τ�@��$yQl$�F`8_���Z��
N�DC�f��`�����ݬ��BSǾ�Cz�c0f��u���X�a�B�R��4ʋ_�+rLͳ�����0i��w��L�dO� Ds!A���*-���3������Qi:�t=e:EB���S�n��
�7�Qn��_�e{!�11J��,f�`���ډǡ}��*V�V�G�
W��Z�WCl�m0�޳�H��K����P�pRV�&��0zV�H�84��t��}7A9�^T?:O#O�f5jeA�z����6~�������Փ�r_IT�7a$�(R/�B��z��큶8 �`oa��]��(���kw�JR�H��IS2� M͋0^��1��S���@r�~ݝ�p`j��=}^�BV�SZc����`���(���t�	v����[N:5w ��T����X,��>�� "��h�:�!����+ZU�*����۵�������x��%����Oޱ:�5��*px9�{�v�5�҂�b�����ba!F�f&m�I5y@��[}��I̭V�+�Q������a0�
L�ܢ\:ޣ��k���'��/��0��aj%�"t�u��{g�?�.a�C#�;�䪅ni	�y���NNƕ:Y�b�G��n�y���Y��#Հ��Qy�k�Vh;� �g���$�t~��`�;�A��K�B�c�1D7X��m�n��K�V�9�� r����E��k�Uȱ���w�Q�'�Н?�%/�I��N��s��?^�����}��Ƹ)E�b�C�
Q�[١�G�4c��{w`�1CQ��3q2-s!��P>�MA:N���d��]��׫tߝV��'����0��ĉa��k,b��;�ɯ���z��B�r_ Ch�8c���%�xj�P|�Qڎ�S�S��:kr,gB���(Hy��<l�Ni5l�ο������J�!�G�@\���:x�f�'�X	�B+�\�Pԉ�4ȿn�������	�v{Mn��5��Ts<Nah;8/���i���a��� �~��Gn�щӯt��gLS��W�|B�C;�P�8��?���s�П�+��x��,wa��4m�O���H���r�rʺ�rQZ��j�������:���"�,��>���}��R����`�;�#��ѻ+|�$��T���1M;#~�:�{�Ъ���j]Fa+=� �܇� �?�4���MZx�u"�B�
Zo:=/�I�5�j6����rw��KϾ�B�e�YG�=ڼYC�mEq�lС�Q_�$3����^P	X�ß��am&W�X��l�yEw$�ޗ\r��o�U��Y;���z16%���j�pfc�·ʶ��˽uIs$����`pu�k�{Φ��٢���º���C�G���lb&�M�C��K�:9�b�隯G����k�1�t�ʾ���xS���O��.�|XJ�L[�/�Z>4�"�h����K��dA�3\�	`ed�z9e�aQ������x��AH}��ggᅃ�5X�"�ÿ������J��ᙼf7uM[�$�G���d�p�ѻ�˿�A-����<�.��r����[��JJ4N҉}���K�6��j���58t�"D�n���?�K�Q�9�h�P8�@V�(�xN1�f>Y�4s�.��L�s��"#�Iؿvp�:!�9���Q�q�z�(��˷F�÷���"�PU\ũ�,ByE�V19��F��9��Tc�e��I@Iәs���ni�Ī�s��"�l�:;qe�X�Qb߾�+2�;ib�U��i�� IQţ���,����fk�m({�u��y˨�LC4�1�S�
�9,l3�)�����Q)�����a]5	���J	����E�#x�΃�3�/"�`.��7��a�����&�o4�a�Wݳ�a����o��l_Յ).%:�:��(�+��t �&G�;R[~�T�٩,vP�LN_T�'�*}��^��:�<�:�(L��"��}K�E4.��E����3$FD��4o��0{/�*�E�["I�����4qX�\@�Σ19=���k������k����z2j�l'��ɛ=�vLƿ-�!�,�����9���5�v-儺B˺�Bn�d�M���j?�ف�kz z�~�h�k�,	?y����N��F_V�Ƥ�x�d�WA�0g/��C��g�6��2�C�ai)����9��VxIK�Eh?M���2rKk�tl}.�U�X������zXQX��0BX�?�l���P�w���-ߔ�M�I�N ��#r���ԹV��0Y�j�{*c�';�גb�2�W-��$;ѡ�o��Mb�0(CD"Y�9@e�����9���W�Ye�B`���O��paE��H�h�ʓ�:�$�%
�C���<y� �����.*;r>��icJe�y8!FNnͮ�Z���XCm�`�$�����`B�$`l�ءd{�O�' �%[\P������m'-�82��w���S�~���U��{��g�#�DD��-h>T]��gB7H���?Q~ x�L�ݴ�}�:����NP	+�B?�/m���*���ogA�6�����k2f�.�^!�̗;ն��E��-"�a�.Wwo�!7H��d}���=�r=1mV��'��DϞ�Ҏ�,OX7����P$��m��Ά}R�����[�GB��[�ذ;��F=ß�x�{��
��[��_VH�#׸��[�zg��x�.��y	����P�=�f]
�<+c,���}� �>WO����)n�@�H鳲)�v�/.�d�^�ۋO��|I�is uJC �	�n�&3��?Ȥ�i}�P�����^Z�(=(A#����L��H���A���HZ���ζ��U��->�].�O������6%:r�sp����N~ٶ��)���8�\aT~�r����E�`���\���-~Ps�LQ�|Ki�7���C��f 9��`a(ÃI,<ǭ�m�]cKn^�� �﨑?F~+�4D:����"C2�)�z�����ŝ\�3��8������&�i�=?����V�g�y��
n�r�~�w>���%��TjD�rMό]�8��!�[8n����3��~Y�$���@��q	�0W.�O�1�w�<���6�I����ܢ����/T��j��%D�Q�gZ�O[v�ᦨN���O=�/E�ś�zc5��N^�����, ~�ڞ���n�l;~@ꔩ�<#�V��29�B3X�H sV�1s����`���i[��ʝw&�3z�F'��_0�&$�����]�Ei�R�dP@�*�f���tO6io��{�i&�%��@x{��]����i����,�bM����u��MLQ&K�-p���ұ��f��_����\�U��^�L����J��[K"�'�Y��oc;%�Y�(\�ɖ��*0�$��Ѳ?�o�UԜy�Q�۝�ar��7���V
�o�V9���R�A��D�H��o� �[�l�aa�M ������4��f�`� m)�HM ����#���eZ����	��d��l��UO��q�j�	�O9q�*$M��s�~Ӝ(|~��_�1;��s�+�m�Q�60[j7���h�³ɽ�;����
�
m����Z�EQ��|F�&��F�ld/��A��Wf�y����,�� ן�KyJm�iU]����k
�00-�\�;�`P(LDӅ���ս�ї��cs���W9�[`��<YF��LWcp�����JΗ-���A�L�u��r�8��+oMpf�y�g=;�Vu���kr�^@�g =._t�f݄V7jd�����;vj�!��߆�����zb=��q��Ա+3ͽ��/�3{�{�����=O�Ó5�e�E�&;������]'P�L����T�4s�M 3��_����j��W�=g����TW���}^�è��S�ƉuX&Bތ��F�Ӹ�����x�x��B�������.f��<`��������|Ya��.���\JJ�ȏ��W �ِ��Q�f�����i�����p�ʊ{@�KS&,�_
c��@�H��N�=�ŝ� �����υ�f�z�5��x�h��'�kng�=E�q��3���i�6+"��`��Ô/?W2�M6u��|��] �����5�^�%���<�R)�l���wN�we�����V�m�q a�!�mB?=���9�s׃�f���ʹ���h�dZ�~���	%l<!��<�F�EpST v�`�~���<�s��}Q)�m�¡�x�֐��s��(Lw���]�Z�)�x$^�F=D]�9ĸ��L�nM�:��Oj��d��p �C�^0����$���Y;W�<��6��YĔ��5&Ă; {f1�"����W<�-g�y!�{��\�9���uҁ�%��Hg4-N��~`�������+�I���g�Wx��$Ji�^�8��(���N�#q(�r6�S���ю�q�@���ziS��מ8�Eg�SI�!�����{��̦1]��E��/ct�\�E�@�g��7�i�z�w�W=mM���|x�dVwJ59�,�fa�Ӛ��~���x ��-�F�y���-�B�M�����'���,���z�>%�0�c-� �GGM8�8�5K	����lU�L�^�Lp�%�<z�IO/�;��Ǯ0����n	X˿�14P(OS*���U��gN-�L�c��VJ�$�R0�IŽ����-���lLk�5���� �Z�X��s��M�o'DcU��'������,���??������ɿO�L9FS�����h��դ��dK�d�S�H�`��jp��m@�I��A�:�Gz��<ٶ��d:��R��"]l8�5/��\���/����"$cܘ�;��ϧ�T�'�r�U��x^�>�s3�f�6�b�X�C�5k%���웳)��]�ƛ��`��j}%s;nV��<��g��
>��������L��-�`H\��0&���MG�Uˀ��}�Nv�$�9 �����kv�>[3�m�+���G�h7����ꡇ��U�*'T�Ɓ4�S9�a?�I��5S�u�Ý�=��^���Q�w)D���-��at�"[���@��ay�5.���|J8�$���`+�U�F�Հ��ܴP�[��ݶCH�N]��9�2��i�NǱ���v8�u�[��`�@���J�p���4%�ϧ1úź���^e.�j:�.M>1HYb/�tr`�$�A:H�;n��|��}1\���+�u�^mc�W	���rm�PH��\"M�b���Ye���|���V�ԫ�r�v-��|� �5p��Mq�q���lը��Ky ��q*M���';����90t�
��-�K
�߯4of�6qm%&8���Fëh���d��Bޮ��tb�p���s?�+�=�W`�ߐj�ǔ,�NG��H�p
a5]�����.��=��"�e���� I�䕪�X
�.J�@ho����5yP�2@vn��R�����kb������O��*R%ځ�"���;W�5����~�]s��Jmh�KT�%����@K��".V�=�eƭ�H�~�m���F(���$��>Lu�_z&3J�o��;����1�x�l��s��^7�:��w�&b	8�b� ~�{6�X=a�q`V���{�
���N������~Q!��-²#
� S�1�,�,e�X��:H����]=X���~�d��H.�ihb���e\^��lw�aTH��|==��/��hm]�r0��k?��"Pe{�=6Q�������:��^wT�m�6��{7��F�(��B�W��ͷL_��5�+���g��S���a0N�f�w�֦�_�=�2���G�.��H�9Iٻ�ދ3�=C�:VYo+i.PE�4q�8,�/-��Wg�<�����@�g�y�2�{N�Pe~�c�r��{E��W�=��gD�7{ꀊ�!j0�H-Ü�v��Ⴓ�!��b��{�&^/�����<���6����l�ؓ�H|0g���n�gMx^G0)���E�ʏj~p�_�h"9��d`9�{2���Y�s��OHLaʫ��g�s���-B����)YZyY��Y�[tM�m��X�����:49�D�qNkGT�8e�p��|N��I��Q�z㾕����-�Q傤�ߡQ�j��S,MT�rIO����0.GLd�F���7�*�m��|�a��1M�w�>����1ڥ�@-ZGDV�I�f4���;���q��!�T4s~��i�{�<�'�[��|'.�F�m!.��-�b��R�ib�V_��U��8o<P���O���n���WY[5zl^�	�X90R�_��u 2K�-�_��q�2'����3m1{K� ��w����<A��� ��)��%�D������_Jv$h���+=S;�6�X@X�q�$����-*��[�)���E���u�����n�b����5b�w:��w�~���Z�*Nˁ����C�l�#�O	.�y����HW�ζx�֩�Z�Ӈ��+�w����a�~h�3}��.	�݇�r� e>snƁH�
Mr�/�gW�̹�8s�y����#P~_���އ�C	f��`��.CQ����^Vw�{�X�xIƃ��L�qet����7߈A��C��\Zo�̿.�\�/j�jiH�϶����8���j)�,W'ߵ1���3�q���3�iɔX2�O����ְN�
�U��Խ R޷W�5�ޭw����������1�S���O}zr�F�z���nB?�D�M�]�h��������%;�!�vw�7���"�� ��"�.�[�4T:=@��S
(*|�,���Gװ���,�� �\��u��@u��J��fJf�j)-|f����6]��/�j���8}Q�3��i�UT���J�3���+;�4�'��c��N�O���72ƭ���.W�AM8����}�T� ^�&w�v:)�ߞ�Z�[Zc_�K��M�����4[Mk}*��ƶ��\#�G���Zg��T���*n ���ln� ���,=؇m�d��������ه+�`�e�I����i°U���������>�:f�}��}.ʶ�_�%!ŏ���N��a���w/]m�#������UvK���c�L\q���d���	�/;��W��W]�B�=�`N��0y1%�?��OL�?�E����4� ���PM�fI�m����(��v� �3��TQ;��@�ƿ�e�C�T�;��\�D#��%5���>	P���W�zz�U�-�F�l�݊:��x,��f] $�|�L��s\b\��]����i�W������*�I��3Q@$]�L�}�TI=>��=��79�+�;�U]��_�1�{t-^3C&�n�끐����5_)Bl���_:N����"*�ו8$�}v�.l�,������V$2�@�n���!?��9��Zi=$�vE�;ݑ���o�����?"�V&�E	����c����"2:�zz�w!�(=�`zq��S\��٫ϺlH���w��&%v�Ϛ ]]β�Y�\�tPv���Ak�+��W�qqڎ��!�jhP1����4A�i����mw��v�fD��'8�? bK?���d�����.�Z�"߸Ia'���^�*��\�E��e0k��*{ynN^R�G�߼�܋;��)��TYٴ���&�y&�[�X߬���5�+ �Q���:�v"�-��!�\�zM��������Re���;l��냑�K��Sja�2�
�[Q�������C��Zx����y�R=JT����$�������g4ύ�4v�x1�m�iA�<`m��7�w�?F^� ����R	v~�%��=I��X��ɽ$x0���d�(û�mG��%I������o>��h���yEp#l\6 8׫�U�:�G{s*0��/�x9rcsT���=w���J���hC�5C.���hY)؇�ȝ��k�\�Er*��r؜����10V ��V�T�`�^à!�:aa�Hk�����J��á\AE0=_k�RCb����2bE;�`��!�S�H���D�yea:��E�lVFf5�'�=��oI��/�X�������jg�VK)��EU��I\O5�D��)L��7͝����/�G��'3}U\q�I����U���S��1��b'�����կ��f��ɼӱm(����o�r�hp��~�(#����B�N��	T�+A=sDpg3TVn����ً�`�4�`I�僧Yɢ��'5�P	�T�qZ��u�UJ'dcZ���	�k�	�A���P�9&Զ��y��'a�
s\�܅��tb��
��s5���T�׍��,��ɾ��á�������˻�9T���(46r��0~QC�j��$�*��U+Vu,8l�Xe����E㱐�ز�{��fuŮ��n)�l�&~pY�ĐϊT�lJ�����������2���)�L��OQt ��e�NR�I�!��y���{ynW�y)Һ6g���>Wu^t�י�F��6&O\�=�2łm9b;�3v�4tۡ�d��b��W2�H�m�Jj�����U��G�@ۿxyM�jH+�����za�����6����ȵ���5�q�i��$�Z��m�l���P�#�E��� {�Zf�׸#3LB��ʇ� $����g���b�e��%7��X�/�����6�L��׎�#��3�1�����P�mąQ�-�^\	���kXm�=5E%�g��#�$c��<�'�I�|ۇ��K�|���չD�>!X]�c��]���2�`��ҥ<��*���lđ��=�~rZ�G�������Nƥ�!��ጨ�#GQj��YMA�zW�3R��}ķ۠6^�J�Q]�O<��풂�E�@⼾ȥ�2��� �Y�m"��"������;�x�|eq�W�/��C���h.�W/��z��x^�+fP��Q���	)�$�����yZ�"��-�F�h�e������R�p�l?7�Ѣ@1�� �^z�A��/c��7f}�n��$�v�p�?�7t��6��⬥p�f^���r�5[���~Je)�&�Y�aA,<�>*���e����H�N(Ҹ�d�'C~f�iQc�?��^����L�� �� ���� !�oE������;�(��}�Y#�!`��������p�Ґ��T� ;�Y@EZ�j�����b����Q���8��@�8��;+�Z��p	�@AW<u�7��{A���5�S"�/�ș0�|� PvG����c�[��奅v��ɚ��1l�~��2-�;�.��>�eu�tn�n)�R�i�eP��}�BuZ��ʵ�C�B�l�Z�ty�uKn!lm��d�C�
Vm��_�J��U6(����~����"�U��x�V0YW�S�4�xQ����u&�͚B�~.ُC<{T�m}S-��4��$��hN�b�?�q�Q#NL��ꁘҶ��Q�����9�!��<�H��X�}���+iKd��op��|IVG��7c��vb|���5�ԇ.c����i4j_ef�U�V��R�P맦��$?�9�#��q)m�^�� %
�5g��#@<봡x�;M_���i'~\Ir�-��O	3{_�n��A@o]�ś�g���ziS�ᓹ�Ѕtvc=��!�+�hlo�p^�G�3���V}Y�z���v�+��s�,�Ϯy���0�vS(�p�>�o`l�P�Զ���5A'eљ�����I��uh9d�yT �,�p$-���s$��S8X��_��.���kd$Cd����:��-�ng�{l�ոXNP���i�q6��yǡ=�u�Bn1�P�c�#����,2+b���oY�-�W�,�y�'�QI��)-b9������U�g����t���N��e�~U��P�:r����ԝi	����Ԟ�E	3[�����QqpȲ�f�lv+yR\���V����+;�Ͱ���u��L��fy0^�&�=)8��]��=�����B�+I7��� H��ceH��𞶍&���s��_�]lՏ(�T61���[�m���pF���M��w��ʶ���R1p6���ٰ:��KIٖOjUE����s��	��ե���)N;�G�r��M:gTw[n\�Q��,:���Ή][l�L*����ŏ0��o�qy���ľF�.�%w��%��5xߋ�̤Xl�=�x>��H�Վ�Av���^����*��,�Q$۬ΔWS6�A䩱��>�s�������~=p��)^�>ѥ�����;��������Y�yRb��@T��x���GQw��N��Z]�!� �וS]h�� ��G��@�h!��]��܍�ݥ���]:d�b�.4��y!؆�~�v�Q���_Fy��
<���ŭ1jT8@�qD3�_��
&UO�.�8��ϵ/�Z�J���>$|���P�bd	W�93��p��Hփ�J%UGE��P|_����]ڡ��A[�X�0@���8������� @3sӡ��af6�b��5{�q���h��R���iLR�։��^�^_�lb��2}�	#�T�#'�/ �[�[�_�z� /�?g7o�z��=޴��������Ϋ�_�&�k�}�Y�̴�a*��h�T�_������&��(n�B�ZM-Ke!�OAB��D������^c�+��G��D��}���	�vbĻݸW�B��֧k��"��l{�Q������������c�I�S�+Z>�/錛Z�m|fR�;�i��D~��l��3J����b�0m�k�^�X��/zwd��;
�%i����p���8����_�y��;Y(y��ue&	�hr{\.W��:/4n��A �4փD
����d��]@L��#
�Y|9�����$�#{�re��,�n?X\#`a��/�:�Yy�(Bq~�³�pT�z0x�(���B���{������'��B�R�}X�/[hB�ySk���H�\��(���sr�B���`B�=�8v�	�s�)"�6O5��ʣ�*Ou�#p���[૦�oPｘẮ����"�xnDC|�z��'#���߂���>��Jc�b�(����ģ�Vqk�)���Ҫ.,`� UH48|�E}�M�ĺ��qb䱰�#��<�o��s&A� ���c��uWc@|<Rȹ�]�:gcN��c�����Q���fȊA���Ԝ��H�иl�B�x^/��&R��INc��|��u��@_�~_�Ԩo�uVQ&<���7}�p�Aؿ_�E�Pzj�F\`�P���Ba4�u��\.������/�����6f��A��Γi#G}�a�Q��%�_�#��I��6���;��S+�m�'�x#��X�t��f�@I?@�$='p
�'ރa����C����D���FӃ���%>��$J��J�fE'�@�,f����.֞L��әe9ɋUe�:<792<~\nx
u( +>�~ѝ�TȰf&FI0�W h��!<�\Ұ��*|2�g�۸(!g�
��ȶ4�I6"(�}qp ʴ���T����W�����0$�A[�w���kV�q�M��A*�8z{�PdFy��'W! �S���2q�����P���	׳]�}�%������X�l]Um+��,�%/k��#H�Ѧ�Z��y�0���B*vC�l{�®���X!6(`@���)(u��TG�:>Ѹ���B��j�? 0
(�����a�Y�Q�i}o\�ה�2��fDr�az�]$\\�� �~+@�mL�p��A�V1�Lc�VД����jl���ہS<C�IH�l���D���2��$�w��S�6hب�l�g��fLP����?{�kMEv�Fe�d��t{ Ȥu��D# �A'���1i��N7�;��kG�9�ٝ�]b"@�>��I�ڼ�!�s�b�:r�>�+�GDT!�ODBr��'�	hIϜ��$��8�L�R��_�|N�)�
�#�Ï���DU���S󏦙��K�9<�L�?X��k4�$��c�H��1Iu�?�0��Z��y�52�b)8�W�*�Y�]�<�r|����/
�}Z���������Z�b�Ū��V�=���O�dmeEW���\�\#dLcj�6��	Χ=�� ��ݽ}����Ֆ�^�Md3B��cy��\���7B����ĲZO��l���E�޹�D�!!I����\��bI ��[�1\�G�G�*��H�iF�jK���։N�l��1M�E�'���r��:�È�r(:��xϘ� �� �u�@�����^�դ��(��1-�G��>;ؠ?��'��E��/Z�z�1�ĸ���ݨ��}�	�"/�=�h����E
]P2ǥBw�Q�G/�t��ٻ��G�ޜ:D��ˬgUٟ�سV{�6���>�!��PO�6���K�����Ņ�Z��$�+�l�i�����ܔ�[�GX��qGg���j�a�%n��O@���^�F�@۞V9r�C��4�bU�ES|�7g}���P4�c���rl�#�V����/�9��ޅ*�M�S���-��"/%j≯�#�0�>�G�܀!�`[�N-�gm��
|���ebƯ ���jEKB'Q�,*�F	��9t��WF����Ī�tI���h��J/W&c��`�yڳ���<@�uR�][j�~0��V 4�$���P����pҘ�+￾�p���Q֙�/���2ta�Ø��m�p�W�3 ���]�M��q�T��v�G�vԟ��e�[Y:���e�{3�ϱiXs���b+�n:	��K�����o���j�g@!��Pt�@�b�[���x��`L�� C�������&��en�=��E���np�_���+��tS��N��IT]��b��)��u�[�O�=Iҧ���3�:LIi�=�̓5�n�2���TΈ�W�� 0T�5��Q����OG���;�sFM\-;��l���
B"��4�>i혅h�!����Y��� "Y�v���47�	^Y�|�-�>9�@�CUX��C��Qt�s��f��1$�^8�|l?�b�F7z��@k��4ةX�1���n�9�L�<�r����Ja�a0��\0�#��+�1s��l��v�Jף�"�
������'�)���2��#��;C��]�vڑ�@��b�;��W�Z#�+F�3�*�/�&��h�S����v�<qgW��`�2p��ⰬD�giDWn.�WPTR�6�$�"�;�G�:���c�%0a�ZV}2a�P�1e�IZc���U��2�J�e}ŗ���ڋ"�.���4F��v{��T����&��9��3�P�-@��[d��0,�^�ly����
ŭ����墩K��2��3����4��M4������pF�@�ź�uꨧ=�����]~+xB���H�=;I؍��1F�.�L��8hY��.vb�]�C�y�#1�cp��4܈�k��LhGP>{7� ��O̮�9X����I,!�osߐ`���հ1~�^w��{A�:$Kbznp���+�� Vv5�v^�H��s�iO7���^��h�;�
��2�0�*��V�Bt��Z4��D��\�~�j@�ih0<�n���c6IA��Z`Oig~�%��JԎ֪��dɂ��B����'������z|I��}m�fl�ւ!�6 }�(�șb@����ԷF`bw��!� �[������P�q�<�]\|��@)���d�6i�7����W��و��ue�@�ukRX���Uc�yA�����x�0K����G�ҁN�I�&J��_F��wW~��=��	l�
;3�T$2DtpA�
GF}-�,��]��Vܳ3a�:A�ѻN�_��B�zV�e�N�YҾ`&�;S�Y�jEV�g��d5�dS�9�b�K���E���@{�ɗ}�����������^>�
R5B����kY��C<�/�p@��>둒w���f����pX�D8{b\8A�&٥'a�kq�.��p��0Fp����#*s�)AEh)���Y�b\�@GFl�V��fg�?1�H�0̜�恥�/�?3���{Uo���h��c�7��g�b8C����	FL+OG�è��J���sg'�w�<�}r	R���'���I����ٛ��n�SX��v��68��KO~��|��L��9!��lҍ��_G�9eS�p������lǆ.����zX���ʘ����he%���%��. =����`��	9/��{OiA�A��е��fm�ۃC�K�!Ɲ�\#g��{zb���@C�J�t�/"�r7%Z�/ X�,Ϡ4��p��H��s��r=>@@�Ϝ��"	����V�)v�	(�S�l55��Ԝ��uG򳮽͵��ih=���5cN��wT��	`&ɩ=+['����b�S[��B�H��t��z0Uc��@LH�ڱɋ"������/�;��H� �����6�kq,�����1������˶L���ڞkt��N�7�/T|�ڒ�K�Z~aQaC�]*���UpРJ��dPV&����5�"^�m���1���͏��.?�p�>�=�^Q]�rA���n�6�+z/�~�!��Y=+�j�':Y�Ţ��s]����
l�J�	��0GG�y��zKS��))��r��!�7����A�I_#��-�N�H��X2�Q��w���k3��ŗ`�ƒ����G��u�q�E��ׇq��H���]-���I{P�Qɧí�f���Kw���%4O�����~�X#&}l�+*I�3�c����E�U��t��>����fU������Qy�0>K6n�.�FI����Ck��N��T��l��!tO�'6��	4��J^�_I ��H�� ��H���{-F���ٴ%�&m�D�R=�&N�����E��ni�̈vS�����7+"3-��_��Nj���s�7�l@{�*{1�'D�С�
��/@
���C�&�(YSF�-�L.j�Κ:w�_�`�a�hGǧ��%�D�b��ZA�+��Q��h@��fA	09>� G!h���k�y��TÅI�$�1�]�K�_�u�MJJ]�zr���9�%LfN�@��΅�X��t��DI�$�nc呝PD�^Y���}+k�Qì�˘��a{�_xAs�����Oa�K�� ����3.�C���J�|3�bf��l̰�s�]�&�X
�=r�oо�/�Ҕ� `{Juj0��6]�sh�x�����Q��U�l6�V��+�tym8h��������W1�zi����r�(	��H���P����a��E*��p+���Ar��6vP*�D��@�16 ��e[��F15����`�����#17�vW��8b�A�s0c�>o(x��#��l��^���.:�B�0ߧj�bR$�Z���cG<6��f�d�g��:h��D�0<�g�H陼�mp�����y��M�7Kl�2l��*AE#R��닠ܬp�����m��&�-4ַl��6i�r�
�$(�u��_D6�-�����c��*`b�--Gqz���f�ǳ�靍Y.X�77�w�-�&���e�a̅���7�n ɹM�4�:"����8��6�X�o�Cl=X�ۍ�q��	���:��#�c&��^E��e����G���no���!��K٫}�W���ء	2;�v�6yv�cDaq���AF�-�Y�g�Y���5`��a�x^߅��;���1ܧ�~5��MH7'l�
��:gX��'�%��_�0u����=�>E�0���z��4e��v���+8�5mNؔ6���ya(�!Ƥv�w��`���)�z�_.��wf�a�Y����Ơ��s�ؔ��L/z��y�pр7�O�1�2I��m"7�g�7W
���ӻ�ㅦ�����t햚��OH7xrm�|��O��wd�6�+$��s�g/)�5D����]�w����T�+�O֓�Q���K{���>�=�?�k��藶��xm<#(�$��<��1�}Dא<��0�g���\��0r)�&����bx��	6_��y�/����L����Ѹt���b�D����b:�K�t�f%�Z��@>���9��}Yޛg�>K����ۤq��?J���)�_ѭ�a��`�9S����.��>�Sg��OTm(�y�x\���֢GN+I���[8{�
v@ȞE�}K:�q�{T�nK�e���iuвt���g	^:�)\�W������&Чm#6a6Y���ͥ쩏!��a��B���!�G{h>J`��6ۘ@1Z�;-&I�-mٞ$�r���e��6o���=�[��<3C0mf6 ����d�\��� k���j�F6V͚�$ɡ���_~l�A���""���ŀ���߻�&��MxQhC^��ü�:�x� �W*�W���E�+I���s���	�g��YY�/�T2g��]��[S�#�8^WH-o��4"�^/x�/=7�8h��" }��^�� <�lƅ�qJik�| V��ZƊͅKW��/*i/o��M%����q�.�,���+�H�� ~��(m�������(�8A�Oud�����9�����ϵ�j�㝙p �C��4�n!/q�����dqD� ����Q���tԆcɜӴ�Cܢ��W3[��-�Ű=���e)}R]��s= ��AѶ~"pSmk����gn������/����6F��V����w��S&�B�UC�|v��p����&�'Cr=T�z0����6���冪���4D9��s�H^e7,���=��vprR,B1�䙄�:���Өޙ��)AE��q[��p"ȅb���kC�/E{��JӍ���i��[&�������.C<������>5�p�S&ǰ6$Wz&�B�aչn+�~.� ��>���F{��Q�\�e�v��鱁0n�Fdr��^"!_a���ۇn�:ss.gI�l��8�g7���@4fq�n��&�K�]��{�A��B���:��%�=����2���A�6�&܎j���S�	�3����Z;t�_�C�2���1�L+��2����U�D���&��
\�<폼�ؿ��L���\�r���L��|�����"x�]�N��	B�!�24��uȼ�HM�)� 3_Gx��`V Ts��B��L�W�'}�[��7�k��p̒��Ir%Z����Q;��s��lO4$�CU%��w%�mt.+�U��+�ܿp�W�8�n�f	��*?Z��9�,ܛ�Ӯ?r�o�Q<��ۚ�ɿ�IU��*4'
?1洒R�]���.����W���Y�oI�+��?+�]��U��L5k�p�vX���A����?��+���5�Q�^���҂Pu݉N^i�f�S�+$���Xg���-�*%�����ݭ���	@K���ߞ9�f8Jk*��ՅD3���ŬSp��)��'�ؚ�7po�����}��S�Da
�1�sY%�9:z#A'�I@$�?�9�w���,֕�Q�$ǡ]O��|��Q����W7(k�z7oQ)���.�kN��S1<6V-3�\��t�y�>��0ת�_fڢu1i(�h��C[��x�Nz����ʥ`��9�cY��A���Ћ�)�@K����Q�i[ح[�UWN�"V�A�e�7_������TIp�yӊZׇ~ ؊��j�YkAI�&;F��U:���V��,W�p�T�39]�O*�e(�mE�޲��,Z�WW);�����?�z�D����Dg�1B�p��&[��dfliY���yEmI���:�*g��X��\A}p�s
�3NW�.�6,
��	/�eP�~�� ��a�x
?�,�FNh%��J`� +#~�����,h���@Q�#��KjFRw��ea�i��R$<�����aV�w� ��lo����Ci~������ ��;��S�n\�u|��?9��U�M�3|��5��+MC���yi]��U�θ��:�N�%_�9[��/�������{ry2*ݙ��'��Ph�2��A���M٬��H��1;�2+.s��S0kDkA�26;k,x�9)'$����T��H���$h�A~�q�}��-K�8��&�Ort_%Uli���"�de/.ĭ�M�d�Ӣ�H��5���+���`l��f�����x�p0�@oV���<����^�܍��p�_�~�k�Yd�3d��rDé�6��P����.rnA{�#�Mz��٠��m}��fT�ߣ�*�Ȧa��A@��!a�R�j̞������v��S����z���X��H�"��m�{�a%�:�^8dз9�C�w)�V���/�g)4��lӲT�`\Qqr�$Cl7x}�Ꭲ��(���c,`�u@�=����8MFMY�%c�/�7n��)��^��5w��a�����E�����C�'W�;���ƫ�o/�W�)��!�8�.}oGl��bu�_lϰ��y��)~R��u�hއ�_%?����EjƂ�0�A%���*��#�1 2`:��#��n��B��PC�^1�@BFT�g�Im-�,�D�b�0�O{1UdM���ٸ/��� 60�?T|��O]�����.�g#��jS
h�4Y�D6�J���!"T*㫏r�M������ͯo�9����/k����@=��0`�@*ǧ�e�����]+��kl�/��	�:�)z~9o��E��ܫ�I�Z����G���b ��� �4�����4�������:�Y�ݼ�d���g/9Ux��Œ̗��a�<yk�W�X�:ܯ}Qټ�)��<� �L����m��D�}�]�\���N"?��Q�<�y�r�Ȩ}��R�5/�X�hjZJ-LK��|�[c�0GK'.�y�	����:��Q|K�%�BP�p��W�"��;�%�dy���j�}�K����h���J9T*�q�U�X.(x��%��`���8��n@T�2�t��JRq�0p^(��R��g����2�O�Y����oMZN-1�XwY�1V�M����[��j}t��=��	+�}�2%y�R�ƿ�Ւ	J�r �ǡ�|��}�Ev�����zֽ�ޱ��Tv�l����K���؀�Uv촽D�M�9�0B�m��>�I+'����Wo@?;� �U��Q��)C�,�_Z��<�M�OGz��2U�/��:$1ɓ���E��Y ��?E ����g]H)����((xZ�>��R^y�5=Q�,o�`��=�y��u٥���"�T�o���l�%��紀�`���	���}|wN�3����j�&*��ւ��1��-�wkZ��X�j�
�9`Q�M��;��Q ׹�lBI�𒼝�N!���/U<�V*�EI@�b�-�Gd�-�a��gs��)n���b�R�X�'�	P(궴=����jy�zC�
�7��^ۚy�9-bz,R��k7�=��E�[]�ȟ���h�G�y�.����3�}h��.�n7�1	�iU+a��nʚ���5�x;`�B�Sۙ�]���5�	.����R��Y�@��:-Al���Eeͅ�탳�v��\�t�.�x4
��0�\4�|��ؽG�a^��܍7�����l\�MLk^N�U,3��y�G���
бU��$��O0�d�i��@�]Uܿ��q<|�k�Hā2����-��B�(�<��4��j��W��v��T�џ�n�S�n���fi*�;�ed>Q�^���GM��ۃ[WN|����:�^��V�����4���
[5j��<����K����}��3Ҏ�6���}��,;�T�֧B����1�3}
��?W��k"��O�v�������#�D�̧v�V�
9��hb�iH'��03�c�}1���Z)���J�xM��:$18uT>��~�R� ��Sj�/�X�9�C�4/�_\~��=��\�JD6@�\SR�`K��]pJ���f'��.��ߴؔ\Vk�٭L�(y��s�;ӧJ+��ݰث�E3�'�T���3N��|�Jb��{��`$�ƹH�f�W�ʘxvI:�D2e���tTjN.cс���&L���Y��Ќo��Zac�@��I8~�#��N�E���\���l�ͣ������hB��iv��������h9�0�������Z��m���c�`��AM���� k0�(���[aid�-��q����l���i��i�0c������ly Ul�0� ��
Ѳ�F���������ڊ������o��x܌���Ћ���.N��2N��:@q��sn�?�C�o�4��<����"e��f�&�د��qG�E֚��b
38�2�y䃇�u�c<0WDR��i�~Ԡ���Ȓ�{��P��.��)�E9�ś3��6
�P͗��Tޗ��S[s�����{���f��u�6 d�0l�n�ᴻ)�&������7���:?��C�tO}1F{K@��y��\���?&W��>��#XH���9H�`�F��z8�,��8�ų�9�Ⰾ`����v��yf"!����a"�ĥjq��O��`{�A��LC�����h��6��`D- *��uQ�KIgrQ��#�=�v�1>+���x��'�3�~?�+Oτ� ��AL���AfNr͛H��6�O���UX/��[1C�m��l�S��[�ϭ���?��0d�ly3�{����)/-�����i��y��#��h����P!��WCQ�k�;�C����r@d�4����vM!�pzY�p���)CA�[x�Hl�&�4���+��39X��n���2��t�ø���HyD �f�'rfc��̹!uEҚ��=Zɢ��$C�#?G6Q�^�������c"�����?���ᒮ�������|&�#\z]P�@+�*%�����������Y}��+��`?Y�Q��=@�wTQp��!���X�N������PxM�T � ����ة�����G�%�����`�69kk�x?�� X��v�@W��Z���bڟ�	�a�ɐ�.; ����d��� �L�lv����pe�8�6��o�,�Aһ��S.�p��Y��z��4$b��F�ȅb]O�b��6��8���g�_1�%د�D\�r�dR���ް���"�N�Q�m���s��?g��q`b*��Q���w~A~ga�F����VC�h�::��G���9�D�Z�z���a_� 2�X8WF3�8#ݨ��OW�죔=(�p�g�=�����A�B���w�3t,����a��!MM4쉴��I��J���P����=�N`y�Iy2�o��c�DʑY~��/��T�aEỲ�����k�L��4��������b`�a��=�}�-+H˻�6�l�.~֛]Ԕ)$qhj����~PN������}���.뭔������Ü�c��������6�|U�_��_����l�D<�bljx����̡����: �$?|GЭN�O���?JX��B�m�~k�%KZ������E2�W�����E%�푪����Tq�TB'�^�XA1�П�l�ԧAYF�s�-�����}R+	8=�-Ӥ�Q2ԃs�� �h��"�&Պ�O�c���Ω�,�C�?�kh�6�@��Κ���$���J�e{6̩ggZ����_���$w&}b���ɿ����0�LY��Dj�;q���%<��A"��C�����T�%G�Ա�S�THL�ܪS1#�$�Ѥxo)]x��s�T����:�̣��q:ޓ�r��L�$��Ye��ƪ���r�����b�$i
) �i�����At���G���3��`�Y�cv��y?�銼���o]y;ϸדט_����^_�e~�v��� �N��v�Ր�����Y�덻2�{��g�1���<qz�%6�1�<�{�B��Kd!�Er�^����?�'n5C�"N�I�*���_�,����]�A2�z ;���tۯ�h�E�Χf�DaW%Wt��M�ݜ_դf�'� �rj������W����E�v͠u�i�~N��I����b�E��j�UA���RE���%Jv旗z�����*�D�W ��{��ʍF���=(�}��a���jn�ƣ�oMb��q����3��Ɇ������=`�$��vU�$\<�7J���d*J����U���s��⢌Io�b�a�9>�("/r5�*�%���w��_�I��n�V7A^`�}w�K����_�o�\�""�Y���Rz�$(��P$�l�M�S`K�Y��'hϮ/�{��ǽ�ȁ,�s#y:��7�x��v��&�lk(bo�c����<�%'I©س&ɺA�m��e���_�/y���9e7��K����:��s���e���Vn���Hwj��C|Ept+�2���"�[���J1����&�9����~>Y�)�>+�+̿0�qx��� ۰�����\w��y�:�G�5�W���
�[_X�������ABuK�WaZM�K,���7����Hp����kpϖSb�9�G\+U#k	��=+�DE����PC'K @��D��#t�n����2O�?FX�i�{
.��e���
�$|2)Y�����;�=ᒠj��&s��}��6t-�YR�_�.�{$�b�\���'D�����I��G��T���ʴ���(�1
�(�ͻƸ�<n��)��O�k^��A�*{�,u��1NQ�8V5R��1"�� �Om&�=��bRO�mM�9��w6�,����vM���	%n����@���/ۺ�1�NA[���l�����҈"&�o˥3��X�J�(���h����4��'���P0�k�t^�f�M���/���nGq�6��7�x���a�� ��e�F�_dK����?ʠt�#��)���ΩSE�ǼҦZx��������x�����N������dO���j4����#� $Q<��MŽ�����G�M� �B_nKݱ�uI�{s^���$ |~r�r��Ļ�^6rr+N�Cbѹ�cl�s\�!U��H��8��V��9���w㉵ڹ�t{`7�葮
��Ɉ&�N��F��=�ƺ��Dr Jg��Pg�j0��U���0
�O6L���xK�Dǟ�x_�#��~��hLwxݖw^�I��vw���@�V	瘃��⮄>Bv��/x�΁�4��wدwݘ�2�/���?�����c��3���ڃ�M,��6G,�~��חD
E)/�&�V�M,|�G:��s9[ZH�uuͫmj��[�]b�/Pvl�Yk,j��h?��O\�p�,t�h��A���ʛL��`)~�(�~2��]h�U�̈́�}�"��Kv4��n��D�~X� ���f7�#(�k�bPc��A�;��;�H�G�+B>��`����L����)Ɣ	����d��2Ƙ���4�L�h��E|u�bY�-�0�ij@k�PD��[p�8+_5uS&�6c.ĖO�<�̺ǣ�@�n��J��}*#��Lҋ�?*>��/��m����ɽ�8�(�D_o�!�F#rY��]��z��b��/�֥ͫ쩷5���}��f%l���}w3����m.��A �j�̔��?i��}_q�*���58_��屮%��xNh��`��kt,曗u�P�^�e���(G �g_�id-�#�ǣ/SX�J�b�P:�� �M+��ދO~фX�T��3p�����$�|�k�KT!je�TY���qE�1�X*d�����h�E'�j�"I)�O̯�^�Z����6@o۹��nxźxJavFdҫҡ�Y��B�A����Sa�
[.�ktZ�O�-��Y@�hOHww�{A4��VU�н����[?P�Iϴ��>��*�t���[����jA�_�4Sj���tU&��mf�W���{�����4��`W�H�Ft�y������U9��@\�%"�9������%맧��e�@ߡ�@v*+�������D��6�jg�����<賑�����r\	�Q]SMb:���Ȳ�N=d�M�ƐOm�тS� n.iw��R���0�z��lr"([� �v:'O�V*����� �[Aى�$;Mi7d�p��4�P|�y��v��F�~�U�u�]�M��M�B8S#�طfs�f�YV��)�v����Uzj�e����R�g� ��Gc�ۘ1nQ����N}6�ˠ��V��+��i���PE�ߞ�#��lZ�`\k~cG�g��ZGCc�$
d�ࡠ�݅��ž�&m��t:�5��� �2;�&��c��P���_����]�7���"�Ը �e�C�q�O ^��3��Z2�S�v'��P���8��>����R�lA�U�m*������"��<:^���x�9��ă�SO��98���PL�8CRD�\y@�?�db��N{\�h�����?Q.TԠ�nǫ�"�F!�B���� �] ����5a���jN�@���(�����'=���t�i �+�g~�7�p �q��T�{S�:��Ý��'�1$G�X��"?g��g:�u��Ã��T_0��mﺾ%�j}{����'�{��B^*߮���-��RI�a�U΂|)Ǫ�o- ���'���}[vUA����U��2��~��\"�@)]��L��c�!���!��8S�%>���X�jT��>�9��`vY�ƈ�1��1,�F|���\b4����".�m<q%�o6��j`@R]��k*��b�A(���7����4��O5�^�)�4�6l��ٶU��O�����s�H�������Hm4�"�<ʤw1�:<A�`p��.�˄�ޱ�ѵ�����6��y����)!��Ж�}\@8LJɥ{X�jg�����l�-�LQ}F5��B���������)�`e| �KG��<��S_���%<�<�vrH}���P�js�}t�.�����\e�-ш��M�+]���{��_L��v?�����Yc���+l[����>E����R�K��t�x(�r�Ω%̀�Z$.�AF�r�o�#Z��g-�<WNG��ȶ���	v�,^,�W1�O'w���q/��|k�R+q�܁�/ ��~~��L������v�����F�#@�#����B�t���0K۞�cKu�Edt����_7��;=Ȉ��t�[S}aF����)�N8]C���a��t����.�Y]P��(u���*nUO{�4,�ʐ�L+n`Q�p�w[�%���=�ڠ$-pqm���<�|�Bb|O��[�����|�����U��q��!bB*»gpP�yhZ��S�Z�����;�����.�Ԋ�!y�F�kB�t��>0U?r֣p
�3Z�ު��xB����f6[�&J��[��������뻥	tK�0��@v�>>�8N"�mP��Z���x�����|-��_��"gD����hJ�cd��
I �N�c���o<�MwW��יT��� 2���jG��N��&��"�1�q1���#�8	)��A:��<����'��޳9n?�g?�����)��>�� �Xy��x@�	5�<|����PO{���%7�+4[4�jd�[��RVg3C�`r������b�����B��d&�ԍ���8�"�˪ �1#�<��!�I~��O_t$�,��5��c7��!���,E`�:H��0Y�%U&���Ѥq�A_s� �L��r?{@�)��=
��V���ό�7�Bf���uң_��m�����|��ud[j�X����Ȗ���l��<G�G�� �Ђ����
�ܘ#�K���+^#�,�5�&I<�`b�a��-	�߽ �`]\d<��x�V��9��=C{���8M,���]��M� ���8ߜ�m_�p�[���H�C��������9R3#�q1iLP��r�&Q�(9B�gn�b�/���庆�=�f�(o���g������_/r���k�;:n��-�g�۶5F(�F�[TÞ�&q�x��%:�K\�ϥ���D醏Mx�"��t
�ۻ8:����}}UR|�lc?ed��'�V�Fѿs��6:���Zu���v���RF��S�4%�**�HS��v��{ V��#����2i��K6xL��.UhD��$�G��G@:� �f��o��������7V�"�r{�i�3#OE&�jV;�pi�iM@�H6�:«.q�(J�[���ھ5��a��=�#]R��P8�.��CR��({�c��I`�ZUf'�ݤbG�{2a`��?e/�;�	�!H�
	���G�N��bS-oXw@���tdhHz�t���D�g�F$+wD�O���P!��/a������c\`�Q��qy�D��}Qԣk�[��L���`��ꍿ�e�������T���ckv�s󛂵�&��{��UT�x1��I�J�~�`�����K"c��_:Z�nS<�I<WWi
��V�t�*<B`�eE75<ʁeW��^�9��4Rc���!qtuZb�L�=�+�j��
�	��47)~��E��������.�t��7��Kd	��!�B?[ԓl�!²wqfP�F_��Ũ�.����$Dj���f��4^��{�gɢ��SMnAq�y��l��OhG���L�74�X���	�|�+�?*A�h=n�`���;���.4�4xB3<����u!�����`ú�3w/>���%2�RT������t��Qߵ��KY�Q�4%�`W�g�rΙ\VKb9@a�8�QB�}�M�AiXS���G��f)�o�����Y���r�Ch9�n|k��x �İ�ʵ�f�}�K����w�+��@iw:�h:���Hˤ�&�^�h~�<]��c���A��:R'=�\i�C���R4i\+{r�r��{t��rJ!�ރ������ya��4퀲=�&���f��	��R�Λ�#��~�H�	���H�^����߄����V��}���_���+~��XW0�=��G��,�
�\kV���.�TD���!�����䶼�Φ����)�!F���@4�3B�;z�h0���lxMb�x��:�0S��Ӿ~}Z���j��dx�(���
�� ����=���a�Zp��A�6����o������y�\��xH{��}�p�wNY|З1U0K^��$���1�M���n�?d�i�$����f:Z�L�~V݄�xU���ɬ&���%mu���@����<��<g��L�k����f����%����֌���Q�lt�|,�<|�p��qa�蝿r���tM� �ߊ�%D���y]��&�6��A��Ja��$.�uh�T�GR(m52�տ���f�!��2�%2>f@s���rvVf�l("Q�\��) ���
\�v=�.�aX;�����b���v>8�8�oٔt�)�]�;�N;�r���/V�ח���>���*P+7���sd��F� 7���^�� OE��_�<�"bk+�A��=`⹷Ԍ�U��@[m�pM�p~r|��xB݋U�r�(����0B�YO��Ё�]9�o[LHO��Nb��T��¿�u�y�Rs;	����^I�˾ѭ�Q�{tX�La�H��S�]b�T�g��K�\W�ŷXLN-c�05�C����p�J�ӳΥ�cr'��
0<�^�/���F��(������K�׀q*8��k�-*U���b��CK��� ����E"&����]���Y����2q��L
� �� ���(Xr�B� ��h��I��\�
X���ϯ���PX�o�m1-��O�'�1ԘDV-��L��@;�\�+M@�z-f=���օ5fr���>�6�m������pE����MI����_V���Wx�����%��RQQn���.�.��ݓ�-��8�q�t �9f���e?pC��ҧ\��[ڶf0E{�(uu0�N+�i����Lb��7�ґ�E��J�����0*���7@�z�I��^�lA'����"�r�
 ��,�gr�����8�Ӟb��:3.��7z�v�HʟZ���\y7�J7���uC�7� ����~B�2J�&��A��q��i :վ�&,��uZ�t C���S�_كm�I�c?�2�M�%��K�v�Tr�p)�N�-�iL�[�m�E��[��ν3��^��ƂlJ;�������j�0�^f�{�z�S������{���BP"�qCp��|Fװ���헻���M+/F� �ׄ�{���9"��cE�� �%[�V�.���/�����MFf-ݱC��V�m�~3w����j�����pu��gk�#�HS�y�f�����k�9�r��zH/[45Ji�&�5�
�7n���O�	5ȽA�޻�h�W˱FQl�v�p����{�7Z+5X�b?� ��w��J����U�gI���?�떍���t��Y�@Ɇ4�&�8�t��Ιߪ���h
�e��1O��
!N�"������5{0��1�J*���[�G'�1��2�Zf��I���Aڭ�K륱7v7*[Z��̞(��N9C�J�R��u����&+f�g�h����7*8�r���Z��>\Ǐ�����.M)�YHx��B��ua�@gn�^DZ[��fcK�YF� \��r�.�.��h�q�5)X>���k��Y���������f9��!q��Č���Cٵ8��U�_�#�q�u�K���vV�^ab��*	�=N�"Gd0W���:_)%N ?>c�؍���`����V�^�]�~'�H�!��BX���=�-���^�d���9�Nsr]�*Y�LZT�����wв�z����KK�d;E��U�c6�j��%eP}�*	c�6��/�ج~���������+e^��UN��bċ���(�$R��|���^V����E���:�ٞO��4��s�r9�@�q�ۨI�����Hd�z�=`��K}�ߣ�N �~=tֽ�z-:�_�7'�Xf�����$E��U�0;u,��`�Dv82"'��t�b�SG�]�>���c��D9��]��T+	c����q`��w���/ma��4s�a���n�;�)�*�)��~LS�+�+&Y�G��7��6����P6�m$�n-�v�!%�ȧ)}�/�;@��uE��X���Q1g7�Uu����^��-�v��f�7�@G�x5k��"Iވ�����t�`9`��<�p0��e�~������˖�	�����-��9^<�W������lJO���!`Q	��/O\%M� ����K��1u�I����Z˶���"��bCt��q��[aw�0�`�Q���}\�t��&@��'P#�D
4o�+uƬi%��6z�]�{'�����Ȭ_�8��i�R��n^b��2��etD�����}.T�E*J�`��K摘c�� 1��S� yΰ�b�n�m �լz��?���ZK��AsT�rf ��(�#�;ܮ@3�� 6>��h�������vy7�O�_B��6/�E����2W���2�O�+���U�OՒ�9�9C��Ɯ8��ŀ���Y�Ā\��Qa�<��/��ĬOz���j�GJ���8��Hy�Ʉd���� (-+%c�2��u�pML�;�:E���as��洣��կ`)(��w�E"sCn%CgPuE;~�+1�8�p�3?���`�b�_�g�?q�V��1%�m��o��q�;�aV����u4�;q�)��v�K�&��3�e�a��P��6mR�^3��J����r�FE;9���g�-P��A��{�aD� �L�=|��}���I��\b��i[��c�  f)���v��� O��7�^�q"V�to����Ǥ�C�L�¡쑒&��x܀[�<�&
!	LΟZ_c��B1���5V��.����W�4���¨x�ȼ"�J�)�9����=���@π�B5��߽���)�I��t��I�)Ab�ߡH�+�)�u�q�� ��$/2����4�2`b�3�m ����x��ٿ��mx�`�q�ӈ?�T��Jh5��r6�Ę%�8A�1O�`�>yD�!���
�� �,��ʸe#�.�<�(Q©?�S7y�*��0�Ҷ�#QN��+�;�@zt:��?�������IU*w��8B��$W��$u(VG�p�$4��:
q��c`9����N.T�j(L��� VdB	�T�)��ؒ�2��0�����L�&"2���w'R�������>qZ�L�,�T9�e$�bdaW�����K��+�K*Ա�І�%����xPK��݇{�r[q��x�#��\���D0�`*�2(5�!�m�J�Ny}"��:�,��~N(ܚ�1md5@�O�p|dH��]B\zÝ�����ϖhk4+�D^�����;*����u�k��d�����<��W��j+c7���p@�_�C"����Kj>�vdI�.�,T�􄓙�Gux��o�9��f�*��j���=��^� ���%Z�Ὁ���B��0jD�ݳNC��c貿o��A�P��B�>�i�8��5��|�[D=߰ ǭ�6��4� ���'^�
�5�-����ɔb�n����K^����s��$;��9��DF4+4<^D�(���Y��)�&>_Tv�S��?|'sa�(N��߰E�4�� ��vA_���~�1=i������_��n($# ��!45�t�@���D�Rz�<�n��"�)m#t����k]F�E�ZI��0
<QW��Xr���B� �@��e'��)�(�i�ŭ���l�P�Ĺ6�I����v�o߸������P���1�A�2����qj���}�̆'��^���
tk�Z�|{mpE�ݎ�޴wz#[��c�C؆�<���T��j���7��@a�~�[_Od]E��"�өr7	\Z8�Yz kxG��E��A�mt��M���,/h��Ig&x4cl�Am���G7��W�d;�C#��AI�,Њ��J�d�scy��4�G�Z�ceiZ�Օ:J�.�*���`Y<�fq e�+/�pm�cA $����6)���/e^T}Z�DJ�b%��h�Z�������m�VS�@���l�_#���Ab�>P;0m\M��)��Щ���j�y&v6:���C�~e@rگ��c�Enn(���Y2�CF�t|k�����k#:2A�|8O�wϬ�
�ȯ��ko�`�	���'�<�%c���1]SH�/ȮoEd�<�aY����c�V}�Ml���f����jG���$Z �$z�M�@@��K^K��9[���I�}���}NCL8�����~���>_� �δ2vg	�"�Jiz��м!l�t���ٙ$KH��D��9,i�oB�gßa~�X�=F��2m����wT�j��m��w:��s��WΣظ�]Y��ĝ���%Lz��t7`=��5�i�=���eC���<�pi�0\}L��y�%j� !ۺџ�̣e9�I���5�=��RЅ�16��@lØ�d�Y]�)���W�2�iL��p1\nK����w�����T�jA`(�AB%�x��'%%n��H!Y���jq�PW��>���O��:֯�)Eϵ �3�|8�p=�����}��U�_H��f2�4�GImt/\�>�6R�3C�ٻ"��?�M�YWeAR=4���6e��W�;���-�8��eM��c��Ҳi�7a8�����:�9��
Nf-�w�F��P�+"aH��Y�K���g�Gy��@!ڼn���*���Y.�ᾋp��1?Sc8����}[F��!^_�O꽲��78s{}�|���t�.�D�=ѓ=���M.���U�f���C�C8A�9Ӿi���3��Z R�����CT+�7է&�w�"�Ron�ο�Oq6r�����Ks���	R�SW��|�WǮK��B��fq�s��T^���P"�v/^/Z�/�]�z��n�^l3��:Iآ�5�T'��{��
͏15�{�������y��Ɨ\$)(���N�:��c2�]2h��8��Ϭ< �j����������V(�kq��6��^	��bx[w��G.���Y!���[�d��B9�6�aB���;>)����HZ�@�u��n������*xd_�Bf�Sk�;L�ҩ�k8�I'$ވ�?�����Π}@f�\��`;e�d	�����@�,���7]6�%;��(+GE��{2^�[x�o+3ѭ�LǶ�-�y���Ɏ`�#��?W��-e�ejQB-o�ݭQ��oJ��^�Y�y���!AiE9�K~f��k�r��l]ϛ���*C!����j@lӜ�	�E�h��J�EŁ�/��̈ﻦ�瀮�)g��"�`����rdVs��]z"����(�v��L��������j�����I���/)�SqsF�t�c��e�f������j�f;.��s]���:���LFi��b�~���������2Y���K5�Ta����Hwz*���s[�������t�G�m�^�Cr#&�PЙ!��YN}�-�h3�"\S�k�//|5*f_�L�	����ն�
V=Y5~]����(5�|Eb�����j�����A���`1�#nt�>���-�|��a���N�"{-��b�j�`m��"�%�#g�^h���ŝ=�C��k�
��ǈ��W�/�aǺK�*o;�^�ng%�}���w��h~z�+�"g��B�)6�&���9������!��X�W(���B\5�v�7��#բ`���=5�=��e���(o���d3l�2O`gJ�HS�C8�����$������9��'��A|,�����:Ap�?\�>YT����.�8IZ��b*5\����r�ΗW�VAw�����7���,)���K`ۅv9Ƿ ��'8�F"<	���|G����,���g����t���	UEOv,J=�^��U*���s�V��iF��*��<���ޱq����^��B�d�SN:p=���n�);a,Ug�D��~oֲ[*o�a8��r����[�r�ص@��&p"��#blRl)�?�ɰԴ1�������Y��B-�#.�],t���&?<��4$ہK�zieQ������mV�a���K>;g���ZG��1��u_�c��FH����&�PE���E^263 ��I�ZC|�?�R�S:n<=���!<�\�`�ȏF.A4%��l ;�QȤ��H+uAX�*wǬo�}Z-�r�0��s�3�p�4����������U��J�52�}?��#��Ӵ���L �x[�@#�ԝr�9��?�~�2��zym;��a�8��-I��%�c�TV��e�f��*J*2�)G�'��+��go0+���XQ$	�� �Üp7��9�D�C��Ԣ�$��iF��6Aʏ�P����s)�fYZN�."��������)"�f�wO]��2��+Nų�W%�����W�.n���m���v��EO����&B�.WJ��[���([
4����܇Y���d:�<X���U� ˁniu�ZĻk�Y�.�n50�\눲L|X�����O����2\0�a���Z���Wq;�Bˆ����˩߁r���nꦲ�m����T3�<<��{�`��D���	F*��^<�F��� ��C�z'��1_͙�v}����j㛬�ã��Es��8��㻋����`����p�Ң� S^���3���#��
:k�TrsV,%n`|d��j]����Ě|��2~���0��^	?y�:�o��e�K�TE�%��2�^��۔h�<{+��@g	a*Z϶�(J�Fo���W�h�k}:H^�W��2���S�&K��b���ϑQ�x5��K�p[��:(d��B��=��JO�וto���%0�Mᑉ�s������`�d�P��d�\� gU����.��:	+�����5KW�,���C��,�^윀wd0��P<ؠ}��>������Id��Y�.-*��{ ��K4�Լ������&d���Jډ���,TQ���O�������$aC�e����V �Nr���	�A	�D����OCU�<�~( ���o�b��M�Y☰����4��ѩo��&8x�h*��շc���z��JOK�[���'��?�n�:e���r��fI�QE����U�*%�K�YB�L�Y�^����m,��*�����m�Va��v��t1PL�%�jM��V*��l&�?F�T�Q�V]U7X1+%H����FMfeX'�b����	�	/*����?� ��9��[A��,ԏ�G�n;�i�݈�~C$�	��Zp�z�����6��/5�@�{���0��U󖗫ƾu�� LA��W
��P؆��Tasr+��/6�e���ίMe����Á��c�64��ה-3�[��=��h"�歂�]K�W�		'd���[1��O�LC�<����j�j� U�b΀w#"����u��U�Ǹ�� ��~�����!DK�'/-�TY����]dkN�Bp��Ŀ3oͶ���C����;�(^1(@[��6����H.ęY.R��|0�/��E�0c�����"�$�8���D��c���\��2�������9��wa��OJ6�lS^N+Pܚ�c�a&�a��k��b/J�����[�\�o���I��
��&������SV������"!cHh*��,vi�}Zi�h�B���r�j��7�X�x0$F��8(<�7��h��RԈ�W��#e>#^k��>S"ً\��Wv��28�l�T�%��4?Ϭ|Y����_St̊���X'�(���8�B#z����w!��p�bK���$�~M���~JEyU�a�����}�݀rOД3q�U~d���JZs#_E���'~9Y�J��9g E�^�[���f0h:��oBP�9���(t<��O��"ʺq���V]��`H�����ÏU�㲻�8>�;˦�ibTϵ�ԛ�i(�F���K�f��1ǝ��al^hC2�3/�A�.>ДH�W����Q��65�TZ�M�r��()�LS�� E�Ϧ��gU��R�EPk�w���VUC@M'?���a0_a���²�Z��,^��-�����Ԩ�@isn$��OG0Lz�r�L��盉y�
�G��O�'H�rRWS������X����y/d�\9i�A�Q�W�X�tZ�֐jϔ�N�Xm|*8�Oz�y?UP�+ڜ*YN�qt����˲Y��J�f]���H��@=W�[Ć�|E�E����y��j줰�edW$�[����S�rr{x�y�{���N�I~��P�KO�;�Nu�7���7�G����,*
>;�ݎ��5Z.�v���e�5���*_8�P�-�Ⱥ��	v����N��Z��U��SOV}�)�T��D^�7���,ݏ5q���n���H,�+)�?�ؑ�b�m\��GjW�Fw�	�,#���~������ziN
��t��0��(8̐l�ƈkz�C��E mM*/�jփ5����&�o� ���h�f���p��8d������nV�b��x�;#��*�������ˀ�1����WIn3�*%-ڰ���|�m�9bl?m��v��qW�������6�)�YC�nT�ޯAb��mCڜ���-�?ܿa����v+X�����C��۟m��8���i�i%a�!Y�_�z!�$'�Ns�X�	�05pK�GA�&��y�m���Mj�*�K������mGf���:e����ɧ�3���q�n�\�m177e(痕G%_%
�{��`Ƴl�^|�ց���V{P��C��W���xvp H�� >?c�3��Tۨ.��#��-ح�KO�E3�0�8�P5�v�1(�eow�T�RE�/�A>���Ǿ
���9̽"���q$v���A���D~x��:��Ð^W<�G?ӛ�ӿ��,�ܹ�&6U�Y)U�w`���N�ѳ*�?����֘H��g���G��L�9�[�/�8;����&�.�g�n���]9k�D�%#~k�>2v�����|
m�H!rd���:^7����BH	�UL	7�Z�Ȯ����Vj7���=� ���|���G�l�B�Y��]��+`iT���c��_�V������m�<z4�^AS
�^���^&Tګ�\K�ɀA���t�t9-?·��G�h�$��_Җ�J�%1X�vn��wN�a|�x�do=���v^~��/������\|u��(��H��MN��1�b}���#
���4h9E@�h֬#ϯ��ް�UH�H�y�z������:��R
��fzn���w*+�twowy�!��Dp�׮�O'�a�6H
���[���t��������P����zn�o�^BRp['J0F��*��N-X�����*y�e4�M�!�G�����Y�Vw\R�R�IvY���NF��`�O������Ics5�F����|��$5bX������������cS��s�D�H�����k�1V�!�Z|�R7�>CÖ uޕ�$��
( @m�'V�(��i�1�Y���[8s��N/C{�h�\�2�2���EK�I�#����A���JU���
�D�Ys��qA�:BH��&���Z�YN�N	9���m����E��*:��͌#��?#����/]`��{��ޖ����ރ��d��&�I5�+��2�G8�}��x���!8��QQ�<v�^y�Q^���ʥ�;�bg蜅ǁ���7�&њi�!�}�uߍ�}ͻ�@{�W���!�ef<"�'\�q]c��q��Xy�H�M�ǂN��a`�����rnٺ��~��)��Tw��n��lva+���ϖɪ�c��YG��-���k�,OL@d�^�\e�1AC�F"���Dv�����t��F�:W��0�(��e9�?�,�	���P��\��=��\us�U��&r�'�I�%���xgf(J#��L��@*mӽ�瀤��Ќ#o���)%A�1��D,���Q×U�Ҍ�I�0]W^�"�w��L�3��ɶ�t{lYHf��ң�����q�T��M�`v���x�U�Q�.)�v:H�+����0��\����_'��\�&�]�
����k��c8���$�@�%Z@��"]�orh�Ơ@�e?��q�1�W*OC�|������3�<�Jے�隈.�U5*/�\��>�t�̪��\�@mbI�H���Nm���x��oKX�i�+O*R�G���W�Y-��ĩ$�2�`�!x������H�2RX}䐻��.���m�	�9��s������΃�1�`,�׽hl���l�u�aJa(����8�_'���-�#Z�[�eb�N*�I��4^�pҶU�����Kg�����ۻZ������O����a$��k[y�v�3O��a����&�ϫ��ڑ֘���Hh�L��.c��Ś�x�����V3\_Ჯ�N]W�u������g�Uo`��XL���#>v]U�$ނ�O�Y�rVd�8�>C��m�ͼw@�[�=G)pӝ�<Y�;W��u�x�M�8�$.���.0���3�[�_�����Z9{ #��:����;(��l���z���m*��XP'�(�SOV�:r6�jW8-���Y#1rl�����9ꭑ-�R���v��!���nt����)�#q1�Z;Ç��6�TZ��.���D�����w6zZ����î)��P���B�x�=�������2'*yWU�~�|��t�ŀ���h�L/�Ж��'�����>y��<&adW�1����S#ꗲHAKc����z���	]�
�M���Z����U�x����p�p���{|�@�?gi����Z�B���0e2bLKP���x:l�p�:;��)%�8Y��ꤳǹR���?=�u��9q辕�m��K�I�`P�PS�;���H�u���9P��2,Ve<��.�x�U�N���:�h{����4r������F�c��U��jEwe^��A&<�R���?Ky/�]��Z�3I���;����&��έ<���{@��{D3&�Oa�n��&:�p�w�[=�@+�������h3����l�7O%3w"`���3e�i���l��SP�4�'�`��f9�@��^qU�1�P�/[�%�Ͼ�S�`	)�R�.�4��W�.�D��NA�*x�¯�=�Ox�q�����;NY޹ќ�ޕ�R� ��T����(w�XdvbvFg@�<� XN��<��7��rm`=^�z�U@�/_�����Xfb�6��~Y�)�dg�JXq�l=�F���Pr*�f��(3�ם��FGdEr��8l�n�k.o��EoO[���#s�\�!��,��͇�e)l<��\���3��:aG��o���m}Ľ�7}�p�Ϫ�{R�^�0ܪ"3؞�Bp�yI� �b{����X���$.���^����$���\X�[0�<0'��_ReZ��Sz0�
��~�	��?S3~�ީ
�iϟ����]�i�����b����g��1�ʄ%%L̍Q.�	h�>��;B�B9�$�eߙ�K8��J6�y�g��9�g=��,�`�J���D9jK1�}������&����9�&����g��D<14�X�0�	��=ۭ��w8��4�PG;��Y���E;�q��46�Х�ѕ������+6�˗�.�����B�B�D�����V��{IM�7	6�OQ����KJ���S���*%�.V����[>��=a�F�g���V�W+�|]�K�f��e��2�챬��-$2�bn&�q��l�;�6�ǭ�X�ܟ6�%)ƽ)V7^Q���#:��OΎ��[Tc
�*K`U��GTcl��Yf�%�_����a�R�\�0rA3��I~ٲ鶏f��S��]�	"��9d� �\1�Kg1�Y��RD �OR�%9�L��`H�;_oL�k��5��C��9��*�
�����r��ǌ��FR"��{'{��%ǩ3+�<#Z�Q���(�Cն ��{������z�7�q�1���݋�(� �~�86���iz�p�]QZ��p�4Y�p�	�@:��<��lJ��j%��oJ~j�ˏ�>�=��*u��"uGK�!K7�y�E�,l��Y���Fu� �%iv.x}�P��0��ݽ�TK;�u		��2(����s]S��:�)b�cŏX����S�s���%eV�!Ů�������jG��r����t��H��Ӯ�*��JZ ��%_v\���ҵ�l�@u�%�>E3����xt�nsr�l�۽�RT�v�+��>����b����R���M�������5�{Il�R��U�:�+Cͧ�f�Ik��yT|㙸�7ɝ*Ⓞ���%�'��:�A�uԗ�)��<Z���P������#���6�ǭ�jқ��VO-6�*:�|S�k$��h�������n��D���w�	˘����yi�2������h5����k�b�,W�IH'x&J+�7�l�,e�4�{��̩��� ք ���d1et4�ݽǆ'�\8T�Zڿ`�R���6o|������r.A�S߇h>`i�ѐa&�����i+�E*���
���'�Nݢ���V�������៯/���
Xo�}.<�U�#���i�a�b�?��6�����>�A��Pc��1i����;]��;�0�~��K+?�ڨ�3#�s(�󒿃0�1O���e�s��@Y$(�3o�^�0b"�؝�.]{���/Uy���Ց���6LƤ���d|�ҽ+�)T3��r�\;�\�YcY�E��#�zJ<����bvь�A�;�Dg�?v�By�R��FO_r�.JJiF���y�7���[��8�{��G7�4�X{Aћ���,���mѼ�s�d
�$��#���+�.�5'c�)�c��G���n8oBǷdm�����|���V�H�,�F�u�[Z�Kb��e%�A0a�8C����)�K����u8+�3nw�{m@oZjd�ϊ_]-�g�7r�y�^�(��$ ��%��^ޝ�����Vȑ7)J��P���Xgg�n�f�4|>����U�]������a8����Q�2߃S��8���f_*3� ![i�e
A��+�JBP�L���B$%l�^/-M���~r_e,;K�����Y�
 T~��
Y"� �Wyϝ
��F��h��3k�� Q����p�,��k�j�7*ޭ2��ڟ+�قFD2��~3�JR�C��o`@��9Egj�G��N^��70�(8-�O�U�Xr4do��Q���&⬞����4y�>+��;	u��\��ހ��q��t�Y"o2B�����[]�t�PD,�Eۼl����<�͋��s,��D�W?�	��>�i�QZ¯c�	C�I7�F���`Ճ}����6���"�P�`ŅU��l,�"�|12%2��e�"|]u�q��js����\�f@�1��x��?x0�m�*3���rleo�Pf$\����O���dx�,?�{6L�P�����Ȋ��rt�؀�1F�ھ��f 2W3�d��Ḱb��@�h�;a��=����uW���L�'�}2���lT��P�崰�.��ɥ��Hn�j�3��g���}%M),N�\�p�d�b����7$?�]%�~�^�`���Dc2���D��kJ�$-�0���O����p��!�Ò]_�b�W���M�Y�UQZ��Ҋ��K�n�+P~]��a=!�	�r��dE����g:�����՝؜�]L�K�ܘ$��H��[W��~H��`��P�#��b���O�̜�ۣn���-%�w��^�����	f�N{xM�j�C�~�،GB͔|#������K�]�6��u�Ʒ ��D�#�|2���}����+*�q�S�g>�ؕ��q�h�5���cQ%"��뾇����TD�S�V�~(o��:(�-�g7��.�\��#�w61γ��THW2&U��Y
�U� ��N���n<4.Ĵn�>4�K��3qw/�e���'%����Ay*b�.Z0��N�(#!p�5'���z������� ���m�b�+3�̦)I?�R���q	3>�.�V
HKal٠@��>��3���E���/^j�]^v'۬WP�%�&lS$��G����R���_*�`���)�d%1�N�����^M�y"p�Hi	O@��b���9r��zu �y1������+蒁���V/% ��>�/_+.����uq�g�9[-:L%2�u��D���hMXv������*@��UL�S5U�q-���/qW�[���)�-a�׍�_b3����Św�+�@�X!4�{m�$cr}[��B_D��3�"L5+�R�?�4s��-�Gu���~|���v�B:>56��c������n�k�f����1��؍��d�r)�!r\�.IV�z�I�GG>TW"��:���2XWe;�l� ~|+�}W+(ĎJ���Wx�^�a7�������E@�V�;�ж�Don�b�8��}ZqAU*�hS�ϱyz��_��.�s�"<��b��>�p�����>���
�<!����1d�j���w�X�0�c�A5��c�x��(�����?���&2Q�Q��0�-���,�:�ݡ�j�mI����',����ۜ�a��l ,D�P����_���f*h�h:��1�KI7«u\~��Hi-ZX���S誄>�����ֺx���?��,��=���'GSL�b�� ��y�a�k�n�FW!��3�c�a���r�fR�<5���<�nY�z.3��f�
1"T���W�B���q���6����u�{��S��0�V >j#��? ���K�A�i)��*�5�(�7��u��Ԋ�s��'��]�_J"d>�R i״<wO3k�Lm������?ʹ�Y�b�ђx���uպ)z�ъ��p�p�#���'P�-��x���H	p4�����_���<��r�9[��x��ui��@�����p�Y��Ւ/{��=U�d]+����	�@b*!���q��w6@��'�^�c��2%���
%������$������� �v�D�G%ʸE�	]���`Fl���)�w`!H�d���n+�b?K�c�l�u7@]N8���=7�\ڕ�T��k�7�g��9�M�Jl����d�	����Q�-���4�� ڂ: �Lf8K��&^4���.� ��&7�_��]f4�D���$�*��V_�0�4%{D7�k3�wC?,n�N���2�����/��6�D�}�*��;�')Ūr#�7�H�&�5�˾�o��X}��x��dI(=�����/D�2�����*�9�,|�@�ԛ��1�����
y��ZK����dw88�;T��rYoeR�8���H��DY�K��KS�>I����L@�a�`Ec'����0���oF��h�oM00U�N�[r�zL?���Ei��{�ô"��$u�ah�r�q�s�� 7n��"%��l�����o�J[w�m?NF�=�h�4u���My1/� y��N~�.L;��Q�W��ı���Мo	�r����"�1Ӝ����м�n��)9˧N'_�>06/5�q@�عE��h:�A5(G_��8߽�G�2=��â	�!�)���׌��hB��6R�B.�%9�%B؅��X�H�k�E�t�]䑦PD$
�T����֒�O���p��\�#lS�����M��y��b����?�Q7%��ʜe��⛹xAd�6�TbT�b�e��3/�K�e�}�T�������kf�d`��вl���B���Um�w���u���֛�,d*��t��J��؅E/�A�� Q����f����p��-���}Z��l����:	�C��lFx�"��K/��?�K�`i %�֮��U����-VAW��^���-�{b�������M�i�����͜�ŕG�Ma]>��)To=��@��D��턈<RF�����.��ڟ9RMQӰ �2z0S��w(�.�
q��`}�`��EV�] ����Y&�_��0�v��,�v�_���`�����	�Ɯ
��b0�����0G+|0T2D�<VU?�FT�q�~l[�[8=J�)���3Z�!�>�'ku��^.�}�i�;ZHE�l�D^�dk�����qy�����ʐz��L��� �V���}��o��ż�$�A��?J�S�U<l�j����C���
�5!ʧ�!hPU���,?�#j�?�9{~�\�޻8h����cW~����Ж��>��i� �	>61������
��ih�G��^��3԰���
��[�{�ι^xX���C_��	���A�~��B(��N�'��U�Ԟ��
5��
��fL�֜��@SY.�&L�k�μ�Q��N�Ł�?ƨj��f~1Mo=y�<ܶZ�sd+&6C��E&�ˠ0/b%�n6$��E��B����Ē:�ݴ}�WQ?�y-lM��,���oi�9ZZA� ��W������\���@\Ia�N���Dր�����A�q�W�U�����->ب��-�t\n4p�N[��zc��S�����SO0��u�p;�T�s��u!�vvĵ���Hi*��a��~t�Q�󮂞?f歽 �ŋY�g����ڪ�\�J�ۤ��X�w ���r�e�G�Rm�ZZ��J�S��G+bi��p����+LZ�5t82S�{d�o�W�ys8���$��uk�,�
���c�����>�o�bN������<��[AV�d���艤�tF�b��BC8aAh*�+��oqC���jR0�Etٺ��ܜG��v���inVI��g�)���t����ɖ����Ec�62��:Dj��p�M@�u�J�D���-!��K���ƻ[���:ۃi��:@c�[��Ї@����bñL��s)�	Hv�aN��f�e�K|Mެ�	���ߩ�'zK��g��O,2�E?<��p�R�}��t��N:l�Tn�Y�=B44u�3���'u��lV�S��&�k]��q��]�ț��m����(s'�^�+������&�d����f0����a7=!4~�c��q�jz�A
'{L�Ѯ��r�)Z��!+vKP����������VoI�y��^<n~̲���ޡj�{�j�艛���w�QM�'�bj��]0����Y ᷌�;��K����	�&����:H�Z�F�Ҙ;@v[�c�S|�N��漧�q2x�変o�ć='�3ƱY������%�x,PΔ)˽�vH"�iX<M�Z�M��\��~q8��K��0M
�cK5�R<(=Wc�P+h�� XxfL��$n	&���N�h�\$��j�A��0�j�ĳz�#D��D�; �-��υ�*��`��A*0�$����,��fT�5��|��t�; ����*;�SuMF�j�4g;ʖ:�"��T'1�+�Y��|Z�U[6 ��"x���vH�bX�
����Yk�Or����XJ0|L������W���l^�f��v���ޝ0�l��ZHb$�Z'��ZPb�PG�����K�5M �>����b�)��!�l����leV���h������5�kY��b�\]bm?n&�њ���� ��W���қ�둉i녩m�
�W�T�,/���uV�%�&�J����ĺ_�	E
�E/��u&�'���S����%p��ʇ�l(���ـ,g[�2��K��j)�qy�1���H��= �R�0D�g&}�� z 裊�&f��D��!s�@\����J�c���nk[��az��9T�!���}������(8&�b�	��<�������s��x!��u�
�K/̿}..Od�T�GT�|Gy�Kl�~P4�\'�.%-P�r���N<R�(�<�h�)���� 强E+����L[��M.������3p$��v����q�]p���,���|��W�ddl��k�g:�9��P�f�27�Z2_�	Gxw����*?W�Pϩ��j�4�ZJ�H���6DK�Cw�A�e����	��mY#��N��RD_cU�Lb�4����/�p�<��-�v-:t�X�"��Ț�h���D�n��c�6��N������6XR[0*;�D��� ��Iw2����xm�V<
��3�B��؛�����4d�%�B�˖Bs8�\�����tw@�^g�[�vP|*#��C@�g�����"0;�:�a��o�>�-��L��1#�jH����ˑ���>��^�9�~&�kY��#�r�7�~)����v��׆����0Ǝ���>b�9L����B$ƍj�^#�֢x�UM��m�J%.����pa�����jj�N����D��1�Eϖ�Bg6���[Gd $�V�)�JFT��|7�*Z\�������ϱi�� �Y��gy�U�"�.�{i�u����7+��g�[C�9[��w��ˊ4��%���e�	�Gn���o����
dF��(�<��Ր�m-&�8�#�;��jkb�A�o�DH�ӂ��yn��ekZ�#�r�������9Au/t���TP��K�CF�ԇ<j�z~t�ow�]�uX���%��ߝ�)bU��C���(;�o��c�=2��8�����7 9�� U��M����_*=�fL�e��Y+�k�ozbR'Hwr�����
}3��L��jV�oQ��V?��84��X�͔]�h1d5�)��n�"wB�0�,Rw�Ϊ�����" �N!�W�� �f�0���)m��nf��/�˧	`<țU�F�0�����6��� �lטãG���sy��Ȓ|�=��������)��
���n�Q�-I�}�!���<����c�c\dT�#�ns�S:��<�W��铭�7�c����)��~�:�NC_Gҗ�|�/-�p�?Hi��ǣ���}�*�bB}�蔡��9d�|�n�fdU��}ڝLd5_ʃ��`
c��Y�$�-�ԉ
i�7�i=o��6���"�'�i7��=� $+����%�1��m�^�(�V/p�R�'�9�=Q����ˀwzK��o?��K7p(�D��\�ȱ9&p��M������H��*;K��U�U]b��Ps��+��,�'�]t�5���@2�j3<��'���i
�"L��3���JN���M�9�=���c����
\�Mua���T���Gȣ�� �5c�.���6 َ���i�pbz�)E2�a��AD,[�֬ž�lؙE�U��(��6��1v�EB	�%�4���hڸ;��½9�,*��<�����"wڥ	�s�VϜ���NJ���HE��C�cho,�)pl�v��bݛ�4A%�TԚ<m��|\߮�b��awg_� � �bI|[�|��=~��#ԅ[ƿ18@����q��e)Y�c{q�}�mR�+��q��Q�;H`NC�+(���@ �	@A)R� 9��(j}��>��J+1�i��Vr���)�^~�}_�g����@ѝ͚��J�y������:�#����K(e�u�����J�����,)uM�\U{"��L��2��DK��ťX�2��M�O`��K l��N��EU>�-��Ss0;�D�C���U#s
��P�pC��3���@I�S���`�k���Q}��+0<s��Ư���k�*����G�fV�ܧ�vO:u�@?���Q�+�
@_��#�X\�w��HZLh�	
�JLc�^wh�����S�^��p݇X�#�opv��17�x���Dd9�) ��J�ʝӓ���ar�6����{�d��_/�VW��!o)����:�LϚ��"��Q��KH�Al�������<�#	i�����/Yȉ�b4����H,�u�l:Nr�n�z��GX��P)�k��щ�� W�K�5.�+��P��RG�{!A�6FL�<�e���\g���������Šx�l�ۮ���isV��Y�Z�|��1ū+[��f��"Y��R2�����L9�I_��K��@�	=�y�\W��h�^Ά<�.)3���֒�ET��g�=�V%��F�i㥨3����i�h�j��r��q�n�O~^t��	4t�]��瞸�x<U��|ģ�#�;W�!6 �#���;��i��Q�𒾠���P%:mt;��Z�[�qM6q�$H��fP2-$�����&���,�Qb8�:�޷$Ug��6q+Y����u��Z�*�8�|xo�1�����7�X��!�s���5��m�ڝf��?�x֎��޻1ב������)F]�F��V�wc'Ȗ�+��-c�_���$nCkH!�:Axɤ�mC閝<؇���������:(�̚=fO]Kg��W0�S�,�dc�m��������|eD#���=�ɇ]u���N��*6��݉ ׂ��+dy���d2�h�V�+�}Öy �p��V򍊚
���Зh�]K��u�����԰&ɳ�A{��!z�?��:=;}��Ҙ�h�^��o�s"[�ħ�[ͨ�Kk�J-6 ,��8�ZB�x*N^����5M_8��N�<�� =~H@�%�p�f��䰯/�FW�#]��k�M��Y�C=.���q�x
�m���2�s���O� 	��$�1�A;x�
Y��El�(+z��'`c,>����J1�f���G����M͙��T��UqߢT��Ox��n��SY������m�E�S�∍ǒC�-n`��1k�[Y�#�|�f{L�!�7�4���0�C�P((@�5y� �{���Ed���x��O�#^@)xb�B�����(��a�~�c7ܭo�4�,)�����	�5gI�����b8*�	�%�ȱ���v�Ԉ�5��01���)j�Z �C��4���%}�M�x�_�]����J���׉~wR��m��ý����L�"���D_� ]�c�د)7E��),Tض���ϊql#�jT�Ǿ����3�`���1d���٠�09$%�V����e��YZDN<�(�ʕ��ƲV��b�B��$� ����K��n\��g��D_��a����:MN0'^��rع�^�� wr_��� ����Fw��髒C!]}R�}���B������÷��G�R�p.l]�̪�?O���t�޽h'���R!�`�h.'@��x�Lv\�F[�͆���Au�1^T�}��6�b�+���4CUZRQ�`�߹�Si��2J('D�tJ����؊��_fXPS��e}�vF�`ԩtl+K_G��Y�տĀ��t��1~���:Its��TQw�H��W�z�&BX@���0'�彖�r���<�u�����W�KXU�������B|ݎh�,�p�4zn�������ʨ^CW�Yzx/QZ���C�j�����?��r�־n�
�:)s�Dz�sMǲ�K-BF���V������LJ8�4�r���CWM�=u��3�'���g��r?�*9���!&�)�9��4�=��b��y7�ۓY
�;`qfi֊��S��g]yq��X:�[���b�럤�F��u�!��jf�0�@����$jt�Bw��k_�Y!�~�f�=����k�fiIcn������h�R���0�* �6�o�jy���Ҙ��4`_�����Z�
��/x��bRƙ���Ex-����Q �z�N�i�;{L�Э�=:�eðk��C���q�E.}�,�h#�/�����:��`�/Oe���Q��wI���^<�#����v"��7-���}�_]Ǖ��8f�yLC7
��ye����͑$�^�Ri�+W� �#����b�]�*h:���'��HB@|`(�SB�����`��b�s�ϝ
���@�H�����Y�i�9�qG��=�����e,�0O0� R�����㖷�
�D&V�OT�OC��Ybƕ�P2��=B������%��S!� ˘f����T�~���L3�9t7��L��dz��� ��6�����u�1TV�Z�X}��\���੓�0��r
�V;�|�`�z�~h\.d^�R�5�bWk����!?�cu9WZ7_�J���g�ÐtH��p#-z&��QY� S���HAۏ,m	��!��f��£+��%0�-�z�a����9�'zB�&B�7�����������a{Ե2@���6i��c��܂\��#�e{�HT���x��SL�^n���Z�7�R 5Ñ�:�������Y-��łR���e�YQm+f�����D�b[�ݧ�/�$n"h=t(o���?�΅q~]ߏ�W��8��QH����W�����ǹM��e�����{�"��j�F�\&�q���ˀ�V�[��d�hr�!��=��S���x��"?Ξ���s3��������|�8�w�l[ǐ��0�PI2�>�oLdVz>��_������Ó4NX�os#�׼	;�z7b�|�FU���5���5����7X8��xo�U)5I''���#��1���,m�L�l�}�N�	i@�@��r��?5[c۱Q8Zoh���� ���σDc�O��9E��rYD<=B������ւ�3�k/7�&�}�{6�Gj�YaS�˒��y�����̞r�EqJ��/"����Y������wϻ�Rk�l��i᮷���$
J��07�J�\��z"'��yU��iU��r�I��S���5B<�[�Y4�+�i�ԙ� .����pt���k5�����:T/��nY��;i�
O���6
�+X��#1�q�#Ѕ�[qgWEN�M��붺S#��j�i�L�rEg�$�X]D�_��c��\��n��#�J��B�\����U�������!:އ������bQ���r�85��@%6A���j�C��.녢�fl�t�k���v��=%�>����Uܠ԰���Ǿ�ީ��tH7Hpku�e���%�-�[��!���Wl�B6o��,��ᰂ���R �h�dT�Km��R/}"�a�E�;x�r��R��6�{�_j��뼲P�􅁏4 �^~�!'7��A�����Fttw66�-�,I{8��{�q��܊�m���β��	�c]mұo���R�	z�Θ/"�H�r���D��u���4>'Qw2�[NΣ��Q��+ɾ����|���L���ĝ�Q�8��h���]���U�d��=<��C7 ~�޼�ޖSͫ|0<Hlص�@�0��1u0�<Ait?Cx��O���pX%���7�p����o��Achp _�m*�2�"$���A��L�!�� �4�iLO�B���بo3�	�f΍_5*&>�����ʹ��cCi{�k@iZ~�@�7`�]|�v�=�9H̫g׹�-�=���h��^��w��V�/��+�u��j�
3���
8QW�-�̶�@X{Β;nq֢9��>�����{;d�A�NFɆ��'�ƨ1K���|�b� ���:���O�Mj$�d�ij$݂�F�q�<�!;;�g��9F{�u��@�� RA'���� ���w$`hq����I�>�t��h}B�S�����o�PLú`J��>��\���5��C� X�f�O��p�R6���rɢWUn*��'�p���H�"T���J�h~�љVMK�@�J�����Q�&��ç����Ii�Sin��ν�g&j�C�(Z--�����cP-�ƙ����p�wI���i�H��Ê����b�)jH�F��k�y	��l�@`��	����^���#���A�^Ⱦ��uEH��[�#�^1�s�Y��_��nQ��[�D1v�ۈ��ŉoH0D�PZ�a�G���Ko��b��Ub�P�������0���,C.�
�[�s�}�U�7�����x��q[t�z�A�a�8�KM�LL^`�bs���CFNi#�'� �
	�AtE��;�$�Je&?��IzV��LL�E+��]��^dK��.~8s �-�&++U̇��@w�ŋ�u9���;��G3�Aΰc�Ě�i�]��.��O��K4�V%������`�A'FV"��T"a�!��4�?��C�F4w:UPS���������:��&�!��Z�T0u�A�4���GDwP�|!?<o��B&����-�$-��e�s0\tw"���hse6�2:�\��."4XS���˒�}gK���8\�#��uv�-��+�b	���A�G��1G������&��{_�w��&%����k��-S����@��q�fR`� �m4��T$���`�T�r�%A=�x��vs8�4Whnlr��v
KT��(�2����]nղ�21Rڣc>��yj�l��t�"�nC +EQ�OA�1Jw��9�*�[�A�� �8�2�B}X�����K�^�G,��	j��+�4V��s���E�k]l�u!�X�>�[�(�[P���O>�҃����֗���2���)�Y�9J�u�}��{�#`ω�)pY��k���p���=Ec�Uvժ_��c�d��z��٧�h8�F6 L%kg	���D��Ԋ$�����.J�ō*�5�2ΧFb��r.|�+�#9Cl�"ֈN�tgO:���b��(�y�Z˨aN�<%B�xWC�NJ^�,�1��޵��l�:�|�� 2�טD���))�m]��F�'�O�:8�g�'����b�P�c}��%Y����P��9L�2������������S���Qe����s�f�����0Ě�eH�Z��F�>L���a�
æ���C��g���A���V�oXE�)��U���z���1o��e
ߚBo-Rܼ�ZQ�C?�����C_٨��NNSr�j�h��ߤ�X�x������$F�s>���",މ`M��ӿ����G��n$�j������sa�D�E�f:�q�iؑ�wӯd3
}��X���X�-5��, !�>36���Vg�X{]��񼦲U�%����3����"�N$�b�p�����;=%�7-�\�UsnL��u�W��\)G�ҫ���#T,m�V�5�m%�g0�]��F��#O�@��_�T��~��g�`���p�u�s�5�oP��Mi��Z�^|��sX�e�~�l.2{�T������!8�@ W��AXֺ�*�o둝a�eRP����!ۼR���k���=�'��R6�(���Ψ����G��{;IzQ,���I��J�L^� ����Mw�W��$p�F�$� �ی̃�f�F�%ŋ#Z��{��\�]B�Rf�/�7����-O|"g�4�K�D���Eӊ[ �Ql�G��F<���3�I-�%q��g���Y��2�����]��UC�F�wN���^śE��{�(�BDDI�^䳥� 6�GCTE�-&잚�卻��p\3%8ҽ;��o��L
	|�p��<��]��=_�%�:�;�2&:a�v��������Yt��JN9Wo�pFҀS�s���Ln�Z۽�ѵ�{�XC�Ǝ7��'o���O'� 0����{5db�W0����3@�N��"�[J�l%�v�ܗ2ثZVT���(sƴp�OK�
�M#��D"/�Y.�y�W)i�i08�#�����/ck���a���B�z��3M��؈D�"��Gv���⻹����J~��2d�d�W�P��-i�J�6tz�x�C�ܻ�@�#h߽��Z�~�[�lC�&�4��e�`�������=E<$�FMS��1,$����.�&��ɶ����LkA�p�[��;��CJu~>	j�G�'�f��fȴs��*�Ah3��lsiS����?2w�0�<-�O�_���!��?���
q��\����"�8�]a���G��wگ8��f���v�N��[����}�6r`b���TɅVS/©���#�L�� �����!Z���$��"L�^E�bA[��,x9�v�����co�zq~���\Pw��2�6��dڳ�bC��4����[5��_g���]i�mz�a��g�2C�wY�}ڽ)��:�S�E��d�?o9=����jh�0��	F��ݱ��$q�j�7wR����T��'���8zE8,��3¨/��҂C����2^%;ZOڦ/���-vԎ$	j�yT_��U��0��of�00��y����pپ�(.~�㤓�,|����d�x�a�m�85ag���1!�C�p:M,�xsS�0��q�����>�Q��*��V��0TJ����OSs��� ��r�N���T�:<O��9W2J���,g�
vJ�d��	7 G]����O1��T�>�SA������K����x�N�4�d�MX�;JuP�9N��`{K� �		���� ��^I+vό�=s�ֱ�߬+�E��k�گ鬚��K��K,3H.9b
�S	)��
x.Z"7Ԁ#YI�z���Jab$�b�	�N��oK�د4�煐�n�dVb����W�5���FZ�r�d���Ű��<����6ޥ���Ixs��l-�-�z��Rj�����#�΋J��������;���)ZW�|��@�f��v��W�"�_�����j��0��)�u\�.���a����įϕ��<�HUK.x�0���cZ�{�7��߹�+�����jD�w"7�|��TJ�����P*�`sqV%�e����M�I!c�~�1��@WY|ْ,#DX�#&������n&���X
�M(s�A��@�Y���%��s��[̋ɡo���j�C�ɩ�J����۾��~���^ahL{I}����k�Y�f����m�33�S��Y��4��+��f�g0ㄱ���t4ֹ���%�k���[���V�WT.
o�Ǵdqױ��+Q�kQNo��p��sȣ��7q���"k|��J���r��̪z"}�e�=h&���7�L;�4A���Y����ً%UB��U�C���h���AO�}a��l�i|rJow�4�38�(^��Py��Z(d�D47� �A� �^�����Y�v�\��&�%����^'T�������F��e�����#�Č����
t+���h'�O�!9�ǰ��Ք�*	G��N�c�`_Q��o�1����z�(.ܗ��CT�OfZ� �p�����*˭]ڎ>�����+�wx��+��/SDD�D_�+5S�j`+��mϢ�%��$�v���=u�� �t�)�J�&ș�8l_��j�l�5�T./��8�۔����۵��[��*;��#���éb�}D���6��f5vv�>6��K��0}�����SYw�K�oA<���%Rn�o|s��
a�����`d����a�?l%KzY�T1�h}/+�ӥ1�~�a��w�)�����}��R��v=���	p��6�����=��?�?S`�/耔�7�Z��@ø�{�+�Ы?Z�P���`�M��k:R��{� y��u��6oA6@Ķ�.�$���(��]��1n`�Dk�c�(���m��+�y���-�ٺ���
X�>t����9�.����$�7�:jR��T��<��0œ���TJI���+�e7���;��Yg���`�`��#���3.����7�r�~}˂���K�tO�[@�`"���qǗI���Z���<kdY���]��	U`bP���V�z��/���ѥ����9�t��,# ��ca�L*�?˞[>��ftׯK�%�l�Hb����'���g!lŅ�Ǭ?`�{B�n|��2�@^�Ԓ
G��'�K�D���-�kpZQ�2�^�]F��QUy>�A�h��l�n쏊�6�e����X�?O�UdG8�SO}ew[�%�"�����AuM:g 	�����%J�h����v�jlCk��y>�~�S�;ѣ���������X	������	�ů2���5�����"�Տm�An���	��P��?+���xdB�aZ�T���B�"�R!�b	)­����f���e��Z��;�����U��
�-���-����-�0��\qG�ʗ�Ӟ�>OF&!�%�������K��7�)�b�����t���C=�rL|�^E��ye��	��l�7�� ��We�C�~�������9p���hK4�U��uOGk������F��10�d�s6�,�K��:��1���g������ĸ�͕��܋��̦1f�"^ϙ�}cn��p�%���E�'��K���L*��J��Y�B���*�UV`��1U� f��),��8�;���zB��h�8��:��g[X��E3�@n(U|��ix)©�oܾo
H5�O���=��~j1��z�m��5������YF��E���6 Q���a<]�&_$���bo8�\��;��=<=�ru��.v��f�(Õeţ�e�w�5�{�:n�\�c\L��J�1�"�H�=����������8,.BA\���	^v�i޲Y�)���gn�;n{�e�6����ID�ac�3�����u5����!���|�Zŀ��3��u0a_;b��3^�n
+�+;�U�[n�sVq��E O!����d3C�[ �!?���&T��{���P���B��L��D�z����,�:_���0,X��	E�#�Q����]�K �䗃9�=(����ҕEd@�X�?:�͆�gO1��ˎ4���ml�lDP���z|��"ڑ�ߗ���7�87��n}���if|2�!��yB�`�l+g�˕�~w"��;4N�Gd��ys�Q��}��A����'´�ź�Q�d� +�T�q9�Á9��|�ew�����L&%�¼ZQp��R�8�̫Ü,��u��2,Am$�0�Ǧ6Zܻ�L�� ��lԸ�m�_C�+��
���BVA*�RF���M�i�5�3�-v�m��W��'[�io�$i�8.j�/��a��k	.=�K8�D�4�NM���� �I��j��u�z����R�4/��3j+.oen6�.53;����'����䑥�]�$����Zj���wp��I��ת�$����l@���䃫��+I~��ͯ��Md���1�o�en� �J׬K�ۂ\��~?g��g�{�2�bsHEr��6kR�a�&�י���|�����7�`�w�[4%�ac�^�84NGm��eC��	H�&���V� !��J%I�|�A��A�@����6�����p�昨���A/�w�����`X��T̘�+�Ȍ|C�(�˘��ſ�����_�ӫ���h%�9�4�7Z�=�VVХp,[:���v%���9wZ���V�u����'�"������Q0���UM�Zl>{�ԛ{l�����ң!���������ـqk�̳9���y��>Qx9-��O'��o�a����U��Qm�������� �����P����xt��X��i�-��˝>��]X�\9�a��|$�k �~�����@�Ӧk�A���Q��2��36F�%���Md��^s�������W$���+�z�3����Z�p����@�X���YeW�+7�!��3|k���Li�{ �A����LEi ���>�ƕ}O���"����a\Cq���Re�֞�c�ؚK���!_����N��cFVx�,�c�I��¾���'Y�E���F����Z�-l"��S�j�nyo'��T��T{�dZ$������4�\�r��O��W�ˠ�*Ry���n�{sxAז��%`�@9�f��y��`�0����)��=3?F}�f�1��9��{�i�x=Qm?aw]B0Ls�\�Y�նp(�e``(��c���bP�̿�_�%�ZJE�Սj[���v]���P��m�R���Y?T[�BE"�����C{ԩ���!�Q<r"el<�di��+];˖�FK���g�ʳk :z���ti�6L�T��{�,"�E59��Z3�\�Ժ8�m\�ۖ�!P�N1%�?�{TUr�[�d�a�� �h�B���$V\�P0:<��{A�-�����?�(K�i��{��������4k��9Q��;#kskAa�-Ր�@���컴[�w�Ø�͎��Y�%\�j�L�wtd4%��@�����1�"���id�YaN�э���+��E�Qb�OU���W�HQ�u�y ���:�b�h��q&l ߭ö)�Sa����\�4��ʱS�)1J��͙c�1o�����gݒ�9�cz�r��_�ڣ[N-�ȥ6<g�c��^� c�M��xua��7.Ⳡ|�s'Me��(~{�j�z7Cmxɼ��������K9�m&O0�nR�۵~}�^�@ u�Hg�EC�"_.���o/�^�ƂH�#�R��~k�� �]��;�8��< Ш	����ĝ��[*g���������#���Y�lU*4�Vli�
����y�JS"U�H�K��u$��{'OQ$�+�Q��}7�*�p��a�{p��D5�]m�z�}��{�Ƈ^�ӧ(?1�bTT�j�n�ZH��� A)��ZY|O
6�g����-Q�5���Z%�pZ.r��D��)G��M:���?!�x~������f�CJ��j~�!�9��k�~$��*	�,%�/
������Ŝ�m�F�v��渧�O�$3��X���[ x��Ǡza��Ӗt���)O����s��B�_������L>��b���BJ[�!?�P�0����<��K����%dq��3�8���6����?l��qCYCy�R�����iqv;
{�E#ɯ�w��y,tgK���G���/fT9��ie��R�ң������=�o(��O�n�jި݁�P �\?����x�P��q�ɐUK��2�"!�Lc�렣�n4���.^w�acT#{�IB5� &�p��&�D����(��;b���ZQW�&ꢞx���� ®$�A͟��@#��f�N1����0_	�`�I����a��[�X��d/�2=V�*��5�@d��y8_��İ2&���#��nE���&x)H}���N'�-�L�iN�$ T�O
z@���~e�le�-S�LлCh�Ɵ�ı�~�JN�a����ԧ���8U�NE�T��~�j�ae���m�L8�0�T�.�!9T$`����ZT�Gc9Χ�F%#�����:��3�{�W��C������^��g��zQ浝i�I��ͽ` �~5��З�]�;�:�aL�N	� y�xC�}��J_��X���`�)JOJ���#a@R^�v�N>�eb�5:�,���L�~��665 K�8�-"�b2t�sl���¼�J0\3.���ۛa�w��{v�ߞF<P?������F֞��рr&�"��0��x_؛�f��W�4��E������ٞ��}8#(%5��%$�^X�JU],� ����؛��G_"�}kV,LV\�<�Y7�6�22p�j���)�9w�&�5��pyc��T�;�u��Η���������&���)�ͻPk��_n9	~A"@Y�-?���.y[e#DB�G��۱<�u�"?�� J�!u��N�HgmG�@J�=�U\ñB8 9	$�+n:�x��F 6�JPd�ي"*�}�Z(Bu�?���l���
x��p�uW4m[|��Y:Eۜ.�mpb�Ίo$1�>�gO��tQ���U��nHZX  r�L�:hA`�z[FY8	��9�2������qibޠ�a'�iџ��[�>��UV���FA�z)ͯ5����/�%J��SWE����#��bɎ�-�Ǧ����"S�cO���/Z%�+����B�f*�EKP�[�4@�@�&�`Хz�z��:�I�����,�k��`�倶���( ���'5�����L�~۠�hP�^r���},����~�a@��Af�Ǝ��A�$�5�pk��R?¥5�W��]��,�z5����[_ͱ�Զ)!4XXd!��k:0P�p��q�'�X}8���������5�wS��?�p`S�=��bPK�6����ﻰ�(0��L*f��&���a�;|�x��������J�2�<Y6����d�v��K�S�*Git��6��_��cQ.P�ǟ��N����C����'T6�o?�_�\u�^�����𞱻���� �zd�o..��~}?�r��_������pa}/WC��|�Z\�+�"�@9j& <>ˀ����v$��S��KP�~�Z���r�$�����y����Rc�q��^�==g��*�� 䰔2��x�5y�.P��F^�pa�H�߁�4Ո`�c$��X�~���ۊ��|.Mg@�n�$t�M^�B�X�Zc�s�rZM����:�c�wk��[ Aa�>���t85�����f�_�� �'��)[̀",㗅��)2���	�YU��+�#b1���-#�۴L�ǏQ�A��έw�[�C�H{F��o�XJ��ky�1���AN�&g(W�Q��!꾴��4���[�I6��,���d*B�x�����n"��?��A~�őR֬›S/��|��[U�9}��(��T�W�^��IES~�Ml�$<�RLuojf�$�碳����]�Ki����,n΂J��,-�W$3�zd�y�$i놑�貯�OM�#�̯��Ԗ�:��b�l�!g� C�8���;�2�Ϳ'��K�1-l����?!��۞�l��3�9���YWi�MQ�5�
9�X��W����MI�gф���J�P~�#؈���o3y,3l��#=};�-DI��s7�wn_�~q̲;���cs����bk�ƃ����)�����	���,�v/l"s_{!Ze�W�W�W��n�"��
��N��+(�LL�Ƅ�� �v��ݫ��v��@h���Z�P�����8[�/��<1�d8�z
�N�Ǌ�t��Ҷe׃#�lb	�&�5�����F_B�;ޡ�k�v��D�3%�����Dh�s���zax�g���4A�.2"�(������*?zZ�TA&$q5ܬF�\����N��;�,5�w�f�~B�5������a�ȁsV\��&����� �
���D��ٲE˓	�l%��̼ƈs)�g3~ߴ���8��"��Uh>�!��C���r[����)M� �=����p�C���U��j,Y�{Uw��<��(G�'W n����!�>"�^�D��ק�q`(�������oXT���@������a���4xt_�3�)N�8���;X@q�^�5j�����3��_&�<��\t0	xE����È�wa>arͺ^�^��e�T�u�ꞺON�O�B��	���*��-����P��`
�	�2nU���k}�R��Aގ����%��'���ǐ=�}Qs�5b�6(S���Rp_�d}�5���(,�����v���[˵5L�����L�#,|<껦𤫐��k|F����pG�.��8�]�ƀg����
9�O!�����3�Cw�D1W�?'����j�d��}a�a{A�v���TW%v ���n"�0?�*�j�z��nRf�0���߳�`��O����P���4&o�U��ЛK:I��x��/������تU����8�]��s/=7N�pQ�Ӣf�h��"�ڳ��{��8S}Ec�5�b��J�S�������G$�t���K딟�,�Dǜ���F�ч���'kG#h��4���L����[)���ġ�=]6ƹl[5!�vo��R�V%w�D	��(��� �$����_::t������<)�x����b U���B]}
�Z,��_򧇪?���d!ǭ���P��`6O0*V��6K8���	�a=rm�l��P,vb/@���a�T�b��
֜̿��B_ |0Ʊ�m�������˃^Y:�0~o�3��/#�~�
ZNgmw���$SM�'I`8�ۋU�V(��c�2.�{8d됤vXt�5�=�q���o��fx�:Q�*�m�N]:�a�(�
<��MH�久��k)*o1*���ʽ��������}��g/N7=WA�=�汫.�k㣳RG&����)R�Ñ��E%C@�7���!��g�R��V�|�mY��tb���*-������X��p�*.�S����_�u%c�#*x�B��x���D7lS���N�5�ݓc�}	bY���;��b�4<��B��.��+�2!��O�,q;l�����wn��t���"��I�?��(]��J~�7U@�z�J���9��#o}�W;�����o�@��$3��� �7�9�(#�+���N�͖7���RF��]�c��iv��;6����DN0�=�v�jF2��b�j�����~8�����kUʨF� � =�uP�S�kذ���;R+�׊��\ʪN|̸�'��!�G��z�$��K��&�JTu:Cј��NI�,�1r���D�=��J.��I�?�BciUB��^��'B��\��s��G琣�{r��κ�|�{�_�a�a��e��`W4�;���P�������1�i�jpKD%��ݹ�բ
����^�O�P<�O���X�8��K�'.��o�)�p�
$�
�h�iȃ[��%[��U�L�{7��!7&:�'�t��_ʤ�}gJ��ǟPc���ԭ��rx�,�;�}{w	[cʤ Ǿ�@��9G^
���t$�4�4}�-O��	,ɛ��$���_��=�7��jU`�	���3ĨX\A�O���[���t���jhaBl��"h5�h5�D'qܲտ��fo���	�"�ۼ�1���G�\<�1��JU:��]��������$��%o�B�+8��v�I8�z�s���z��#�$-\��6�l,�dloWiz\4��5ϳE��`��X<ɫ�CpS5��j��J6���V�Aa��CZ	'M;�?>�����Y	b�������^T�&
x���Y��g�|�Z�[�w���xJ�2�a+�>MJ�<���y����PZ�N���B�a{V��0#ǫ����P�9������?���D�di��j����F�qvjݨ|V�|;���QY�H^�OP�� c Bb;��ޝ��8�Qۑ�X���l����ǎK�֥Һ^�:�S��xw��Zm-�^�|�mkK��EvnBS,�	u�Sf]�w4��<B�hۉ�w��dB�<@Y`�B�6�o�h`o�5`�!�Q���VV�À�oV��\o"����#�Gg���So�2���_^�:rG�(C��t3Gѫ�߹���ң�(9l Ev�_��s2϶�~¡h�E�ٞ�S��M�\�W8��# �Y�����a�Bx�(�]|�^�)P�lAܯ�^1�v�����ڃAY�nC%B�{��W��S�������3Z�������Z�Mj^���QEk�?z�ݰߒ�Z�-q,W3�Mȱ�Cq#�N%  �c��j��X	au�W�Қ&XB�&��|���ҷ��R�������W�\��������zMgr����5��r�*��d���v���N�K|pL�"��VLʵ�y����Suհm�i�u	ƀ� H�7Mb��M�O���MHC^�x���96�}�+<0M'�W�v7�#��_�-c���Z��!y�G2'=_[Q�y!�v2\d��K;8:��4��ޫ�&4�e�A%�u�A�r��YN@���}���1QSf�ں��0�qq�Ӱ�%�>��s��8���x֋V}*B-�׃M߳p5H��g���Sڋ�z&N�$hA]ڡ��)�"k_r��<�� jf#��
��9�8�W�7��2���1Y��d��E�ڊT�G���V>��*�+��>v嬸6+u�L"��n���!$��!���?+�hs6�a���(���"f�p)'���r�/2B�M�2�'�����ç���0$��Y�ω�Y����oV#��-rL��Z��D�� �h1���l$��`^}q�R�9MA�9G�<��^���߂ݙ�9�̽y�c{����P��a7�w�RĘ5]͒{���H`{;��{�h�6|u[�ޙ�,���@=;C�H�x�?>36�M1���l�g��y�R]�\� ����M�򧨹�-\��̿_K�>Ѳ���[N��n������Hp�LQ����\\<q/D�Mn����[�-KRD7?�>țM{���WE�t�Rt�3	/�s��1B��@�1qb�n�@R���R�8d���%��حא�F����l��W�_� ��V���zY*�����`�O�[�x{m�{hƈ���I���h�<�k�B�������4���Ջ/�_^w�z�ơ����$B�{�Jdn�����A֔$Ԓ�O' x(✀���%�Ѱ-VU���Ak��~X�J�U�\Z8xu�\�~X\�$�ܰ��������&�KM�Aw����_=�lln�m��0��d�ӊf��]�n4�gb���� A�ЖU\O��2�����-���7�;<��H��>��͉3�H�d�*��̺���I�u����M�I�.<�j?���^[��N ����Nځ��{�#���ʳ��&3��e�9=����F��s�ٟ�η���dg6�RMҷ�6�CR��K�%=Ӻ��l���CB�?}�Fg�3ݩ�qU�\㶏�U��[�
�!``�Q�z.��g�2�bC��#1��-���I7\:��Ě��0�x�Yۈ����b���R�!�ua3�n���y�����oEcH�� �=�����(�-�N;��0�n1ac������)<}��}*%
*6h�!�iT8
��T�#�B_����PW��Z{�ʻ�!@2x�Ng���3Q��0���ݢ���f�^Q�M��B[��篪_�ҘX%sˇb��� ס
��M�k�2kNmh�8M4�[AR�T]�q0���/�tS�.�m�ᗖ����{�t���N��7y���Ԍ��HՏK���oj˴�]������Jy[	��P3x�3�l��W�����w c�IIXZݕ2NE�����|P�����`�h;��e���kʘ���Gmܔ�����jŭc��W���:K�i�y�gG�aJ�y��kqزmZ1�N�l����S��#&�5t܅����*�m�A�^����~��h��o��´�z��lf�Å�qRwf�F`U�����HS~�G��_�\��cA$M�o1]c8��(�>=�7�v�gW�{v٣�#�/y#riR&�k��n�JA ����������-�$9��/ɾ->���N�ဢ*�c�a�A|��K�M�i��m��� �SIe��X�}NQix8�=՜��cA
�eF/�����zR�:K!aU�fl�q���{�&�U�NI�B�s/��"a3�4�����4�7�v� ��Xy��h��Zkq�;�y��7e��Z��t���Q��p ��</<�#kgk�d3,GU�Uȿ�lN̩%��s\�����M�x�E�w;U���*|�aK�%ɹ*B+�^~fm��,�&N�s~�BH��O`����]��_[��-��1�A
���+AG�L<X!vr�;��iN6S��7���O
L[.�*	��	Wa�-���'q��32&�B�&|�[vd�SE��P<FN�<9cUZ�Yh����0�&����9m�J� U��S�����e":���W�D:�כ��&˂�����P����F�R���m�pF�'�׬�1��>n��vh����Ƒ���~r��.��u��� x�5>k[(�������D,,�-������Tt��srF &�S[#a�m��￫-[�D�a7*m�w�:E1���v������0bl�;K�����
�/���;�o��n{���Q~S��&������A"^T�r��26X��Q����nxG�Y-M�e؍R��&u�k�1�)Oj4�纂T��|TS�����]|����5��ܜэmW���q���#��3DF���e�94:���ѻ���X�fG���fdT9�́/�9���P�e�����G5pMl׽Ό�9p�F�G����xC���#�(�{(�A��Z9­����Qߞ��dq��,TG�\�]�8ޯw�� �3��j��{�7��Z ��x�p��y�i�~C'�m��4LE��@N\� '�Ty'z��GP�w>���|Q����K�����g����nh�J�
���.��l$X
�� X)�&��'�0��`4���l���i�A��v��S��Ж�w�u.l�����ޚ��+m�j�w���J�fZ�Y�6�j�ѣ\t�m˥��
�'�;/��"���̚�ϔvi���S�ZG��6CJ՝j=��Y9+����2�g���jV��u��rb�ǻ��i]Cf�E��J&c�;G��-Ym��o�ѥ~[��`o�z��gC$�$�k{L�"��ʥ��2�R��6�A�X���H������0�7���P�G���X�稅689�S<�ۋ+�" -�C�0ҡAK- ��%i�2��C�0!X��Lb��-��\lx~��x�	[��F��R(w��JW���m�dN(s����@'��(�KK�S�z�l����Bb0
�QP�ֹ}B����|ܑ�o�? ����ɻW_�I�,�
��%�,_�ln+�k�B[y��+u`��*��(O�F��w����v=�´?[(�L��1�p���#c�!mXq�?ɻӈM9Hى�_sĸ�Sm��TXH/P�*����Ԙ��a8����`��}p?%:�~]��S�B<���3�n�5[�^QR��BA\X��<xi�muf(��o�s���Tq��ݵ���O~{%somx�߅R�%-�` 	b1@�O��(�� v��1߄4v�Z[Y���|ڔ\H!���J�e%XK���5�0��'&��K1�1��.������R�Q)�ᦠև�|��L��:�����H�+O8������A#�<,�ljd<�V�G�Yq?d��B��
uƛ|X�׭0c-=�7�X��[��^���60��0���2�H[5O�kp	s[����LX�0�k+���V�ju�%���ӏ�&��Þ�#I���t�"�ܯ���;KH��c0�`)<�Fqؽ��p\"��� � �3{����*=�U���:�HYAߏᯭ�gF��7���0%�QUY}�5yE���a$Pۯ�
o��?�%���Ҟ
˼���A�K5eN��g/��D��bKtD/�~��m���KS�(���u�*����nH����eF�p"���xm'G�;�Jm���������K/1����(�9.�	��n�m�ǜ"ӫg���Z�x=�&u�`H��/
�'Epbv߹}DQ }Z��x�nh��@�ì8┄�����뒧����l'�+����q��9\�ޏ��0a ����)�~tk�o���&�c��2~��xc���.�w�^kz�"	O�SV�B�	��(���"������j,�o��4�T5O"���}�S�j�@�6�`���~��N�-P�ϊ���g�#�15>x�r��Z��xPW��]QN?>9��c%�%���/Փ�he�ۑ�����u*������DjlPk�okw�m?��#�2O��JX=g��g�]����&U��'�3��'�/�W��� ������ �b@S���kV[�� ��m�uu?�d�O���Ug0&��k�j�}���t}��~P�(7fX�(��tPX!�:AW�%�Zg������eb�ȃ���2��F7�B�eGE,m��ښ���ܧiL�e�'�
g��6J�ˬ��r:=�x�ZD�"vPN���Y��|Q��Ύ�lM(��;Km'�������[x�bF�>���d%(Y&��|�3�v�}��b����tJm��M�Y���{}�I90p0�(FC�o
�{1��.�����@.'*%x�-�kb!�#�������VW&d���&��Ƨ�����(t���j��r]���
r\b@��\/�n�z@hf7t�bEYp>�'"v��p���1{���ZD~U&��i]��S�}�UEp2��&�#f��U(���	������u�,�y6ҭ�4����v�����*�v�<��
�Q(�f��a��,���4�>.�S���O����+*�VB�T�J媊�{v#��:sO���˱��֔���"�hD�	��`��!� AW���� �%K�R�#k���&apUKؔ$i�X@��ߨD�>�,`bmHyE:� ���Z /����$q�gAl�M%`*]�J|�B���>�sF0�(�?e����`���]����n���I�W����WV���삠�Ŗ`��v�������[�W���_�%�B&䢵���w��A#j��J7ϳ�����z�a>�ys`2������r�0s�#m�;+f�h�8���΄�̰��Xn+�mP��ge���A!3�V����.�X¨Z,w�`�V�Z����?F���Z�St��6����B��pL8���F���u�SF�� ���˒*T��h���K���Z��!S�>ÑM����nHr�?&������j<dx#XB�<�V@��b_�Z�K��3 �A�B�b$����� �f�v��=��R����+��T��ɟ>4����U/�ԙ�H\$EZ�3ll����c���D��	�E k��6��5u=�҃%ְJ3�ʆ{�1�Pޢ��q4���ƻt\������M*�N$ �F2�ΩbX׌q�TT�W�*@
!�҈��^�o�䨵 ��5v%��Lx��>�-�e�3>��!�O���q���|`]P�8�8L�L.��P�md�	v����Gq��v8&�h�=F�N(�Dn깨D�唂���(�H^(1u�H��aF���yI[�*s	��������������T\C�b	�_YlS�����l�f��XK�f��~Ld3o?�7>g L/�%~=s�/T���#�z�Qg7�#�=8^p���t@����1��F��7�LD�A6�RA��P�v/�c�>ET��6�>�tla���
�D����L?��4{�^�ĞUʐS�'7'5B�����S�Kd�lP%.�p�%r��+VĠ�9~.}�w�/�gǺ]�G�"A\+*����i�\3z)r�WG������}������88�?�����q\��ی�>\k��R�'S�5
S�}�"�~�%Q�Z> ��nc(.|�n�R���-h�{�"ԩG��(�������f�`�*�����7���M�O�N~������Wi��͔?��<�_5����7ϧ���u9����qk��=����|�'^���}V�LNՂ1n���+)J6�߰��\<
�r�Z�xm�C��mb�F%-<��o� l��:A8�/��K�0;q�.��z�eR��f�;)�h��fλ1/ʣ�w!r�0"�~�ř���!�滋f1��TWA�2�p�tm����I��nv֟��e��,a��t�q�Г|�=�m®n�{�{��� ?q��a�9�r�i�Va4��?�;��r��F�o�o�&A����|�d�$6�f.g�����J�?2�4�2��j*�B(l_�ĽM����m-x.Y��U�{�����ĕ����6����s�]Pr�;���+���+qlN�z�bV�p�:'l���v�aW���n_-K�z[�抡vfn�Y$�W���mYB�|��:���+"jī����ڭ�8�����Q�OB��t����eӞ��s4�8�O�=�>Ֆ"%���Cs��}�4��A�'���������?�0ɏ�<#ã[���n%����#y���E��93p�Wr�oma���ڷִQ��J�D��ϣU`�-�FK���n�pDp:�y<\ZXY������� >6����=M��(�9��;&lА�
~�տ������q\gc�t^F����V���U&�faƷ�EQW��<(��Yn����~w�ݵ�Q���`�̖v��-����i�+ ��Mٮ�b9�a�E��R$��
��Y�*��q_hE������~�=�����٢����%L#�]�Xܗd6��!z?�����!5�y��,L\P}������D[ȯ�b����2��}�I�ѾIJ�*��ϱ��6��1 ��j�MD��!�J�*�*R�u��h���c����ۖ���n���@����P@�?2�P�Y��/B�$���h�+a��2��T���_��)!#�6!�`���|�f�\�<��G�5�Gi|v�K�ܢn�2�"�A���a��x�3�%�C��~��}��-�G�T ���%p��Q�k�=��!L�A��C��0]��$�]�Ps�c��D��X6Rl���"���7�[0/�0���B|�x��@�����s��/���䦙I��1j`Ox{9���m�� �d�����p�Ǆ7"+�[��fsA2�ED�n��f뵤�eǠ�Pc�>W\�&Ql�:[~0YƠ�:3,��ơ�/�f�	f���r��E�>�5����P�:�kU�A�/�s� a�T���:�A��JD���JU�t��˔�+��NҕD����Yi���nj�WK�rPN�aa[�<1W�f8Mo�ᑤ�K�*�⪅+�S�Ο����6hmz�XC ����1�u�}]��疂���qU!2�4�{����؝��IyT��,Q���/b��gq��U���j���O�$!*�^�}AS:o��+��y���=�|���cT�SS�-ڋmҭ0���x_.�J���-Yɏ����,��&��ۑ�e��ߙL�"�l4�W�µ��(���%ƃC�s)s�2z�'HR�:��]9��`��U���G;��l!��D˕+�v������m�_��R2�\��l�k����0�84ƯD�(t/�F�H�Kx��vǂ-�C֠�� ��l�- ��f��6�<�<!���M3<xJ;҈�-m�ySk� %Ģ���	px)X3w��a�`�����1��/=�Ȱ+�wt	H��@^�%dp��V��p��ɽ��\�c���XJ|���ӑ���|��K]M���;�6 �}���7$�egAU{߳$[s!U�%Z*�)��*%�z¨B����K�:
竊�Q����E��8+�K��&j��."�'#��WI�p4\��1����}BfJ9�裎H;C��$���7Sn~ڷdhpGr�\ɠN\�?��{ˉ�tEA�w���mp�1���͉Ãa`�V�h�V���.�D����c_��q���kYĠ��>(t�[��#�\$��2�'+���8LƏ�-&~o�:Z�"�s���B�c�.?ځ+��m�q�]
�L�~^�gxL ���.[���-I3�vT �b˵8�h3�]�zE�Qy0^Z��4j(�Eͯ�˪H�ry��EI;�I���l��u �1�,H�A��t�?��W�{.8\�>��k�����Ƞz�s7G���{>���}W�-���[�;�-E��C:.Ө#�lrIy��3��R�{b������H��y/3��o���*殕ӌS��#5�i�dADBF(T(	Bpi�OOI�8*J��Q�}�Ѿ�����p��ʊx�����
�rd�<֦5}
��{��`N�4�ZȷO��Mb����oa��)>�Å�!�Ұ���f �.#��s�H��a[����S!�lj�Q�>��Z�iO�ӣ]��XXQL�ez�X�ء�M�0����(gJu�X��4����	�Iyj��9�e� ������êCǥzK�ގT�!�v0#��1,g4��noV�߅�X�L�k!�୾��祈w��[D|���e��㥿X:2�v�OS�jNw<������E	ׯ� ���s@#@K?L^��<^��2*��ajV�Q��\_`Uɜ:Tf����0�����;�.�PD/QW$�%b -���1[����͔����ښ6I֡��)q���B9�{.
7k,����?k�1�?�FK�H؊�>����R;���\�V��~ڼ_�= m��|���#�|�V�!2=)��ڸN��Gt��
&���U�!Gl��n�������sF>ּ�6C�R��b���W�<�@t�S��{�ߍ��s�^���M܉�뙧%ݢU��W���c�Ѻ�����W�3�φ����[�Pa�	�p�j2(�������Ġ� ʈ��P�0���1�A�J Y����J�M]�x�a�ˋ=��=�<ɻ2�ab��B����,U+p��I�Q��|��$��	�~��ō�iGx�%6B���Hw����8��;�.C���>�!7Oba�+դ�UA�ŪÁ��F%�G���8i��e&�APx�E�v��|Ƿ�Ϛ�Q����aE��E�c�N�6I�ռ�15�N���Ӝ�8�h���c�r�ТK9�k���+�i�X	~���s�I����8����#n����;l~?>��x���I&3Pۯ�@���L��?n4����"�$���n/�����.���tv$��`=� �h��c4�6��(��$����� ��]��^"#����|��1��
,�ϑF����⋍.�ރ�fJ�8��-+�_��	(D��4;�m=TP��kR��l�G��m��Iy"�6�����l/Mkň�PgMȷ�d���ϥ1�p�k�1Q��[���~����7Ϗ�^GV�����.�	7oS�3T����^&�wf_ղ������pA�Q���v�ij.�8�0�� ��#�ޮ��JQ
�Y�	��,��Hz�`�bȾ�x��T`��e �et�'�W��Z�=!�P����gE*��%E;U���C,�U��e����|sDM1K�nѷ��G��3��f:�ƍ�z2������d�r)�`Q�4 �9[�3K�HG*w���[�9��4G7�{���������֙�����?v'���+��̩���;��XJ�t�{hU�Q܂����XM9	���c��S8�-�&�(�z">]��L��?��@k���z�>��1 Sik�}wOh�'fk/��M���ϰ��j�`~w�5e2�M��P���&r��"2�7�϶�h*PR�hZ[��w�(��uؐE�>D�� q�L��P�@����"�U$9�5:/{M�3L_��MA�ُ�k��RAe�1g4���ǈ��(������Y������<�izf)Y��n��?}����x��8���B�b�dዕĲ�!��,}�u\~!�ΰ��b�{Ցu���W�P��[F��f���ى8׌�n�۱ЮUL�n>VU���I�v{���e��y���J��*p��QN�^�:9��^�"�< Q?��S�.�#���M�I]���+�**���!,O=�5L%'��,���ֱ�s�O��ť)۽4o���Y��7�d��=�6���Ӂ	�8ۘ�]J�i�"s�B����a����r�ф�R�+��d�Q���R^�	�[�q͠��*���~��o^zJq��p� e@yG�9/���;yߓ�&�wҝI���,Z�Х˕ҫ�0`�	��px�9�3�����mp�Yd��z��s�ٜ�����fYMRD�o����F�c2=ں�
P@�Ej㱽SP�72Cx��-؝c���c�"�/nÂ�:6�����Q;H�ci{{���5Hl���#����xhQ�j_�g�U?���;�1z;$�o���j�M��r�8�b����I�����D�?R|��Q�C�e��z�z�Sv��K���u�!� ��,V��)���ߴ �R����VB�C���}�:��BĽ8�v����F)V^�e#�#H]���e�e}��/�WT�3Rm	Lß� 1<��,���Y�����NlT����b�ȆT��4���n���W<���CC� ����;iB�L(�,<�{qe?�̖��e�M#�RC���7�e��]�z�CWJ(_/�����9?�#S�Hl	��S9�����1��{��ՃЂ�`{�Y�>S��媣K1J�>%*< /aU	g3�pl���T�x@'��F�%�50����^�����1���w "��푵�9�a����tj�|��,�epK�)�HB���3� !L�4�f��m\K����E�7.����4�����,���v�A��Yo�.�G���x��GP�b�
6�Jk�jOy�k�nWk��NY����Dz�����K�T�b�չ�,M��8=�r��z�]�p�ԘN'�[W�B)��\S�B!`�_�;�?�A��jJ������I|���Eep���8�~�|jk����]�ޢ 8̊�j)����i�T�*���5���
y�춲��UOxj�����;�XS.��W�!����`Ðs� rJQ+a�'���d%l�~F�t����E�Q�lY{xh�&�X���u���_ÿ7��$:j<ӻ�m��i�r���W{�#[���$�������b]��B�_�1�#�B�&����Еg-��}w�+�Ģ�%n%'1����V��\�s�bq�<�B0������7��G��yKv\w@�nNR�� �Ɯ*��Y-d"���t��؆�K=��C�n����/��У��I�ub��H�H�C�A%ضF�e�x↜�V�=��ab�1��r�%V�J�5��#�[����y�e��P��p�}�14�:�]D�T�/y���˦��d�)���=��?����D4>O��6
"�Jhx{�m�d�YY����@���R��I��nj��F:�s���-#��}�VO��э�|�ˠ �����)��ryU�xOz6w`��5<���Ŧ��e�1Q�[�~�)M�?;b%��q>qOd�,��1���L�K���MX�$eW�ҿ��,o]uzV�*��e�d�P�����/REK�U�8�.�V��M����ړmt��X-���ja~4����`�/�M�j�󃯧�o��ߑ�@(�Nu����O��w՝����&�e-K��W�g��t�o�߸�n�>��(�x�z�$
�s�¨��`Ǻ�[��ޒ҈�v�rW�q��cz-p!X�:|�ԜW�_��L�P/�ed�,U�PL��|�(�0�l�F<���G�M���{
�� �y��R[ư�{հ�Y��>�73�ª��|�A�]5+�֨^���/f�+�Q�ӭj�/����6.Ў$�D@#(��g��1S����S��V���$�b9Ž�6�=4(Y�#�;h��L�-�Y�1t���1��*4����wH�b���F/����se?���-8^���.�k"ao�-�9��A����T6s:������
]��F{��rSC�Dq��)� ��|@�x� ��_����Z����u-v���^z���ͻ��w�:� .����M���F`��Ԃ%��w�	.��IU�K��(�D��#�At(��=�����z
 �!��d���m�H��;�֬� �������������`�,���Ƶ�=L�>I�\ ��!��4Ȓ[a�_'T�T��o����B��5�<��e�G�8����8��(ca~�o*��z
k��޶f���餼y?P�<]v17��%��E֨�S�ӊ}?m��� �8�+��h�~�<��7F�?0n���E��+�����JݼĿ�<�ң�x��e9�����[��K�iv=P5��?�.S�#�����k�H�-��i�ӅmY��p}3J�Cv��]�����!s����xw�`_��� :�-פ�RS�����Z@��
�]�+���Tp4��z�:���+�'���1�3-����ړl�϶�˼�ʄ��	�"$��h��û:쫣�GX�'�9�P|�_6	w����v�1t�g6��9%g��x��%Rȑdɞ���$J�:�O�ږ�a����L�ef�-̣M�FZ�'�By1��^.�������L&�;�S�>9r4R�D0N!d"��W`��HѨ�ϱ���̾���%��C��un�WN������m����O0Y��.{���Rr\^O�p�!�+BK�H�:�>�Uuq2`���=2T]�fFϾ�8�4�3��XF03#�!ݺ�U��%�[o"�"%T����F��kol��B�/:+�߄~�Vj�,sk�����կ��nKj_�����b���0��>N5Fg6�!h��=t�"��1����-�+7sd�@�@ߤC8�	ɦ	`N���ob��S�C����晋����RY������g�l�����m�y~��TA8Z�W����k�o�^�$XM>���������ž��߰����峳�S6m��a{��E��~�� N�,�o�nX��<���=o4K� ����tR��`m�9t<�w0{p��[ýd;��� ?��a�����j%���`𿶢�(��}r��Ŝ����A�����Z�;���vu�2�%�l�O��n�R>Y���؛b=�Up���Ec���.uǅ9��4.�E��K� �`*�c6�}���I|^Y@�b��C�@	I�H��T)���[�g>c�4O@�EX*!��7��
��Y�/�.+�����E�3�&=I#�|<��D��/a�5Z��osd�h	H�p��2.��H$�!C�	,�H��r�!#��<聀2:T��B�݇�xnDB���상F���+�?�ŞW����%bv6��|"ǈ��٤��DG��w���᯿��e����<�4�[#|��DYq�FܜJ�ķ�'�{P2�i_��.�K�t_J5� '�[�a0nU��%6t���I��чAG��?�2-淪&
�SO�����㒪d�Q��7���Y݅t���͏o�Շfз�I9�ZR�_<�`��:��QD����ƴ�*�-�F�63$FQ"���Cv��m�*�,�׊�숈���#��̜W�-����*�@�`�V��/s�ek�q�xG���*��]�Et!�4?&H�8˽�mr�Ι�+�*X��/�Q7�p��B��)���y;1] ��&�\������=�i$$�J���?�z �� gS�,h5S3`8���&u��-�t���҆��C1e��'�ꄪ�O������<{��P�e$zq/��v�-��.��~f��1{�N�	T��U]`V��ԊE���'�$}>@`qs͖�6�
exhL�����Q'8��G�p��?�|8�57�C����`�6$h*&�5Ф�/��-`"���R�k�]{�l���0�m�y����g��U_���HJ���v�i�+�Gߜ���P2u�'�|D��v�lI]���%��6��>q�1#���,�S��/�ۖ�eT��?-YЕ�VyK�zj(���Be�q����I�6�%���L5�{2Βgd�ˡn>��=��ۇ��д�%RPB�]�S~2��<�x�*X;;��R?�kԬ7#&�\�n��󪙓��"����v���I\����;kDm[��W�?<+��'J�g�Z ��٤��׿��Z��3-O�e��j*��4[<�����6�Ǆ�}kT���Ш4jj��K���
T�q e �q������ޟe�69(�����Z��j��zf��,�8�`���/�3�B��6Mζ�nw�ꜜ�fBi�h��I�<
e�Ӹa�=��J��ZVXg�b�N���̬TH"��b�X���2/H�/Tv�1m��hI���U}A>݉Ϊ��L#��*��@lst��1s��$q�4b�i� 玴��|�ʟ���&��ll�s�c�_��Y����]��:�>�sf��i���5$��kS�`���:�&'�S���"��şǱB��)`ǈ+�d�[7UJ�4FRNs|�9D��{8��n&�;8'[��f��m�l-b����ђr�l:?6x���MZ�$�ǫ�U;qJ�Pҕ�dw���p�Ə�Jz�my� �TJ�G۸�����e�#\����	��\wٸQ�O�B2ςg]���4\�	,�#+A*���.W=��p���3��`���~�g���$���=>.��|<��==�bL�Xe�%D.N���w<�f�4��W�iV���ΒBQeK����K稓Sf�
S��(�z��?���:�����h��s�Uta��D@�pBg��lGnì�O2����wS�{7��9�t);.D�aӞ�+Q\�׎k�J��l���Z���?�픗L|��oI�����/n���n�"д�zUK���t�QuC'���r��B�݌0A��.��sF��|�$S��`W?��?#�>!�Oscސd#
n�Np�H�';�o�I��@˟���in���ɿ���y?�Z���y ��#>�7#��,o ��;I�$� �-������V���`4�
*���a`{��n�Yxz�!�2�=� �#Dv��%�i�_��5D��Й��Äx���j�S/����Pr�$�Z���gz�c���k���� ����Sp��k��5�w��h�|�i#���̃1�o��s�&�L�x�S��.W�)��PV�i�kFA�&N3�!O�b�-9�J��|~Q��!ӏ�~��*oP�y�>ߎ�[���h��!Vx�bi��g!��M�MB���$R�O�hKyE�|�D`��/\��w�g �v��}��7B#�Ƣ����*&��*�}(���� ���ɾ���yo�oU��|�����J�bWz��@E2{�=�Ĭn8}�o:`g�5)�M�#��޼Cc��~},P#���\@���8�sKN����������}��׀u�Ü��@�Ӕb>��;NB��{4S'IU~��e��(�R�0
_��㠲�Ǜh$2��Ko[���M�C ����E "~��S ��{,*8V_��60��:�Q��� �OZ�ߏ�F�bCʻ��i��n�w�ۤ6�R]c�I��(���N� ^�ڮ�詶>�R���U
�(����Г��!UR��u*�>���.��������k������1����ѕ��*�u�W�����n2�ct�&b�flȣϛ6K	�^�T����L {��4[��� WnݠW�Q���锂�W��>�f"`�9��S��-]�R��gj�(Ū<U���ߐ��(F�iObq&�nvƝ��W`�����Ǡ<n��F�����܉`�R67���;�9 �-�0'�>o����9��~���?/�b{0��`�I�7j;�,��v�_)@�-��)���F�Fp�ø��j~Y��rO�F� ����7�,8;�]�T��+��ip��n?���Qnֈ:����}B)��֝����ϋ�@>���lM.:��.֤�B��5����5:��{�A�2���%�UVe��}�Z���6qt�-����f����O�h�4�"F�:��q�|i�����O�o����\8��*���,x���,wDJR��a�ξrD!6��T�'��]�Ľk�Ps'���kZ{!t�R�r���I5�Te�Y��Z���Y����A�BN��6~����x��W��N4�\�O�0]�q𘕪l��=���������jH��a����0�3�gFqz����$;�z�zA�Y?r�$)�0��1�u����N�Yl`v7B�Z\��=�Ňs�C+K�>6�k�[������3�䷂?��>�PY53ۏ�`�C���G?%>g kan�B0O�6�0c���F"�|5�����pY���M��������SG�V b"�<%'�����>�5Q�)ܲ΢Dz��DS��ޮ�͜��R��~4�����
e�i郓���D�슧*��?<+U��rXyF#�`�K��V4t,�A��8RQ�&�8�' �_~�U�ы�4r==��G�02+�ì�eo�^	��_�Tn�L��ۥ简��"Y��Y���F8��^j��k\A�?/�I�k�G|wc��>m�x Y�Em}��2��C?m��z�9�e��'ro粻L�2��-�6�Ƴ9<Q��QI%	�0���1)��6�Ţ+a5M��	��/7q��zs�ֻ���)�q�yc��D���f�h� ��)[�h���h0��|����&��p����KC�{NE�g�� \_g��%���_������W��pl�w���I1��}��f@�2��`�a �=;-o�(�������Lq�Jmjk�!,V�ml�,��88�I$s�^	�����N$��޺*jⵞ@%�c��Z2p���kؙC��d��?��e^�
)&��'��κ�UQF���#���H�MSC;�U�%���Q��|�-��Q�UE���{�1c`Uj1ev:��i�q���si�4�.���ow�Cwze��\a�Af,4aK"H[�b0��8g6J6��_ˢsx���T[Y�1���sC��xu	dgBMO`���6LF��]`ͭ��{�I���q���X(�1�EM�W��Nа�j���"��z$����G�\Tl�ͧS��Ʉ���S�����H%Ъ���������9�e����b�v� �,��.Y\ڿ�)͠�Ns��/�RO5G:7s��7���v�rf6�c\�ϵ�W+�"V�PB���Z�G̈́
Ш�I�G3`�(9WC��B2ٯ�񗨎��@��i��=��0��rOi�w�r�2����|����+�lW��R���l��W㥐ɃK�Ȑ�Qj[��b��5ݶ��W��J��$ɉ�f����o��|k�e�׿T ���N���?�ڏ
9"Vf�Ơ�A�6;U"3���4�J�t��F"��õ���j2��9ѭ�q]:�$d�6����G��l%(��μ���Џ��MU#���fH�ƃL�u�]��%|�Q��SD94�7y�<��_�˸��褝�~v�Lxd�J����F'���nK�*�j��|i*W�k������}7I��LǠ�\jRf��_W��$��8���⇊(�j�p�QįF*�&+?W�?�Ͷ�˳h?-�
B�������uV ��ٰ���)j�!���@�QwC����	���'h]��>���������z�Zk8lc'T'�����FxC>��7W���I=e��vOϽ ����l�gߏ*gK��\=0�	��2%ˋ�4�]��R3{�����_�W	ǵR��C�9��X�4*��,��-Ȣ;��I�h���c!	��C��q	s������MxX��1�z������q`�z�B��*���YͬϢ���1��ު2B�R�-@m+p�HS�w�m'���(ϗ���g���|	*���=n(m^�g:�a�OMok3��c�ً��ٍ�;i�M�aQO��bI\n���",2�L3qM�ބ^gw=��3B�����̙_@DnO�~���Dg���lس����Fa]�Gl�o����&+�`���6ʳމ��N����0����⢽�/>�hI�R�3���W�T�]~dݟ�lx��ZV	��p��6UZ�j�KV��Փ����4�S"f1#�U�.0 X��32�1x�~3�Jл�ؖ�7c���u�]⿸6|��rb�������&FS{�6��S�p-������ÝJ�N4!�m�]
�gaV�� p�Lt�S� � �C�j������綄��^▋����q�~�Q�jsxkd{��G��K9�X?�H�1B(,�EŢ�Н��M������~�K�h��W���R�A�Mİv��'��ƬyJo�l�C�SZ��&gI�kO	������NQ�J�(��T�r��M���+]����1�L��8N^�-����%*� �u��>��2��T�$z�V�ͥ��c;o�:Xd[�D���X��=�w�0�)d=Cųԋ<�=��RY���9wE�2��.�p_�g��^ɗ��v�3��(4Cn�t���28<��l%:�i�٢or�[�2D0� �Xv΁s��5{�*J��4.x�%�	*����.0�X�_M�>�k�R6B�v���2r<e;��|x
`o���<+V8��0��!�O ��Ă�_���$	��x�%��k�����
�R��<����rr��#��������v�/�{{��A��Ë6ō���
��B����5����{���\�8׿��PD��U�����P�M���<1$g�9!�bYͮ���i/ǭ�踭��e����صW�zGU�z"�������0V�6���Wuq���>�/}�3���������T:Z.>}�ο�CQ�,r�"au<Ԍ�rPUuo����_�wV�#�8�,�?�%�ֿ�mh��x_�@�>���ei�$�V��MjO���^ԠM7.9��3}�t���u�ho�!|ѡ��"��g��p*)�K�Ma���}����"Ϧ���5$��z94�E��M��ʝ:�~0���$m\��^�,Q0�}���G�B����3�'����rB��V�����V�3d�:�W����19�B�2åg!EG ��#���
�N3y�ic�;�)�Y�漙�Tf��,�dn���P�=����b[�S�r�)3QN�s���gW���d6m�a��n�Q2�ͩ�,��U�/��j;�~����� �ҙ�3��"h=t"	~r�\��j�?aY�ZYbB_�ْ*� �gJ���`,��ⶄC&�kt��1���;��8�#�!5������n�-��Cݲ�a�]䬲�[�Y�rP��ԅ�¡�G�����������N1R�
9]n..go�y5�~�ght���PT��*Y bJ=��ޡ;t=����a��e�
��ƭa=5w��t�nϖ��>x��I�&O���_E
���npu�qP���8^���n~h�ew��A�WmB�fGò��aC7����H�y\��wAge+��t1���"X�~�?�c�$t�`P�M'Xv�Լ�|�sC�l�V�	��[g��Q��#��ق��A=�_;ד_�2P�0I�? �u�d:�3 @њWw�.7e�t_V5����}�r�荐<�(��𧦇�J9��6�J�,�V�w�,̂۫"����/Pz��U�$Ë��j\-~�T��)�f�����X�	h�����+@AU����#L�=ȟY�d�d�)�Vo~���y!�H""����lS��K{�T�b�>�/� �rjP�i^�X��w�O��:#f�39[�9��2s:�.zb���!ǁ�]p����s0P$��0��P�qK׍*r���Q(�º���t���o�Y�.�ڿZss�v��ʋ?��VG�>����F�,=��a�ӧ����Sn��j5&_n�����l������QB%�i�Cĸ��ضE��v:_��x��3��7��v?���c���4�۹��J	�+)[g����o�.f>� ��m�v�s
��J�{����&}-1�+YY�y
�'�(;�4��B	9��,��B�ύ�9,7��J�8I���̍C]2��g{[ogd�=��O�n���Zݷ��0(�z����h��}���ߐ��m�v3J�iûf̑�z�S(ӰD�u�O� (j\樄PSO����,�i�Ҩ�y�=�_[���ãͰ=�q�<����6�ӳ��q#/
%�j�l	7�
Z9d��:bV�Զi	;���zL7d�&��<��L���Ӑ�wL�VX��k?��zcb��L��BUu������d�_�T��FB���.�V8.�
�XX���=|I-���M��-juW�Uo'F���`�J�֍��Pc�׊=G��O�v���A6Uob�E�^��mA��+'	3✊a��i�D%�]�p`]�35<��P�!�>aME䥮��PTj��Gf�j�L�Z%=�r��#�H�C􅢊=������!���g<Mw���4R=��*��c�h��M�uc)QZ��+0>��].��HK���G��]���D-�R1�V��I���oE�� ؤ9� �F�|�wsĠ���k���{�����y������J��\�ʼ��_Vr�
��k���2{�R��������ϔJb�k�x�:���E@nxo~D(bQ(P����ጪi���+���J�7�]&�VO�'I��0}�t�(*d!+���cc��f�)J䗞�\��0����+^L��j_��VIF%/����:r��಺Ru�� ��%:)����T��>~P%��ẇN�/"}�J�F��$F/��CXE~��q��{;��>�ל��*Tdr+��� �p�G�����b�H�ް���N+��<O���G~���Ɂ���ʙU㦾z6T@�UY �R�'�uGe��yW�5��p�۔i�#�W]2U�0�*8�!$Ji�?���]�pKZL>Ws�1!�5�[�8���c�H���|á�Uo @׮Z���x�{C��C�
�BڷAz���e��kxZ��(=ؘ����D �S���[�'��JMUX�+VJ?g�C���@B����Sp��;HYs�8���(b���Y���Uy�k�G�|J��b�vO w�� ���mP^�� ���3ސ�8NK�1�D�Qs����XGm�G�l��ڌH*)K�*��,?�٭�7���S�A:�7���*W@\�'U��#:vF<���Oח��)�M�.���D��� L;�-��(8�s��g5�7/��/��5�/̿���o0�@WY?b�vA(�`;#u_�I�Y`���_x��j0��f="jĀ�ˊk�h6��z�e������_(�4m�v&�L�>�h�k�}��F�.���{���O�ޕjf����ĸ�b���r����x�z�OO���c�L[�}�j���N�����e�\�;����Rtr4K�7��]VkK]�N�t�t���+�ZY�C+TC���V����xs�~�H�>�wp!z61Ǫ3����J' #�BTTb�p�\~�q~�+�5�,�4��Ax?�5�| 	B�Ħ偘���DY�χ)7M&�[�d�l�p�=D�>���E-�a����C+�h�|X���+֧uUe7�Q�Ohըfc�5nI�nSv�aA��4t�x�"S֊M"@��$w�fZ=���F'��#���G�M�O�0�1�����	1S>�Øpi���ƫ
���E���]���YP?�ExF�W�-�G�8���\f7vZS�A�o���8�K��Ne���ޡ�)��>�*�ٟH�8l�a$t�f��!0J��I���'��v��L�B��%�x=%$�c���Y��l]+X�����t���t���8�/`C��6��(�ؔ�]Y���8��ƫ7�����'�0�]���|>�è�^�{`�-hd���Уf�w)�r�E����ąZ)"�1�omx�ƌ���3_�r�ѭ3��&��˩���ý��l(_4�����>�ja"j@�O���W���ƾ5�g����~�0|k�1DA����P���� �j�bT48
&6����$H���w�+� e+wq^�P�����
rĳ����dF؈�/s?t�rA�'niof��K�L@_����a���S�pؔ��0���r���W�J����'��nK�U���3��@�8<%S|U��a˲�p
�5�"|� ����$��i
vI�"��"Qeث��NY+^5��Ș=B�/�����-K�(��ǜ	eK�$ӷ��To2�3���p!��Z���p�i�>�-�F��Ĭ��Cj�6�M�rSOEb'�VUs��e���6�ԓ�*}Eľ"���0w��.�IF���l�(�p ���2A���8si�Q"���1h��5N��<�	��B���ƂA�5A4��훤w�C��I3�L oe��� ��V���!P݌LQ� ��6$�;��yZ},� �&9pi(>1�]+�hN'��$��F19,�CEj�B壟8X�Z(���*{�8�=~�m�b�6��ǅC�h� ����V�E�����e���^����$(+=�R뻓~�M�g�^�;��	�L�%wq�X]��ދ$�Y��}��4ĴuI1W����c	�����:)�	V��	���p���|�2�+���,�CaE�5m�:\��� 1Xsa���o�w~L�´3о�<�b��!�nH�I��oPE��I�t8(%y���[v	���v�
.�ϧկ�{�����!��t��r	������2��"r�S(կI�����Ηݛ	�a&���
 �wLVco���p7i���Sy�g���u��?�8�7�gP�AU��+�(fP��<a��䃩.���O|h`���J?y �1�0eB�]M���>��X���B?ݳ��Y�k!O�&����ke*�]�t��ցV�ÁD�����:N$�F؉Md�-��D.��Z{��T��EKӚO�\Pq�w�?���KS��nw6��S�3!,c�z.��ڗ��AF����R=ڰ@��@>��@�\ס�I����H��T�E2'�{>}�$F�n�S�hpd�#|Q��Pt�aG��]��~�Ԃ�x���B�6L�C�譈TMw��3OA����|r��`16_�&���u�2^�V�S�#�$��bU�@M�Z<3�0/|#�z���%������vE�gA�Oᖦ=�T�]a��'�n-.Q�[Z�6u/�ɲ���v���t���~�)q�P~�LV)���B�p��Ы9��D�̹�'ւ��y�3�W�p�(���� �e��~�P(�.��F�����{V9@<9��K�*mx��$4f��T�#E�[idN1�AcԜY55g/�2���h�j��!t��b�K�<]q `���\���sF"���]�lR��j��Ԋ���ޔ �ƑK �:���<�JFf<�X��G$̰Z1�W`?�ލ����bn7CkL�-��
���$��?=
ж����T���x����#8������F�Mw�OG�`��$��bzwߛŊ��,�H�Bz.Bl~u�^���j�s�r/��ыD���oS���5�zY�)�����N����E����	��w��������<|�sH@����z��8c2ĄH[A(K�
�ΖE�e0e��k~X�}��(�6����0d�w%�W\��x��\�H��xB�nr��)��؃����R��x_�uʏ6_8]=<�ªX���u���G�WMk8pzpW1p����~:�2��y��Ѐ��H��C��U1�]��3���t�Oͦ��(�+DG����uv�.}��U�9�:�v�9b�������a�U�v~�O�ag��K~�zA^�ZL�}�QHVnie�@������^���8$a�k�7�Z�pV�i�#hK��I�ME����1[���w���fQaq��l-�����7����4l�lʯ��:���!ߏ����Ox��(X�\����ck]�òy�
�,@������0q�aS<p��lO����x[3D�䨐����i��& T1xg��I�X�HMT� ��b@H��Af�ˉ���$A�x�eY�HQߺ��m��s�w��2���{ګ�b�-��K����b�M��Gl��>�_���63����y���,�8��Dox��Q�vq�7�C�1Y��3o���X$ė����]*��q@v�l�)n�t��(ԙ��`��3v���P cJ2������Q=���ϗ�%䪹��5�l�}g��dLߨq��p=� U���gn�u�ү7���ڱ+,%�+�(��]�����l߭<2E����o�=�>D4;�62<.ho��d���	��Ε�7 fz�̽Wd�"�g�{�ո��f$N͝ͿDl��rG��]H�Y ;w�l��&�E��W%��,߷��<������O>6K:_����X���$����N1��tW'�P�����FȜ����\��������T-͡���"#��?��+�Y?'LA�`>!+e�+O��3xYs����c&�0{��"x�U�M�x��q�t���'nR 0�$��(�rxDz$�8�1L��`���e�m��2`w�A^�p�>;�p G�E22�韼F��S�*Noϭ,��tGN���=sl]�����i�\�0> WJ5�'ɬ&���m�:٤�.(z�9Rڊ�	��Z�Nu�AY�~�a�l�����G���D׫`���ǎ���D`�/E�Z�Qe�=�H�v���*MG��L/ˏ���QW@F���0XJր�x���C�. -�����CV���sΞ^�ܳ,���}��(a�����K?9���1e��hk7�~���Y��;b
Ģc!ΗR��9�~��
H�����į�\�G� �(/��
M�����fG�6=,Z�G�z��>�� k�h��=#�Gzү�с;�h�c�>�l٣�Ec 'E!o�"�R�V�s��
�l&��b<�	ݒ�vUKl�њ��#C<c��#��X�yj6�������ÁhXu�TQ4��q�9j�h):�k������t:���_j
�%Ұ6<1�ȡI�;*�`�+>R������[±; �g�X; ��dĮN�]����2����TηދD�hJ ,����[9�"�7��Ā����u�+��+;>S�Y�?���g��N�V�r�8	㹷��I$ʻ���j���%��fnS8d�SR�tboAe��!"��TN��Q��!t�� 1���/���}�p!/��,L���N� ߠ8�w�G�wD����iۨ0Ǯ�"�$��zWd �xzZ/�J
�<_����-Yx�+��+�L������.	.}��{����z���%��IC�N
�@O�f&��6������-����(P�:�$��ka��Z��3��֨�C�Qz�KA�q�,R�a�Q��֟LP��PVr7 #K�N��N1�*Rs���I&j���rbJ�d<�F �L��D87b��H���x�RZ�O��V�)�%��~�F�Pj:*�pO-/�H�Q�a��.�����͋\R6)��k��u��JF��O�߫-��'|�+�q���Ø���X�o�x�n�\ΊK������˪��.�g�'��`��쫃�炋i�Aι&�M`X�(<q��{;�A�8Q'�d��n�Q��T�p��YY���v B��9�5�Qw���C��;{�x�_�Z�� ��<����Q��YD�/{����P��� �� #�Ep�ϼ��j�i�Ƞ�0��|8tܲ+"��ʹ�n��>���V�PgQ�e��y}�DB'����Qu���OT6y����D�_y�|��[�m�T|O�~���2
�w����N�:�%������U��d S�u�&
���x�8�fF�Yt.�ii%&D�@�ר�+W-Bo����C�Ǣg�O\����p�� j��wh��Ƃl�3#@{��>���Wݥ>-JE���e�LL��LOTn����YL�g�l�*��N��bs)�)�J��X8%�W~&=��J�8�$�Kw�yL�ИO�o�m��=��5��ayF����U�����[~���̾\�X�$D&���b�'�c85�� xnh�'�'��ˤ�Ђe�Tp��l��`�߮��c#d>	k�������J'��5&H[+튎�Q�z�)�DՓ�*]*���JfRAX��Pc"�Αl��?N;]�qm�!s����I)��/�P�2G���������F	s�<�,e;6�E�xv���6y�*����yB��%��u�37����=b�mJ�o��x���3z��ϐ/��qd��x�!���V���CqǏ�n�2Pd����S���aU:"��tE��]1(١`�-[�����0NHr� ���X���5Pio�l@�)f�o�����/��§��,~4x�@�RuΩ�~�NO����4��ye����c����\�$l��~Wc����4f0ⶨ
TI��3'&�f�������[����$|�g�I���iїÔg`G�D�Ͼ"�0�|�Q�K�"��$�X?���_j�Ȥ�t��@��Z�蜡 �:�!U����]��z�z&�@c�k��K�/(#o���� {?��h�>��N�T���a�.R��!���u@�vu�b9�=h��07�D��[�Kh-�\�pq4�Ɖ����>9��G�YA��Æ1*�p���Ӧ�!ɛ�vJi�f'�U.�����'(\&���W�n&m�?�o����d*��3�ӵ��	q�������`4�Y����c�({d��B�X}��Gr'R�Ntgl�n�eB㊛��u>+�o'I�D!�Pi��+�!XB4�4�/y��F)�GN�ϳva7�D��@���z1m}�[B�xI�d��&j?�U�K��p�-`h�K�P��4���4�r�2/.7J�,�ʰH*��ȿ�,W����5�Z|2�><��~^%o�g�?f�N���_�����>�������G���3ǺKpv��e,�h衐RNv) �9�gx�(���R�Z_n�I�ȟ�6� w����W2e�ܔ���oCS�F����ar���!@;q謤�7�S�LU�,�ю�i�j�h;��j;�䁸*�[8�@���ڲ!��Z���~zmӶ)L7�Ɲ~����W\�]}S(�v�b�E��s�3S!`]4�=G�c�p��L�E �ԬP��h�rτ� yt6��ks;��v�E�b�(j"UjWBck�Pe?�?)R6��ʭ+����y��l�{���x����_���F�2��L5��z�1��u� ��c���ϨǱ��,�����:|����w�3R\!�
xQTF(�Pbj|f������S%��h9�yήM�9��oc2��� ]��*����y��.+�,�T!��dw�49�����S�����5���ɯ~�ٱO���Q`H �}�K�#c�pa�Q��8�h�6	�}��Q��a ��������#7ѶQ�Ω��HU{���.!���1�4c�3Hk����uQ��ڻ�]e�&z�-}���:�5���ʏCL�Q�
[i�$��D�N�@KN���\�F�r"SS�Q�uA��Õ h���� �-)��Ԁ˪o55��f�jSt vS'�lb�W�7i�g��iM�	����}vL�B{�~Z���i(�q^,�CbNu� =Opy)�~���fu�>�[�d��H������6�0G��[���<����O��}
����cj��n��n�g�\x�/��\hz<9+K��hO��^i+��˖5�}~����;-h�H�������Y�C��y��κ6�����
��_^�%m��>�3�����M�d���'�0R�]˩ꗍ��?%8K��qq����ʰy�.}fYIx\�y|�\���ozB����F%��l8�=O	�
��Qͽ?���qx�L�_:��<SX��	\�½�\rW�M�4� s:��X�UA�'�����JM�:燈��P^�*]Q��sR�N������C�m☠�Dw�sPr8�vsy�ww��Tz9e��(����I���qkؠ�{N�Kp����Ћ�޸ކ�k�~���i��T���.��%���9��q�+3�_^/�#D�P6��^����������#Ζ�HŚ0��#�VuaLJ�?�B�GI������\ŤM%�qQ��3`�gQ��!�Bd!��oԽ�av�#aܭ}7�_4P+ @/f��Lw4"<�|날�qۆ������������3!'��j��h��Z;��.��
�����5R�s��ʘS�d9�6Q�|}; K�%�g�~�7�-��T9�:�Oz���xO� em_Qj�|K��_weXS����0�hc��Ƣ!GX�B�`��x���R�V�8�w������lqm2�+x�b��-I�,�|q.� ��wٛ��3�vX�Q��yVY�_��@�Ʈ%;�fZ���Yy�;	J�c�ݒB�Z�y�w@�'����*��,؀HkE��:��I��I�r���hB^&on������0���B,��l0�v�S,9<G�aT ���������6[����@����n��vg�@b�rp��G��K�2���+ r��S�<d W�0���E�Zt}����5��'��5"t�fD�=ܧ��NuT���_ @a)���7(~%`��0�o0�h�F���X��6�F�e�8�O/��O�&���?ג�,޳G]�����g�H���c֖��sZm�d�4Zq5�X�5Í�[�Q1J��&_;��6Q�psX�u���R9zV�*C�O).@���� ���ǹ��2����v���蟊
��8T� >++����zg��@9y\��6��`��a�����%3�yh@d��6G��\�$;8��V�s��N��?8����q��»i�@34̼}�)O�Uu�u��H����UyH ��`�k��`P�Z�%���Ɇ�x�SS)5���<7tr�<?i�2n��O���A��ʵ�i�����H�ZD��:�� ��p�k�~��'��\y�9,ɛ�*�G�dh��j�J�I��w?hSQg�	���ɓPCgZ|���F�d�)E�l�a*��/�mZ�%L�D�
t�{�|��h$�*U$��1�|�1g�t��4��O��mր�QdKZc�����P}q�����e�SYXF�#B�P\�����$z�@��+^$��{jUv��n��\�� ҂�#?��>��5�.ތ>�SLI�Q��D������I@���028R"�l�!\�ڠ������5(o�����Å�*6*OO�b	�D�5b�Q~�ם�b923\�Ft{n삒�����l�A,h�b����6�h�_�1���D͖~��V�G\3�k�4�:V=)u�~+�����J�p���V�É�D3x|O{q�eh�c���;1%K�G0`ʇ����)y*��Y�jS#��6ұ� [.�J䃲$��Q�4��S�MϦ��nu�}��]�� 5O/�h���)L��mu(�hvɮ�$	�V������P��
�H��������N�������W��!���_���ɑ5�*?�����Fe�#W;��ҵ�����h��R)��;/���z�Oph
-�ȖIm��rq�c5\l���9��P�n�m��x�o��T��dʒs[�����4�ؔ��k��M� ��Ӽ���s��I"��t��:��$����m���'�y��R������}T�?vU{AsD�^�1AJ�A��)z�t澌g@qu
xr����^���d̒��A�I��P��C�C�t49x?�5���IՊ4JD�CPA7���_j�(��(cBH���g����6�(��OɽPϼ�BC��uak�������1���	�YVTr	!l�33��:+�ɤ@�So�(�~�{��p�Y*�4�s�!"�\��<�a�"@���"؇>'��<:͔�ź�o��:ͭYL�9JG��N��4�B߾!�u��#�+3 B|	�1��ʸ�w��R�S="���y|��C�e���Nx�k��A`΁����(Mڱ�^��}i{����D�P���B3��m���D���"�Z��~��*��ah))s��1a�u��/"!/�����)��qjs�_C3�}�@so��/y[aIc��ᮋ��iW��ԛ#°�ۃ�G���޴�^��`�/����.T$��
�aA���g=T���h�%O���U�Z�Rc`Eu
NB�$񼁞�`s삐���O���L����9�#��u��D��8�G�C p�묋V79�F�Ś��W�x2��w�[��S��;0�W졫zq BE�0���f� �����;z2���T�~�*�"q�4�&�.캟Z�"i�On���]��#�:J���n)��槽Rm(�����	������7��D�]WZOT-ߑy���±��P�)�(GY޶z�w�7+� ��N�U�g3^��l:/lܮ0t�ƪ&��?��1A-CI��m�ABjGmM�q"�e����Q�6��Uh{F�]D��J����9��]�| ĸ��c�D�呌;�-c�f���u�f'��3���f�wV����XI��"��%Lâ��nF�u[��/���i�Z!H��\�t@��i���9���*Z�����Ԁ�/ �=�G?��h��~�G�>���*6eo~g��С�Nd�`��mV�s�处�=,30�S�)`��./h�v��N*zcWC�kC<�T'��0 Z�6���3Z|��I��� R�ď���[��[���a��u�^�g��[�8����O���2ܮ��7 ��~%�{�|T�*�k���c<����!t����hԃ|�.�m��+� ����֢�y6� ���IL��8�V�N��1�k|h8c�Ɍ[�s若�f���]ZWd�Lm�{��s9ԁ*W���# ��aht�B��~cL���v���m�BD��ehi�=_R���UZ���H�0���.E��E'?4��U[�Vr�([la-1
r8qF^?�G��:�����S�L��{�8�q�fs�d�hAЛ (t_%��AIt}ڹ[ ��joN�c�v�д�C�40.Ǔ�MHy����L��4���t7�O_�˫��Y�8�y�F����9�p1S�	��L��Ϊ�
[}2�[JZ�5���A\��F\�9`�L@.V�܆�����̺6>$aM�L��QE[�&%�n���4o!�z��N G�����pX�e�H{���Vn��[���-\/Y/��K��e.�9�������֢d�s�!�U!����Ue��g���j�����0>���!w����yz$TH7����#����ҋ[��ё(�Nw��T�z������?��4�����oJY��t�j�,��M�)�yJ�$����w��ˆJ��^�L�E8ԟm�bS��b��#'�Bh�B ��te�`kWq��X�:��Q�����L;��������~�)ac4����#b��g��<.>�Lx�����{܃|U�a����K�3|+D��� L/��Y{��zX���< �-����ex<i�c�B҉���n�֟gNO����'y��y����Z.�O�߳��~l�{���񓪸$�t���'��W�-���]�V�J�=6�)�~��L�Ѐ��n��|����Zs��.ɖX��^���t0]r���@n���;�ܠ�� y^A�*��g�T.����~(nnƞ�'@�q;�[��I���X��'�Q*����ik\`A�Q|
����GV�"���DD��q)� ��e��h��[�0N�� �;�E`]�C����p�e3��Vϛ��;�c�,5[W@���?f�:p4���J��#�ՍK�!T�(0�m�G�z
��y`��"ɵi�H	3,k��!ē0-I���c���kbxx����"Eo$g��ӿ����í�>�+��海�4��L9��H��@�Y�,�����Җ�p�ݸ�p�X�E2P߆I9F�o"E�XCKo`�u��wH7 ���F1H�y2�/n�ؓSEn���ff�x\Η�cO�B<�b��	/8�9��J�&�F��̛�%I�,e�M*Axg�`�:�EZ( 2 �g�k�v����je��������k؏aVR���b[C�;I4�uM�jB�g����2S�_��\�-�N�o�v��rf�72��9=��5ܖLYW�[�9<��ϟ���fc�I���L��b���T�V	��"��'��蘠 �sD:�j����ӣۧ���9�R�ր���(VO3���;33e�mt�������M+jY��� G���=�9A�$���=_�AΑ+>������bC��>����a�o�:�0i��J�+��Ki����;���Gڈ���WS��wR*$6jB � ����&�ȕ`K]"^X�Y�5ʫ�uA��lE�n�M.�,]��W�DS�X�I�g3-���%�3��t�����`#��0�w^�ŗ��/9��;a?�O*��d�`]0�JUM70�1
p���[ ,�`AX\L�h�b�2�ٱ�Vq7}� �<����?��Q�Kml���D�W9`ܟ��+t���i�4T�� 7�	�`�u��(B]�Ȗ�F�i�u)f�����t/�d*&�x�i����,�O�3?I�iq��U�?3���,w�;�t�	��Q�;��tx��a(�>݆g3L�I�%���e��vR^Y3L��`�$]��٪wɝ0ڤ][�W�M�vMgũ��|��[���[k�(2�x���2�+�"�) 8��?2�LHc���`�U0.K�"7���Cn���EC&�t�������ŗb1��]m�B9� x�6��2P7K���@d�)�>zޫ @/KW������c��X-�毐�D��7�$;���4*�2��)�������^��hZ�i�����^�!�bף$5rt6]!@��C�%$d�y��?��;�s('@��E2�z�t>!���1�ə�/������4�����$>������ߨ͆�f$u=�a���_���Y�޳�ǯZR�A����o�#QM=�m4��VlY:�]^+i|:�h����N#�Lg��@�/��'��ta�D����f~pK�{��j�����*����Fdr�-?���H�3���Ŝ9x�����2֝+5p�`��]1�����MAt層�F҇^_����7��ԧ�$A���0j�A��cY�z�_����4�\0�&��CF���������Z!9��C�������;[�q���6[��9�x�o\�/R3�G�g9�+k7�A�"j���:�������n�hd��c	�[?�Ps��,�2@^nU��f�B=��
ƀ"�����I�8�O�x�th�}����5yu��p�uM�5.�.��v-q�8��-�if���~�VӴkD=>�^�Z��R)���Sp���CK|q�+����t��P� ���z���y��	�~��z��f�c���M��_r!��S�lS�m���<7��M�[\���}.�;x4���&Ě���Yq�,�:П<S��r��7�H�� ��]"�<��c�����C��.���:��g'�`
a=� �E�$����E^Y�y���̱�bIe�fG�)O\��7
4)���ʛ��ҿ�8��s�d�G5EU������v�-��#Z��ǙO
c���+��'BqC��8A���#㸬�	�_��|��*n��X;�� wŜ���>�&P8B)�Р�<;�X�#ձtCV6-�����x�<����m���^q���[��KvC��`���DE�RfI���ɖ��G&�J}��K/�!���s�kgbh�ϰ��%KV�M�%K0К�}�pY>@̝�0�� ��w/�9����.*yF*Xk�+T�k����!$�dg�����ӵ+�բ6���!Ln���~{7�+%�2fc����k��w��fP�S���d�ם�PD�2AI(=/���	-�Y���ѷ?D�?}9Z o�Ń��ū�q+w�� П�\��2�F\��� ��*^f>��"VN�41`��Ftl���-&ꚳ��%
��F�1B����T$��'�N,&��h�M��3<f�Xp����9��R�LK�x����@[=vqo6^� �!�H|x�L�,"q�� ���<�t�3C�*��2b�T�	�)�;iT�g��ڼ�{~��=����� 1�����8,�O�\CS�fx�ಝ-׺P�9I�̢m.��鰯n��s�}}h�eh�bU���Lg\�V������+�&��%)U�'�:�w�g�i�Ĩ U-l��	8I����"!�0�5Z�d�:�g�E�\�	��3�a:	v��r-g�@�8Ǿ%�ڰ^OL��'��/�`qc�R*$�(�9}��(1���^v
���*}+�0�;;�����	�c�v���E��
p���5ƆUa@c_qʶ��^Ċ�"����;�)�y���C��@�v�y�<�nE)Sz��T\�u�z��aocH�9��V���-*p<�ICA��� ��?b�$��&Pg�ᜨ�d7d+̞U�Ƀ�X/$Z�m|ɮ��Y���0�`̽�i)�>4  ���f��w�����3w^ی͜�9�ɀ���D�p��_m=��R?7�1E���Mu��ݕ#0/��#��C�Xk��[��\
���c�75�+�yWvhEI�]p>������ꑟA?�#U�����T�J�id�0������@c��(��i��S�5��PS�QT��d�^m��"`ZUFgA ��P�D�]���B�*�y��#��=���n�e'�eĳ1iY�L��i�(�w�k�]Jۏ�e�8����C�M��hf�)o_�29��dR�����.�
;�Dx*<�<&�|���m�\=�Ñ=�5	��#���&�ΗlG�&RJm���DlVj_@.�~�ʃ4Cj z���h�JCZ��؄,�������#k�o�_���a(F��tg!%=A#/$k�~���6��+_����6(;s����^��Yكy�T���{-�4�3XU�L#9�, s_�[v����M�L��;vW�0�C�YW-\t]�{؞W��=rw�}Ƃ[�Uq�c�{�/�(�o��?��۸��a�l��$*7��oX�|!���]��<�$n���~�I��� ��&Ha��M�g
�E@�^N�Is��}���R�����K�H~�?�d�ِ90�t�n�Ț�*O�[yv��Pgc�n����Dj'lǘ eHc:\���\�ݢ�@Z;X��@�Q]D{W�bۮ���E��벌J�?|3R��/�NgG�[w��H����`__�iI�4��Z�M`3���z�{^7>%aY���	��B���U(�.��j�,3�Ԅ���f�?s�ӧ,�&� ��.�0�⛌�W�FC�w⪙H�@d��0ǐ�R��:�Ô��NZ�����0�d��z���������Xm̫�F�R�ǋ{؂��d\r�R�6�(�1;^�z������,&�U�C�3�ь�?��#e:�����V�Ę�w���0�y�N}`i�C,��q�����y@Հ+)�[�l�� n��[�/p��O��4�C�[�lw槚��
��;���7S�1"���	��Ϣ9���ի�f�n�;"��H?c�I���u���5�K~ۇ��.j
��i4��XT$un�J&�v������X�&y���<�|m%��H�oMB4KuY;M�f��+'�_���4t?�5R�C���l�l����`��1�X{�nN�n�dd�{����LvƁL�;|V�'U^��A�s?a9��S�`�9�<lT��w��X�vDO)���n�g|uH{���Pb�#��ar��u]hX&�$b�yN~v�������=����#xEzgZ�W���q�|I��	��/ͦ̒�ᐲ�m���ŭoU�������o����8w�R �L�NE)��]�a,���E�ߟ<|_���ơ�Lr� ��e \��5�����$�N�-��lI��Z����D���6d�M��b�5W����!�4�Cj�6��Y�ה}��ڮ�2�zG�e�w�>h�8I�R��ގp��7fE{�	�@޲y���
�o�-�I3�:��u�H�fF���_�S��{���ñ NK�3�9�'ɲ&��MHT�jo�<�5VCo�B]7fy^T|�;@t&�$�.��I���j�_��ਚ'fIQ���Om�8=�È��XJABx����C�M-j�����FC�>�'4����ǥ�-O��%��J�-�.����Gbs����$�:H�f�xuhݯǆ�Jn��՝Ԃ	�@x����D3�_�ʂ�"���ʉ*�,D�N/0Pup�։�Ue���!s��oH���F�t[� x�&���a�w�l���:\yB���Y��:�����é{��[MKk/n��r+��ƾK���9�fJ8�)mDLWo���h����9�.��|B���'S2��blGv,3���*���j����"[Hs��^����}n@��íuԃbpxF�����Q�4��V@�q�؝�_ZVLm�z�i��}���;	�G; �=4@ `��<���$+E��Lo�N�^�8sC�����z�o�G嶸 ��^ee��V1	�E2� �U�4��H���e*Y��gꕸs������΀x��#R�>=�=���SM��0���*~8K�Ji��dYWxӇN���?8`__����TQ�^�Jh�0��r����ċ����G�<��:��N�֮[v�&0��9����P��W<,�5W!�7�ɤ����Ί`�5Y�������
O��]�R����%$�dRȵ��>�)���8�^ ���E���o���%��-=�F(#�6lV��7���],��|Zl:�(2�6�����0�;s̴�1�S�(M��?e�ֈ} $��|Iڎ4X�������[G�0/�y�o�Y�a��t{��{⵶�����6^ݟ�>��d9�;ӟ�=[�
!s��ф�~�%1	��i�ԢS���v]]�Ƨť��Ð?¬�oJ��}ܧ	;6~e�MZX
����h��z璏�-�6O�lV5k�`R�̓��1Õ�Sv�*�xy��T^���8=�h?'R��:��H�$\�](rn�S;\1�↞_1^ԩ~�r�h0S��#�L�c㝫�mǫé�jb c.<�R��m(��k2�yi}]�,C��b~��%c�z��&��|Ĵ����`̃�!y\��\"PY9V��qY\M�޲�k�R}x<�	)���<�zl��>΀��ao��q�F���'%���)���0g1�_k�)6�C���E'�<^^�"r@�U�?�c�B��Dha�ۙS_��hs�5��b��L��#�E�q ��S� $�b)T� ��c�.�*��AB��g;���v޺��)�2(�Em�i�˓N?#��Yn��M[�䦷��Dh���i�͵/�it4��iOx�	��\�5�a�f����U?�����s��"PGΆx�t�T~�������Q���>�B&�R;���HK�-y�1<���Sܫ°W�-�^:�s�Qs^��՚�Om��A�77D�sB�R��4��UX�"������m�W�if�Iڡ�w��MN���c<��p��я2k�R��<A}��I�"6?s3�^���U�~3��,���!)�E�ܠb]d�3i6�1��������wA���o��R�#�xs`��ҩ!��U[�T��G������h�:��0;j�ؼ���-r9�=���^'�]�?8χ�(��A6`E���p��OO�$>|���)n�҉�Ny˚��s�5OO;弐{�j�f|P��8��[�2ht�CJ���l�/E��8k�@�n��^���or;��ia18�*��U򰀡�,�*4�PX��R
`f�h���&��O3Z#�T����W�#����(���i6`����ަ���Uë�dG��0����g�L���,b���WG'v���"Ȟ�y��/���$q� ��g8���l��l̤�N�QP���ԯ��nK�Quw�屰�8���;^C�5�hu ����U��D�P�Z`&�1��4�a�kZ������{!4�&�M��k71�õK�VG=�=f�����R�	F7�DrG�U�`�M �{X�Yۛ	@�f0b��0�CumP���?H�o��A�~���"�)0R�A��i�E����ӡ�)����C�����F��T۾"�O�cLMt�<����p�(i��N�,c�K)6bEԻ?
���M!���6)?�%��QH��8�_�H�D���zr�יS�z6�I]�?k^>�f�\G�>i%\��bM��\犛�kX����sD^{L%�SR�]��#�|�@�:�̬K"숈���y H���}Б�x9,��|���(} �����|�� +�ؙ-W@�n�aj֙��qNS*1K�=p
 `�6d���:]�tu�44jIc^Cdl��r��k�OB��:���,b�m��7��>�k0�c��IKV�&�(w��*йՒ^b�&-1+�ӌ���i�_��WźY%��짮>�� @Yo"|����S}�1�A]f^�fr�'�Q�8�[�#��Q�3.�˼��!$�`� =��u�l���b�Q�X�%FSS��R�S�����78�Y�cgISI�d��BB�O�0�� ]E��?��,��1�{FT�^/󁣛u褐	SI��ds�Th�yi?Cs�.P�����'��M�[�(���nl��=1-&��:	{5��N��O�Je���+�o��#��;;��ۿ��HIsұ����9u�T�5Ȍ#���?sF�����[�9b�1	��d*�Z�F��n#Q���2 PεTj�g4hX���
jaR�(t���{�+�h�ҪcPZ���%���++�!9��X}8��y��99>pq��'ψ��+Z��97���E���fE_i2ڜ�����3a�Ƥ5����ݎ���obV�g�P�k��W��˸�� l����,M�đws	Oʬ��f�YYc��5���{��\f�C������Xρ}{��x�	:l�~謁�	��y��2�{���J�!�x�{�2?ҞY� ��#Rd�GP�����:������:v�u��f�/�֕���N����u�B#�9mz�;��6��`)�F�[�f�����ՔT[S��R��m��m�q9t�e��I����ֳp�����c����+R�U����|8����1)���Jh7P�� s;W�ؑ0��MZ
�(��DXF������'�Ɯ�z9J�RI�/.3n�)f$�'�w�C�e��t��z�f�}�%{�(�Io*��ˢ���������5�A��� .^33�CG[�S�I�<�C,��r"�4���Zl�#܁� ��w>�xֻ�C�YyIU�'�֥\����D~W��>K����ހ��z�1�"�R��`�[Bʻ������n8�\c�m���K9���s_@X?�SB����N�wހ]�ߞ������6�%a=�}����ש~Y4�1�_�����;8�r�ѪI��V�f����sЙ����G�ȥΣ�(����B�OĴ�*1wi�X�o))q��f����SO����>2��8�&�Ѿ��,/�&��.��d:�Fָ���.f���^h@S��7��cϚ[�]����`ظ�c�L|�.�#˪��q)�9���(���a�}�&G6�r��ba=�D��i��X��a*<�&4�>L�"�#�d�I����dY9V;Űo-}�	��C�p� JN�ם�ĲŅ
��w"��@W�ŝOT��/Z��?�d�w��<�������R��R��
�Pm��5�cH5�|�Q���Q�����C2h��� ��l������:�f���t�i������g�g��oc�rCi��M,/Z��;Z�C��.�<�#��0z��j���Bo����(u��@���¤%��NMͩ��G@��-�nh3K�̲�����~�)���[�K'�ן饭�f�����>�G�Kq�p�@��u��P4�f�jΞfE%�x�E��u��2��00|��߀�Ls�v[eB��!�*�LEs����xU Z�G[��V�i���N��k�rK����sù��:S�#}�����"˥B�����3] >+!��;��p������"lPq���F1iƑ�~���s0q���ěi���~(q5�/_[%���Gx1�K�����"��Q��'��?	0�1 �H�Z�06X��sl�ퟸ��$���qPp�ɤ�1i�/�ZMJ��+��\+���dÐ�)`��a,Jn_��!��y��d|D#�!̓��&�rvb��D��\I��C+��@%)qDH\w�ta�!���]JY�D�_JO���:��r�����Sub.^��H]����.=�.;��G��P2|R�@���j-���T��k�P��\�\pf6�t#�SèfC���1�R��j�6��.�!T���*���ŧ��E��4
�Z��h��"����j���{̀*����.���رIY�d�t�ޡ3 Oh"��p�z�C���)���CK���p���/���>��.�Zp�W� ,*Q�m!JmY�@��8���i;iF<#3_�|�
�þ��m��@�l�� ښ[s�j�I����>~/��=�I��Z� $-[4([֠��:� ���0F����FJ�4���6G��d9�۰��fc*)B�j~����W:_�ҹ����,��5����\(y�ԕ�gi�Z��姼{dB"f�-�`S��'E��b����ǙJ�6r����>הn򥚶��T�w1G�5��مt�a����ΠK�2o����������Z��@�2��
L���d~��Ŗ#���cR�"�,,m�x�γ2���e�h�����h�b�����JI��)�EpI(6�fh�N���3	(���Ã��D�Ԝ�j���Ey����
����L5)��
O�f9�5�A���"�堪o��-���d��"h;���-#�Z&�ܞg.��pLQ�2��C�I���5+�3��Jք���`�5�0Ԗ�cR0`��vLy,�GB��һ~���:`�(�9c�����~����Xb���b�"��;�T_�E�~�ZI�Q�ݥ��%��q7��=�Zc�̓�&a6�����=Z�A�	��nw���)~�I.%oPŽ��U�Q^^��is�1E���@vJ�,ܑ��7�)=����|/׊}՟ݕ�Pb����nT`��£Tu��wJ�$炆�v�%���3�V��[��;����Q�"��:�ci�5}r�Aeml�������V3Qݞ��	
H���䒞�)�����:c�;��SHB�@�q�;DF`�p��9_O\a@���N���]C�JCK��*i�T��A�[+M��U��e��	bhN�s9�^����h�G�n��Kv_�� ����Q��cj����r��dZ�Ez���j'33�,�5���_���5k`)��cE�����J��Q����Z1ʘ)�Jvz�����J3�gC��]Y�F����Y&D��>�~'P�ا�ǡ}HY�Z�I�4l!�B��`�Ѡ�M�'�79�T�B8x�U0���{��D�$��>�7G���4-q]ij|a���H�0/��"���
H���ջ D	E��m5H�c8��H)�-�g/��oA"�nhu����۵S�)X��$��c���%�Mvj�0�_�c��y`��g�-V�N%BW��䫇�S��I䘣iA��Of�0扙�s)�]'	�0:3V�h@��ZXh�������J}�	Nhn[��{�ͱ�
k(*e��D��hA��i��n_Wϗ����>B��#�4cF�H��ꁷ=5��Tb�~�ᏂS��M��ʡxD��Q���#��&��9p��?���Gד�U��*�݄��z�@�"g޿��+�`��7~�z��$Xx����w*�ŝ��kIC�Q�U�I��8/'$����욛�����D�u��-U���u���t}DfS	�.]�j�Ā�w"�Ԃ�g��ٴq������.��Z
���k��~5�H�IZ������o>��
%^�?$M
���� �?et�\A-���ꜛ?�S<,[y�����1��k1��I�o|��T�(3::5�R���^<h���,B���T5 �o�Eߺ`��L��Üv_U�ˡJ@�H[<�}-&g^mbZ�� �e:!d�9�es{+��R%�lA���h�;� ��㶶o�y�t���v.�Xk�m���g{���%�Kz�8�n����a��lx
>6t��{�|71�eLx�å+݋�J(�>�_ff��		�{�zr����;p�
��j�S�Z:I}�R�ܤ*�ZR�b�#�,��x��8��̓��Kǵ o�]�t�I�P��C$�%|��`��i���x�]�M@�`6PU	aׂq�ܰ^V����m���w`捻EQx�����X�fa��[;���`o<����K���mt����ǃ�5�("�@V�B&呗*U�J��	�e��/s�5~!s�u�QyA�r����s��#�cu���/T�S#p����ե6ʝ�`h>��-FujgÑ�~'�^;����{� ��26�!�?^�\���YD�~�R���\_j�DFD�-�՗�5�qϤ*Ȱ��޶`o�$7���K��$Tc�.�Լ�U��ؕ��F����b+�ND�\�"��dq¨����8��%��O���z�"t�ZQy�"����ђm��nT�wQ� ����"��\���_H�>b��\:* ����h*o�{���������+�a(��[oL+�R8'�nuQ����#o�����V����t�����F�t� 7l��N]`"n���H���:��U(�F�@�t�/��$ck�ž.�4��Z��#˲N`�����i#`7�B~f�@B���mB����F�Vr���@����]����>"�2�r�����bW���W��Xݺ���sی�:���&�/�����N��~�Df��� ,Wo�ߚ�Ah�A��@	ZAU��aI�)zm�w��Ya��k�ʍ��-b ��a��a�(���#2�Sc>_L�2���L�ɥ˨g��FwR���.�;H�{$�O�q�~U��{�FuC;�QH�4'R'y�2p�V���"��c������4�#��c���Y��I�Vs01[l<#�,ᗗT0�E�F��>�pV��ғ��xo]��{"{.TgL�HU��K�P"͵@��}ۙ����]�
�&�S��;��S��vКE��Ǆ��r2����E�k
3���W�8��	"�q2k��6a�IHk�Yp��wWV`��=u� �z:�f!iM����В�% �#�.��0I�v�%�H0D���_�I����H�p두��Ͻ�7�u�`u^ں��O�F�y,�o�G�α���:� '���g�sh@�2��6�!ͥ���|�[��� ��`�p��?X���KFk���^�[��M*	��\>n��9f���unp�[Gx[��[O��\�dmA�R���Z�$V�$�?Z%ؼNľ	|1�uX�Bv�&�һ��+�#��#��g<�A���R6��I�o�.ҁ�	m�Wy\s��s5��4�o��l�C7#«!���W��\iN��c�����](.c��-xӊuw^��6�Y�(	�2��d���y����Y����b�2Ȳ�:�Y�'O.Ѕ~ꠇ�NmS^�%#���S�4��p|;
$8uj��k�7��|�!-ه���?e��0�*` ȫ�/3�mЛX���"��}8K��u���>V��4y����be-�$�d*>���w����|�G��k��*Ծ�]♯ʿ�ok��_����&��VH���?�������1�VN?*p9�ny�B1��{`a	a>����>�3�MM
[d:�D1����Qe�s��%�����/�"��F�����*�$"������CZ���ǋ�fo����;�z
��]� ����n��=�h��ؠ�u���Ua��9ZQ��6���ip��vip��+�޿+��R�B�7Ȇ�3�;L[�#���zy	TV:B��3�����btS�ʋ˭���|ľ=��B �]HݻB���ᛣ�ݳ�y; u�`�x�d�r���ө��}�0 �
�~��i��U��-rQ?������o�6+��d�t@�4n��7�٩�U�֫I;*���^N�Pxhn����E���qRK�X�����d�4���3�:��=v�����G�v@�,i�R���dN�7k%	F~�͛fLp\��3q衉����|��L@�!a���>��F��F�����v}ZΔo4���4�~?0ާ�S�1k��K[��X�c���(���0eM���'���-4�l�!��	�)do�s?�;�J�d0�R��q��Pu�8*�x��+[*_&��~6}{������i{�����PS�7�~�-����i�Գ��Nۥ�׹������D:K�4Kmx��ӕ'�}կ{��m�R[.�9��<�S�ZY�o>�P�ţ��Ual
m-� ��ހ�bU����͒)c:T-��v��˚�Y�FH2�P8�N`4��#�G�#���]!~
S���[����yzB[7�9�?H�Wk�fP���e?S����̲]���9�B�Q�R��u����+�Z��
�jşt_�#�����I�ò`u���&nR��~մZc��$��뺮7_<tU1siv�Q��#���Yy�T@<v/�������K�5>O����c���}�V@,���_z�R�>�"�P�w��6������f-{N�-*5�p2Q��@� kY#$8��[~��*��. �aq��M��硚M[9PsS�Ր������+�!�9,������Ey���O �������)ļ�J�V�qJ�I�pߕ���#:��q�L����%���Z����ڲ�/?��E/|�7�g\8�ļ)-J�"�C"���������d>~n	����}���/���pt�Ku�I����S��ó n)�;���iOC�PCFW�^%��V�r�p��<�jL�p�[;IR���`(
��y�1�:��΅ ���B�$8y��,��/�^���X0�bZr��߿`0�H�����b�)&���95U(�.�ҋ��iC�.��\6�@�tYk<�h���{Mm5�g�6���B�
�H�	�����
��2�:��.[
@L1�;�aƻ�����Av�m�@����z՘	]�f�F�)u�b�a�TR����D�����N2��;�B�8'��=����S�/�� ��1^w����NHoѥ�Et�7���|�+N	�06���A7M��4 Fɂ���&<��>R�e,F ��K�c��ڹxe�����"a��]jb��Dp^0�������$��4i*ڈ4��� _l� �<���,�L���?��,N�6s��hJ
�N�h��Gexx�p�4����+�ܘ#9����/b��=���!��dF���J�Y'���.:a����7����xaM�I�|��D]�1$yZ���j[�R>v���?mY�`q���+ݑ��
�#������:�ve�)����S6���r[y>��&eI�H=2]ª��^��s��Ġ䪭�Ĝ��`��[wֲ�5'̴�Cf؁����tCC����X��3�0#�,�<�5M#��z{��Gl���#ta������d��FE�A�M ��&���:�a��-�.��И{�,�p2�1�ӱ��>6��րs�k���8��w���ͦ�6H�R�.���L��-'��.��6�I�oVaw�9�Z��E��e��g����wP��3h�¸"�u��U��-���,��b��S'��X��z���9���{Z/�mv�%sFk�����7	��e74��%KTN�he|?ڣ�E��xݗc�:���,��~E��沃�^��ꛫ�"�G�p, d�0������#!Z�2י��4T<"������t�����Y�gl�������E�D��M\8��r^�������~���I��4�n1���%�6���$e*�Į���B���Fs6苑�;�׽/)x�#O^� ?���A�]aF�ǟJ;�u�4]S���L���(��Ӎ�Z�n>�0HM�ÿ&�z�Ͷ��Ʀ q=���՗���?�(s4����wOĐ���sv��ϣr �*����~1a"��� [���6���eUK;�[m��$<���!M�jH�8�M7t�
^�=�E+ؘC&|)l��qM�#��c�.�;������X�����8$�
�G������7_G�h���vwhݿ{�6��ji["J�j���Cޜ���Kku������?��2��8����v����yb|K{����"��r(��V�|�?؏2T�PTgG��OX�y�����E��'�@F �Y�*��u$��� A�y%[�#2�m왲�����S� cp-�g�h'w^�$�C�열�ߣRx�6�������Bx�i���4b_ZS�+��$�����K�/�ڞh1�d!<�ֶf<3��'�,aVc�k*I-��R�hȣ��^JY�C��\�g�P�q�"�[{��l�Nn򴫦:)W{��@�em+���Lýl͈ A���w�#�s���Zv��*aƕ H��r��g?�vt�#�8ϐtr�կ�iI����I�偮ǡS֛�h�-�N�����ۗlC��',v�Ǎ�~.	c���$HxW��=oyCw�*���=���o���\+rty(�^gc�K� ������j�ULG�a�7��������?]��]ٔ�$2�J�C��pF
� �F,ulՃ�Z����\���z�8�j�R@�2�<��{�z�o����g�@&��Ӆ��u#@gӶ�:)�g.B�� ����.:��/aA�{!{�b�P��2��(�&�R�C`Q��g��N������f��H����/Ǵ�7�ܘ�Y����q������	��Sw�W%{5��f��a��s�x�R���{J�]�T�/7p��u��rQQ���'%P�cb,���2�_x\��mF�U�C˜y\���e�s��r��7u���KQ1 "�ܯj	#ji���,�q4[b,a4y ���jH#3O�[��٠$ͤl��)H
�+��{�׍K�n:DK�{{G�H` V��Lmi3���dϨ�ɻH� ��ֆ�m��dѪ���g}A-s̖-(�����a���䫦����,:(����|�BSS+#���JV��=�m%���Ҵb��c\�?��� ρ;��筄��%I�آH1�B>�i�U];�p[�p�Ij�����l�N)��|�+U�>\��pGA�N��^F�察���6���߹�s�1�w��vK�,�C����"�՛zI@���:.cf�����fe7:�tB���ѧgw�<�m6
�R�5-��Y~ݸ���h�8����Þ|bI]j����Y-�{VL��n���i��v`x��z�R汨�Ng����š����,y}å[;[B�E���0��s��1�Z��*58q�P���q\d'ͻk�@�:{�˴%;����c4T�]HD�{��G�p�&Aʃ�2�>�������a�W6-{:�Q]�0�����U����[��>��

����S��s��,�׏_�_�5�ns(<@�s�'g����V7W����K��Wt�ՙ:&��Wi
�E<غ�G�ۀC=w�l-]N lCW]�����9�,;�ҽ�1%�6�͊�jK��D���z��l#��~H�;Z_OΕ�rXu�f�-0l:}�a�`Ō��V��`�q9_�̊P���1Sq�xw9���#����G0����&*�-�_/!�H�:}�,c��j<��9����@��T���a�_�b�B!�Sl�z���z�����T�J�)�T�R��BMV�;���ʌ��-�l (��Z�Z��u��R��D!i�I���sOa�|�>�χ�.�wRFe�-���z�]3�Z3��2�g�ֿe�H�O�/��c�W�l9�������OO�0&�Tֶt��\��Cn����p@�/��c���I�OD����)�A_T��!�������s�����@j�AY��z���A�Aϑ�"m��Q�ph,��;+ H��}�ZV�%�s� �bPg8���2��Q'3?ѹS��7UD<����+��QŐ^��h�>��fx�o���� 	�&b"p�����/�?:&G�J8~��C�����0��{�D�Ds�nĪ2i�����˒$��͑�z��b�i��Yo(K���Z��&�tCc��q>D5c����civH�~ɚx��E3����C���~?�z�! �o��0{8�@"T��W%u��n(�7��0�Ş-�Ŵ��,��8����ZY\1�G�Nw�>�e�=E�qj��í��"1��4����5*2l%�*�wEJo$3}�B����;�HIM��pk��-�Wnq����ʯEe[ƛw�b/��=|d�<���5�:�D��l�/���;tg}�����/z��T�FOqIN1]����-x�+�>�0�m́<]ܕ1[<�.S�6���sf��i�^�G��LR�����jla w'8���g�A�8�y&L��:
�Y����_Vр��E��KN�$��7ݯs�Zy�ޥB�r{�9�i:s���y!��r�ǽ�-��%�+��{�8���~�EcPhY���|���:�� hC���Cl�[2��!�l���҄��9A׳��0j��͝�Q��Rw�JSu;�Z��Ǥ_B���q��œY̌߳��W�-�1�D���a�ۊ:yP]�e��u%bZ�ErP�X��dЃ�G��Fm�8���Xy���f����1����6�̖$'��F��l���[Bώ�������r�#x� 0��7G|h�Jn�G��f/L\�J%���;���b�b���H(wql�$\��u�`���j��w��??�c1A!!��j�� }��L�}!�Bb��:n�p���F��� �n���<X��=��bd(�6�| ����}�O��m�AP[����<Q�K���.�̺���N�[��-cd^���@��vL|�
��<+��v�Q�s����4^!]N��r,�2c�xR�'�g��q��so��j�3�0H(;���>� �u��E�P(u9�O`�*z]+��N��a5��i.����%�T��"*q���}�E��B�}�&
Uqy=<��b�T��E�'�~�!wi�)�oܳ�7G+y=��Y�Cu{�T�����Օ��۫*�舮�Q�/)��-0�ώ�A.h�k��`�8�6�I����*�ǽ����_)B
t�P�ɰ	HN�l_�>2w��e'үf��"��/���:����
J��������4��"�ِ�{j� ElW�pD<P^�-�]R�;������5'mW\A��w��e�Ȇ	��\b���,�Z��R���J�A��+��cIi^d��'��z���;p�R����N`�s^o��Aph@��s��wd�ש�M�!��k{��ݘ?�Ҁns�},y�㮖9���`��σ���H�nS��=U��9���
��ὴ�4���NA/RV��)?��C���6�ؑ*�k�St�3{�kn��Ce�>l��5�"3����D�.�;4s���
�c�G�Xz�@���*O��ЋM�p���:	Ʈ�kU�X,I�R,ep��[�M����Sz�Z��ɭrvN�RH1��v���:�,�\{���c�0뛛d>��|a�ew����9�u6OE�V�)$��1x��H^�V�?ZJ��I�~$$��! �`�V�9�;m�U����c��'�����д�?�>�%@G�q� ��IϹ��Ro: f�`�b+��"�v�[c�n�_CWj6#uSm���Rg����-ɂt[8O��c=%��p��I��E�B�$E�e�����_b�V<�(߫��×�������:g�S����A��b=;r-�Xq����_DVͮW��P�m�vuT���z��F�b�.X�SM�$�_�2����� \�Z�l�����ל�wf���1����M)G��Gj��S�*΄|�=4�����c~i=���/~��>A�=Z2Y��ޙʊ��!'a��pd��w9%
���qpn�ux��,�Su㳕㦼ٙ�P_�f��r<G��Q����g���  g�=����.˂ѡ�`!t��2RWM�Ez$}ćE�-��c���6�m�Z=1�=�sH��jk��g�ic23���W���KD�V�D���^)�����%�����c�3�b�/�+�Nkw��%�⤉�>Z�}����� �.�Ў:˝�p����rE��JP؉���?�Uf�;y�t�*[iF�Vp:&�	��C�Y5
^�f�s�1ш�oq��zR����'���Fk�T���/��������췦9o�;4�������G�#��Yx�����Cd��x�o�ٯ�C��#��fo�'��ʽ���^g�4�hd�m�j��t�~9�i\�7[~m97�u���Q�u �9��DI�yTC���pK�uB��y<B�n�*���Q�:
��!��P�jY�K˘��9�oX��F�b�-���A��jIi�`���K!��Ǆ@�𹧷��w˹���4E�`Y�E7޾���#��T���U��5��R�JA��j�4������P6Q��(��<�N��؇��/R�0�?i`
�)$&��'�������]��T����9id��Dw�m��8N���	,�3+-
�(�5���8��OPR0|m�N��`3���j�w�hyh��Pa$�3�宨�"O�v�(�?�PN1~k��j'x�ږ�yK���s@�y�@���I�K9m�\�nho���O�
�K!E_'G� 6���/\�"g��$K�'(�af�ݾj�o<��Gr'�R�<VY �@�N����{3ו.���8�j�s�'~G|r�!w
_T�8�B��?����|6�P���C���}O�e���Zy���-N���q�ٛ���j��8�D)'+g�	��QO�1�S�X��ݯ���q�P�����u��d=��s��hEwl��M�Uķ^�탸O�!��kC�{�+=|١�g�I��ژ��poM�V��ؑ�{P��94�-��v�K�t�.pp�� Sիw%~kI�|o?F���%��/��oX/7�}�T��N��:�%'/�o���;a��2�p�nόAb���z%,�K���,����܀��"[{Y���u��\:�#�Ğ�Y�V���6�Fҧ��s@�WI�)
���uY9�lDc(+��'v�fi��8�8��~J�EDb��P2q�[���X�fk����l�Ɠ�\�% ˍ'�4��Hr��?y��O���k���#�5�ڎ$�N���z��<Kɜ���L�C==Fwod���f�L�N��k9�,[����T�ƾ4���,�m";�:���{v{�*.˿;��^�b{3h�W���rT�S�!Z�֛X���
�Ӊ��w�i����5��ꮥ�/���]sӭ��	�e�N)���vvw�R�D��4���Q������_]�]+K0��/���h�R̖���l.��c��Jy�??�G�$���L�4q���j�y����-��Gԏs���f�	��8��o s+~E{�i��2 &c�"䯒3��z� ��Xx�{��?!�[�Ff���x���	�$�TxB�f�opl�r\|�&�7Ђ��S�������%Cw����*�Ņ���t�(ԟ��ĚcD�8"�|�������~7nwH).o5s����qm7KS8gz5?�0�C`)�5��I�gG���)%/�+�o/�c��_�6Qf�%�/(t/t�Ya��~�\y�:��d��'p�,*4�q�� %�ʙ�#ר͚���-`��ށI�Hn3���y7�A7C�1�
Dq��"!��i�������b�U@/T~j�F<�6:��Ǡ�re�@ᡟ���=Df(�U�ۃ�M�� �����<=�I�w)ty��-�f�x�`�o:i#1w��������N�C����}_��P�����89D�eKĄ�1��.������NB��O��Mn���} ,| �7��Q�ߚ�ƅ�N�iw�Y>��[�r��u=�t5����.�&�̿O�U�_��-(��Я91��-��[D�4��=�C�hױ�
�←͠�BK�ÿ��He79۽Zz�[W,��8��A`�q� �5��:Q��.@����y�DL�]�6����~���������6�p���D��	 �Eˌ�N�ۺ��d��o7�֗�D��?�@���ɚ*l��"%,�@H�6�t�h�����:�$�B<q�Y|�Se��qA ���D<�ݨE���N՞D,ym��l��R��ʆ�����&m�V��"Nн��ӕL�Uܐ�ۂv���w��������8�-7�^|T%;�-e��s[��2˸�����%r����:����n��B����ߖ��,�.�f1�t�/a�?�v{���H�Kp:�<��q�OΣ9�!ı�&SɼA�����.�ץ�%x��P�׀Rvľ�{�R+�qGEk�v�o�&����T<i�F��)g8fm��U7�A����Ѻ0*�m�*���A�õ�p����`?~�k�O�DYƽ( T]Pd�y��Q�ݰ��E������@KW�H�J� �d���[A���������m��a�x`X�$.�3陠��n�#���V0��R�w�ZKM40�w�8GM���G��D>�J���M������&W_ ��%���)��^���^,vp7�Bp�D�<��|��o���zK���\���]��n%Rc���!�3.���nP�@eR��8Y=�.���ʸC
�+: ��N�DV	�D;�@���A�j�'S��|F���w��rxhH���	L����Na%d��;�����E%�}�C���l��⮰;�}�,ݽ�>򰯺YO�[�r�Ru����893�XB����L ��^f�N���T���B���;w\������y�Z��J&cdL�(���l�9ɑf����Y���pR�(]�_�S��j2z�4GJ�m����,��|���Z>*Rp������Ჱ�h~ý�F��ʣ�^+������@��7��%J��Ԯ����	���л�%��Q�9�nW2b}��GsTV���J0����B� �������a+�D��o*�7KcXM�Yk�8ei=phǡ�уbr�[�X,# ���l���?�����X���<��2�ۡT��	�_(\�?����0�HE9gl\~|e�a����m�����"���9��{MA��f2�Ӏ��
�]�O_)����ZW�⿋��-6���>^9���37��(|��������jK(�O�����������5�6���kN	C��۴�2�{��Y��WGt(Q�s�x�eЌfTyО�!\�ɹmH���<	�����䳏�Lŏ�}W���?����v�(`H@]���x�~�H����o<	�k}��r�[��@C�)�6m�KBhq���#���S�c���n+(�e!����ͱ�)ǑQ������aoDy,�EprJf;C��f��zYic.������_��������F}F� ����":���� v��D��*%.��SD���p���as��>��s�E�r�j��<���gq�0f�i�"�oj��&��G�`X�O,�#{0ew�Ɣ ϣj����@z�����j��]��1�v+��Ʃ�y�6=,p�Ú��BY�nT������r'��]�1	�e�R#�/�^��2 	�m6��q��[���o�B�	Zp!���?b*��SC@�M��>Cݹ��%l��i��*�(���͕wk��׀S.�2�Y���@M�X�NZC��{d1�Q�M�P���� ��#}�^J�0��H�x겅�g��b����:�k���q�X}���Uv9����k�J�.����{a uJ
=4�jx�0��h%bo঳[!���F�@ؠ�<|��l8����UA�7K�J(W^��<Q�+����"
�vi��|��ʭ�d=�n1��T������U���ӪWW/3��56`�&`���(�������Ŏ�$r�[���u����d͜7J���}lfBASG�扪�lB��&����aM��g?h_V|&�2�o��Z��شMZ���D���]
}�/�����:��e���b��.&Z�D���G��}�҅���k�Г��D5zo/W].�Vh�ݶ�x���mf�8�\k���[8�����ɿ9�fn�ը�k�k:	��mv6�
y�R3sO�#4����?��b�]�7����n��q�󹒳Jǌ��7�g�8u���=�<��:�X�5|�\�,�H�X��� ��c�ɹ콩^
宓B�|D�2q3���?*)$��\�>���׾or�%��y�?�pP�Y���$�b�u���$'@ρ���T}50�I���|3]�[7@!���	�N+׫_��h0��m�C�V�O�����-�W@��M���Ud%��q�2C
��1+"��"8�}���l�o�)@��ql�@�7絖���O#��㒥�5�S�G�N��@��%�d�4������T�}���Ib����0v��1> ��{[� z��ޣ�MO<�rY7
����<�E�s��#Ԟξ(iL�`�}��2�[���MO�4�'~��v�j��ϙ��־��B��^[e:Ĵ��B����"	�9���~�����c�Q�z(g}a�VO1L���O�#7��"�sR��c�Cl��T;*���T_���	��V��p"`������K����3�C�B�v��qz2"��\ʏ����V��\��-m�.bo����a�����37�@���1g��4�E�^5���v����^8��x�}��j��(�>^;�����h�8��"�%ϴs�5��5�O��y��v�t��onD�ڷ5���k��v���� 8����b������1B��� �s ��������5�T+5�x�9W.%�:d� ��c+��;s?�(����ĳ|z2]m0O\W}�-�ڍ�Y�|���$cr4��ߴ���n�L
t�=ܠ��B%��k�wzL/Ѩ�~���bͥ��N���g����Mn$���?�K@��g����*�Q�t�G�}�%�� h�x�+Nf�NF�cC`z*rH7s��ܩz���8�}7���P��p�;�(�k�հ��da�6��<�:?rx5* uB�.5�W�$~�Q�t�꿓�ҙ܆�ծow�w��:�6͉a�s�*{Ƣ%:����jp����)��~����C��7B�y�[Ss��߹�d�� �a_�F='H��l�c4[�8��B�%�x�6�UyP���`�:L�ڵ�����D�o-�mv���*�lB��	��hb�L	�l����o�y� Ձ��%7���룦��BD�t���f}I����pB�LE��e�`��>��������X������.���2�f���/�(P�[��l*��c0dʶ鿂"����ʊ�zh*9��o���£o�����lSwZ,��.�H�f���TW���iePw�G��sC^F<	�t��,��G�M8�G@��b63D�����ؕ A�,a�͒�e�8vP!'�^Q���C���H���+꽫)S�crJ�]/�_��`e��&ȹd��r�A�`"?�0� ��4�Y{bnu�۶���Fr�l&PA��0(T�ZN�O���m-�W�6��\D��c4�\ lE���1nw�2L���a�	W�(�f��<�'�>u�����i-9I{�4�WU��5�P9�̣�Ǖ����1u5����P��O���L�����pogb��4�ʃfN�C
���i���&�׵�cB�:��R�f��Fޫ�
�Mخ��o�I�<�֠84��gxKkMQ�S�(��'��#@�r�Ȣ6��P [btMR�.2��3/�=R��zIz7��kC�`�y���N0(}Jn$M�@����7��=n�j�"?��r���(�E6��bI�ǐp������!c��(�q��Y(�1x聢�˹�P`Q��`���*ޜ �pI�5D�^S_�c`���!:��zq��L�&J�}��BV�_>�\p��n7}�s���)W���+�<6��T]��3��$��՘��UԆ8h1e� ��r�Jp�;"B�2N�J%T���g�z��7&e��Z��uI�t��������l��%����QSk��'���k�jx��=�%~�����������zKSK�=]�*;!4����NA<B$ˎ�ʚG2��Pf�r�\��T�����<"��o,S���n���/~q&З���=? ��B����v kg\cK���E��܊8��@̦�}Py�_XY�U�2�م��Q���j*��K�����Z)-Z�܍�oϤ���s�V�'g
m|�K�"�٥wP�}����>�y+�s0b��N���7 0oX�Iō�)��֭�f'�͞�j����Q��ˀ��ſ1cI��)��lk>!e�7a��яx�G�K �ŀ��c�Kyd_ǘ�����4���H�����˿�ef�mFrһ�e��sf�?�w�9O��%���$�3���=wD���1���{}H҉��^[�ؚ�&�D�Rc5����"�p��[B�k{���qL����7$�yR�rkf��ڒ8�:��S��a ��Չ����ў�}O��ẙ�~�Bs�5�N
B���q-AtqXZ��,�Ā�j���A0���y1�D�� N�M&4�~�*
au5�U ��9������M�`��n�<�T�� [���ôN�{PL��.䩦;��S�t�m��K�@�+���%�&��Չ�{�?�eR
���i��-���"��������|���3E���?Gn/IՋ,����Zs���Ŝkz
��Џ׉���o;lA������a�/���S��,e :K�e����ƽ����[C�Հi��g.rC�<+0'P�\s�iu�b4�&��JNM[�u"[��b��b����}zF-����]�
��|Ԭ���}���^� �V���������5ZɢBUߑ�KX�NEƘ�E���i�'���>k_~g2��F|�M�1@�V���q���Gg�;2g������}A,�a�L4�K���軦C���)��$"i5���>�Խ��.I�x�@M�|�LEެ7��N~��FHBg��˄��S�<�N��g�������oiHRJ�b�~g��NP�&)��9B��H����.Q)����Ɏ�T����ZW�+NB%�\&�;��B�;� ٌ҇�����Vu���c��/�
�X\�=�-N^p��N�6('����<V,z�)�TN�O�{y��B�.�ԧ122����ՋѰ���eb����S���X,�зr�!�J�ɶ�p�eD�$lzO��Q�D 9�$��-��ǌa;sN�'B�n�,�9O%�{��
���м8�b�Ħ����?��u��S��H�5���=���2ur�x����Y�#�p��l���̞G�#�i�q�"G�	��4���<Ц��W�s�3��a&�7��\#}�$����ll���{�Cx�v��eP	2��p�<T�������w��R����7����M�鯽��^��4�nK����ᡠ	b�XWL�Q�54���g��e���t��霣ݳ{�=��.�#��AK�>��4g�뽆Q�0=��t䰰<�3���n�!q��_��;Q�fla������e]x������r�Z��H>���efE��V3p�͈?�@˟R�2_
��a�h������5M��x�f��$�(T����d6"51H�<GrK��4Wݎ
�ϟ�6�9i���� 2����ٶ�X�{�+N�����*}�woM
���~��`p�!I���JW/�s����i/��>�z|jp��mBc2cu�㝛]:�Êvc�Y��_���q'��fkg��\n�zw����P7�a�Nǲ�?��5��v�.oL �.���K8gp%�$�6mb�R��*�.'>h�"U+6�N`�3rL��s�uUS��k*֠9f��6������hc���8q�9�
G���w�?C�BN݃�q9�nT�N�Ыx���;�^]�֔�=^��3�m�WZ�����НG��>}-�ȆöGHڿ�W7��[�®7[��7�v2Dz�8�d���C�H�p����ճ�1�L���;M����l��V<D����t3���~I���jY�RL�݆|�k����h��f���#�� ~��c�BJ��V�
��GQ q���>�+�nJ �؋x
g�|G���s�y&ڲ�7o�"/
%��Ѯ��E���{+��cW�-�Y�=S�ҡ�j��'��OT�T��ܖ��T�CyL���ڌ%�x%��j�����E�)���fs{{��k�>�`O��ߡ���h�߇@	��q@*?]�|T>��Q���g$r-�9�H�`��)��W����&*_�Q�e�kRW�fp��8XF�O����2�p?F�gr�'S�
۩I��A۞��+Ƣ,��x�*�e<�&, �xl&x-��y�9:S=�����E��������?u��榛)ǽ�n���Hl|P*3d�����8>^����v�
�C�D"�!��SJ��Y����S��U�=b{��������ϖq1���X������9	��;��]�E:�:CcQ���E�g��b?�T�;yM�V�|��1�.=9Kw� -��-hn���|}�w��Cg�gJ�U���ե(�җʤ��`�~=����@��o�Ļ"aig�T��Ag�ޫ%M��Q����@���"�Em3_���}E~c:#�İ��H[�����2�Szߟ1>��{~f�y.�=�ݪrH�P�H=�uo&@D���^����ӋT�lt���mU�88�����v��Й��K<r\�Y<�ڑ�U�R�gSXM�5)ťZIŔ��y*����n����Q�0C�.�<<1�	���3.I��A��+�_/� g%�[���~4)��_�s��.}ѹN�n9�?�R@�1z�/`����l���LNy��I�I[���f���ւ�<s��{a[�W�ċ-l�zW��u�b��z��yL�z��t�)+G�6yZ~M��U�>`�btb�r�\�S�MO�Z��&f�����ͧp����8�m��DD��<��)��9��Q�L�ᱢ�c���@��%���֜ke���嘏��x|��c��z�|w���/9iA�	�.3� �L��Z��D<����8�B)a"4�Kk5�H��S+j�U�u<�����.\��S�Q��� ��g���b��a,N�G2;��e�Z=u��s�SL �����/q��~U��i&����ә)�+���^���������BD����P�T���nzI[g��k��{��d9��傫�^����i�q"K����Q�\�r���k
�����OU�)L�2'G���`��ɳ�3ڧHL.t_��Vπ(��>�����|	ɧ�:
�ț��vL�Ʌ���7��N+rx���;X���'�y�g�E�ͷ)�s3o�����$c~;�I��cB�t��,������m]w��)�w}h��#�%���#�~��M�3�0E֗�:��5���/��h�P�$�|ᯭ��ebY����N&nZ`�����	y_P|�-]LQ�3Y�����Bj��
����LX���p����D��4�rp��$>K9�#����yy�c�aD�vŝ���aG��@m��rx�u�Q\��D�ѳ��I}*��=��(��h�5O7�R��'t�g����]�b�TM҇C��Q��^ŭ8�>��&�	�R�µ�Ǖe'��Z�@��%�E���Ψ0�Fa����"�"��$�D���t-�?6z�(����H�#���ۡ$gF'P�l�=��SK�:^�e�=��Jy�m��4�kgʯ�0�Ī`3���`�}'�dfK����>@�Dޜ����T1���<z&��[�C��r�Q�H�]^�y%Em�{�\D�h9Ej2YeZZ���>'PS��H��Eδ7���y����K�k�����m1�����e��^�w�_�Gj���XgL�����	��y O�x��t�پ� ƞ!�}�Mz����{a=5�r����!�2^�d/��}�`�آ��-�)�B jcGe�-5y��EP��*�Ąf�t\��FoS�ͫ��p%Ʒ߭5Ҿc��{�e�h�Vg��%._bo��Aj1RFv}�?Ma��J�V��d-UUy���r�����L����}1���ʣ!��R���|`hi4*6s>���ӿF��D
4�`�u�~�a d,�p]����*�j�be��S�����#���~#�}z�g'�?%Hxk8�����+�؋@1�1��
��1q��P����)U���ɡ٣��cPB��䋄���4���n�,��{���g�c��mת�j����Nע@�;UMbz���ǋGp����g�y����gT�,OF��N2v����l%�>k��~v{H	/�pt'�8��	������u�J����[O��`e�_:Ul .I�@����ݿ:O8�(W��+-���A�Q�Zw?xx�v"�$�3��<��k�[�|�Rٍ��!��h0��g'J���i[9҅��\���V����h�I(����P�|Q�v� GT���g{r�� uI@����`�Cݶ�	���l]�&���G��(��:27M2�x~� ǂ�Ц��K�����_�4��5�;duq4"�(�D�n�{�5�
�i -߉V!��5�>�׏�^0$f����������<>�)�X���8�q�k�(}�����*��.����>�lH�L�aՍl��i��]�i��fp�x�d\�]I�+����H��q���e���	�\7'"GȦ�"3i�b?���]#S�J3J_���"]���oR�^�3 ��N2%��>�[ݕ��7�2��g�PF�n"s�_}{5�S�G&��-��z,K�p��?�B�I�p���g�>��{`+�5�3��ӳ�D�^Y������E`3Ez>�&����݋|�idH�wg�և>�$���|0?�t$��벲����rt;z96ۿ��,�\V8ɟ�
bz�f��H�Ag� �0�^��*d��{8�fH���+�䞸A�h��+���M�լI�)�<�D3��.,t�����k�?Ԟ�TQ��a+��\���u��_]U����&�kT}�A>�2ץN�:�ϣ�k/�.ެ2x~��V���l'���� >��;V �I��� ��4"�sT�|�5�l��IS�z�2ZEU���Z��:q<�s�]G/��r.��9���Q�TZ�y�!D�`��9�%�ӫ6���4AF��Q��o@j�C&B��3p ��S~�&�d���J��t�I"���1��ʚ�F�}�g�cs��t�0T-�6P�P�����q�o�GX]�+���uh�V�ԩ���;܊�>���gB��3��9��@�)R8u��إ�EO�E���L9�1^�@N�G�����pm�PL�/.�%�fi]%[�%w�k��9�|I5�' O���A-�Rv9��g����!���(ƑV=.�v�C�~���6c�Ų��l��T�����3�'仝{&�@e�M��S���WN�I�#O�A"^��J�c�Xuψb�7\������ ��V�e�/AL���ӣ�z.YP�w��D�>Kc�t�&����=�&�J��O�A��0ӡ�5�k������&-f ��)�_� �<�J�*×�(�S��9A��~��.�I�»&u���C�ۦ:�h@Yޡ�>A�\qK����uT�G�Қ)�YWO�LT����ԡ��b�#R5���so/��u�t��|>����/N'�������se���w��	�!�`!4ZS�m����(���M�z�и?��C��*��h�8=~`���咀]��1eÝ~l�f$'L	���v��{g��R�1jR�ɔ�82]7��[��|�L�g���Ee]����F��/׉�K�0��9�������G��T�� ���h�OZNO���|-��l?z��2�p���`�X�' vۚm�8�y�0r8���yj��is�r�a�����Z�B �z�vT�A�ʐa;�#�������Ya� ��O*�kā,�.A�FN��0=n�I��$����P�(�M� Q������Վ����	L�5�!��
�&ԑA=�IK=�D�Y����"����C�q<T��/]
K�N��>��B^`���)k�C+�4����p���6L�	�p�u>������6�!�|T�{Zai+UE������a��N��K�����	�iQZ%�O�x���N}���F��aEޚ}�XS��J⅝Cc*^�6����p�O6x{A�O��Ҹv�Y��mX��	~�����m�,�.�?�;Κ������G|���4�5���N5���зҷyR���-�����K������=�Q�	���Ds)����g��WZ��p�l��4�A�
ӎ$���8Q�D��VSS6��9����[�y������դ�8EQ��*�8�Ʒ-���=��M���u��:�v��f�E	56J8�����5H1��]AM��s���:��ٮV���2��-g9�!�C��iy��?|%	.�h��&t�L�PF�s,�I���?�b/���|P��s��y�.�*$��'�
��|��^
w���MW��p.�)��\�枬�>���E��G{�^�3��b�̅x�J�Й�uq{iׄ�������;L�̠���K�Ya�z�7ن����Aq~��Fq��:TM�3�l����b#�\�.l塼��v拧�J�+a;�X�g�cEg73?{hk��GU=�2��E:��dD9��P=�d����!5q�K��6EK�����_�ף98A��A���/��?o)_`��hP�q#�)���;?�{�Y9� �>���{v�����ҹ���Qu*�{�Z#�B�z��R�W3:ii�L��"�:��[��>�`%�e\-s��w[#2�
BkP�6��&뛞)�"޿|���m�]i��T�QlkN,(��0�:�'����h��y�l� 0�ď�5pɦ��2ׂ��=T�i׫}q��,��8���3r��B�u<��U��jb����2-D�s���>�ꩻjZJ'i3?\Q�%��敉ۊ���qZY�Nɬ�~�Z�ǵ��}��<�NN��I�Y1��s���MS�v�J�c;^����[�tِm���wpD���y���������p�Ce��o���R��w�S�L�O;�ðu�e_7��Y�����)�)��_S��\�صm���v��`�+>%�$|k��f����I ��v���B����:� ���纀 ?�0��jxG��υyc�1�/OA#�u����e������1G���"n<����Xa ꬿL��xgHU=���t �dߣ�`EX��e���cź��fKc7�0r��'��֐��9��-�8�n�(g�4��`2���,1'ѝm���)p�XKϭD�*��"�a���+���'�G���q>&���c3C�i�܈��:6�Lb-"̯��g6�&�ش�ښ�#'�R.Q��
coJ!�|��{V�֌A�+"Y2�# p���+H �܃r�����'4��m�C��ȹ+�$`���^i]U}-nB����ǜ@���$�T!ʞ�W }*������K���3���O�v*����Fc������dr��#K�����-�f�:�S�nrʶ�.���_�GOl���Kg5�����r�a��ކ:�~�{7�߻g�WB�5�(���f��ʠt�-&k��#�����<�{�}� �\�f����`��y}.���#��N7;��5o̢���pI혖�ݟ3�?G����JAw�m/7`��$�"�S>��XY���yH���zP�GoJ`*�l';>D���ySqA�.Y���T�nx;�Djڏ؝tO9P�u��$1[�t���d�I�����Z��e<�܍�D�ty)��#�}z���Q3�#���p�e�>�ۂ��%c=?�Y���?�ʗ�X�l �����z�>�m�F�}�6=��Afqx�A�Uq��l��RU��2~��2��b������Ą����?�9zF��r98��1��-|��Q�z�q��Ѵ�SD�.P���x�I�����I�4J%��?C^Hi�r������~��_c
����og�孇���?�d~i�p��}�r��;]�U�֬��eb��t�7�i��5�Ԑy��N�u��QY��J�U�\%�G� EA�g���0 nRT��'�Z~])��$��M�K���kR��z颰�I�@R��A'���6]I��5��s�����'���|h.3�s��ǧ>�(�R��|Zb���|�gM�8�S�	�Y����؃�Ɨy�G�T����
}rXMU�@p/�������J��1c����?���}c/�RZ�3�"V�^���O6�|ga<�T�K�G�I+�_KId�m��%����%7��V�!E��V�'����i������D�/�\cׂa���Ge���Bֈu�,q��E�Ϗ�%�,S��1� �"aŜ#լJ+� �I!Q���d�%�F'�U�D��܊#����Zxn�+R\9�s����M%@']�A9+j���kS�����V���x/���'x�����/�4���;�f'k�/�<��NN��=���nkp�j���8;�zB�Q ���E�$t�a��o�]���75_ ��IEzc�;:�ӷ��Y�Z�N2]�Z�swt����˧t�`^��Xe�_m�TF]�4/8|��Y��=�������AJ4��'xu.m�b��]u�.��J��n?���FN�����R"��#��8�CC�&Rx����q�%��<�
J�6<�h�3�enZ��OI��ۈ�r����D���$�D!���M��"�?F��s�6��챂�#�i(-�A 	P�ߓ���t��}����S�@�9��i�r���q	B=�V��c��o� 0�^mT]R	W�!��I�l���X��}�',S��WG�'�xx�C��.�~"ӌ�ÊՇ���r�Y�*z����T���U�%�ل�"�Tep�\:��4�S�Nr�6@?�U�s�ݙ�|t��ܮ��3�A��b�!�:��V��#nȃ�Q8�8����3s�HL'��Ɯ1f��ّR}\��==�^�����B~{���\/+z	(-�Ƚ��[�k�Y5.�U��AL���%j�,���R��<�^��5��?��T䏀d#o~5H�M���'	�̌䯎�6��G�mp�NT�j�D3Q��2q��ҤW�5^tip:��I��p� ��ٶ�t�K��<KU��s�2�&�
�qt`ߒ=��A�jeC�Xĳ��DWl{_#2]�"^����E8Nj]�#�!�-s�����"=`��:�ʳ�K����5C���;U��@��}AlT%����z��nsF�����P^M����I����*�U���c�w�}� 	a3I���4��xLBҪ�����h�j���#C��I���Tg��r8�r:�@�Q��|߾M��ٻ�^�7S����*
h 1������B�F��m ��O^7	~ʹ�&�w���*G�D�Hh���U�q����7#3R����z4Z�����PZ���L2άPB�-�𹠤g��:��(pӡ�#E���a�	��ˏS�]!^g���sI��D�m���|�\Tc��Y��'�LU`w��������|����;^3�imҙ�@��Q5��3���a1P{{L^);�G]8�i��u���A�~FB��B']M�[}p�� V�߸rϵ�ݜ=��:Ld+�y���Q�ft�xy���-��6���l��\?[�����ܷNЦ�u��< )���.�������;lb�{�]��~TV�I��6N'��������Z0��8��h�<Б�2%(|�8����-��ڍ�Q��2Xb�ؾ�ȁ�X�hG��F4o��j׉�k�?���/���|�ɤ��2�j�:�|��>F�v�RZ���ьlċϑ���"a�4�Cj�����i�����i���<�a/hwv^5��>Q��ƾ�������;���v�Q�t�Nb:�Q���<L�%�����W��M+��`�u���Y��D�aX��yGK��a9�y��Hx8K�i|C��f��"�n£�X���=Z�T�M��$e�}{�S@e���$`�)�;J�6���M�p3N6�`!�Jѓ_Nb�kA�{�_Ф�W�5}T+2Q������'5���Z�B�����cQ�q��"GFFeD�ʺi)���L���|��{D��}�
6Z�K �Y;�	\��*�y�3���i�Sؐ���E�� f�M�!Ϝ*>c!���5O�E*KF��쿋�φ�.�.���N���8���4�>�����ݓ����M,�8��T#[��H��Q
�w�a/:�6�|g-)::#+��T�IF���X)��yQ.Tt��*dոڠuNA2G�'ҘQ�x�]�{?�A��'X���b`�P�r�,�SY����0�x��d6=�Ȟ��}`�.�]��<7bA��?>�J�S0+�)���&lZz��L��0K���1F,�8p]�M�$�l?t�*~��jw�oO��-��߮�%����U����ƻ�����̠ku�mޠ*�r�s��?*d{ј<��C�#���̄6�]�Q0^뜔~���l�lg-�{0�8k3�rs���k=��:�qχh�������u�)	�،i}}4 ��J�)��[<$�(�_h���fy��h"��2�+�j�n�y~��AkA��  ~4�Ɣ��~��[��;��	yd~���6`x-�>��pT��]�L�N��H-�$���k��^�t ���;�M�6%zHmGXY��;�ML�"<�D���L��[E�#�C9�L_?�~��NF9J�P�m3�&3��1���-�=��ŉ@��ܹu9O@	d�3k��[��Op`�;I6��^ֽW*VeC��(L�eB��!��2\��vp���m[`v�3����iʪRN�u�ls^h�g�tV�$h�Q����'�bI���)�S�1Q��g�&�R��P�Bݎú^���W���Q�#�H�iY��O�p���oC����_l��BFb2�J���|���������b��hc��^*�S,��P�/wG¿9p6���T^�J�Bi�~�(���<�F�?[y��"�ƺ�Z����.$�7�ˎ{ވ��`�Ρ�\Ԉރ�@Ʀb�� l\�b3��	k@;�D١a=�Z��.�&U��'��T��c�j�}[~ؾp ������3��餣�/�����
��8Ʃ��1e��aT;�R�.Sm�ſJ��9�%H���{6^�K|�iaL��)�[\�a�u�L'���UA�?I	�kwg5Fxg��͑�Y�6=���/⥮"N0#v����%��-�5�W�l��C�"ywv+J58��M�ƈHZt��$(������Т�#Lq)'|�M�Lf(�(+�]���7#N>E�+��M`!����Zĥ��y5�M����R��R&��Ml��16vhZ�y��(�s�sdN��SC?알���S�<C"bۜ��;j��M�1�ݑׁs���� �k9o��@����,�.�vX���<#�TAl\��pH��;��=�*q�m�X�9�.��d�D�A:U!���T.J�:�Bn��j��q8�n��(~�Z�+��!މt�5���&<MV�Xp)7�V�0+}mJ*>ʔ����Q{Aֶ�
=�nH��1�ȥ��"���NK�s+Ei�(�m{�0eBCK8/w6}���_G,�HR�D�Ǔ�r/��3�>�\����[��9��u�d�G�6��11/��S�DZ|g.�1���~=j��X���d%÷������4�������{����P���Ťd~d_2M/�����㩘h�Tl�YsTN��LՓ=P����J��6� �,j���h��en���'T����:����$��$U��Z�U���m���J%������*(&�1�Ą��D��J'� �y�d��E>#����r�6�L�oY�CW��Y��m�P��������+��S rڟrB]c8r$:	<Ǿu�$�e��,.�9=�rb���~ArREQ^yR�������yp��~>�?"�v�@,�$�֐�[��6L�@ E.ɭTx�=�x�1)��!��;2(��\߈Y!ٙ݉;�3t���R��Ω:8��M�̗��p1l�=H	�u���u��Ȁ��c,�[nvb�un\�QD�#�>s�Y���DF�����R �vjX�T���4O���Ft��mD��e����"�X�F�Qo1�����2K�Y/�h��p����
Xgpy��;א�hU���'�Z��r�}��eJ�$]��Ch���H\<
kvH��D=��Ҭ��<�p�g���,f��RB� 	����<� .6x�����t[Τܺ��H
?b��JZu�]GH=�X�z��9;�`2HVWJ0|HL���w��,w��$��	�bq����/��<��:
R\�s� {�W	�\�;EL"��)`��?p�)�-����D]�S�����z5=o�,����@���(�G�җ%*R�5�����00Z�~����Z�S���Y�h�+��%q��s���i~�1N6������ ta?5�Α�K0�qS�h��iN�2b��w2{�� n̐�}4�4� |�jNQ���XT)wL�s��P�@��,��c�y�}>E��C���>y�W�gd,tTIg8�
�I��F�&Gk��H�����49ɗR,�l*)���a��R����x�01��Y�B߿K�����w��J�9'XIxz�a�LO���D}����_f�\G��\�H��^��3_Ay��0[O�ܲ&@z��T�6p�7��^��R�%?�E��R�%쾻P������}I��x(R^0��ޣ��g��oܞRQ�eǐ�M�̘��Gg�HyE@�l��v�K�;5��.XB��a$���H����,N1(1���L�{p�>>��[����7�8�lHkg;GGΛZ�ڱC�|�ΰmWw!B�[!'3]��d�E�:X:���t���Wf�̮�'[�����1���Q��0��S���wW��i=��-�=���f�n�i�
蒖���,��F��W�Wp3�It�0�)W���XEޛGE��.`��p���\U����#�^�n�Y��k��t�9o�!9Wc$԰'��=��%4��nn n͝����$#.����V�|��4j���<V��bD���BIdvK+�H���CP�"1[�e�RFg�7R4�	+RO����{�𰇙���6$��tK.綥-�o�@��n�~2�2��V(�I�I��x�'�;�e��
0�A��1�ȇ �
�@bh@�-��-��3u��F?Vgx@�l7�2�uY[�s@�"�5��]z����Hg���t
����v嗗@�|l͜����� tN	yݪK��e{C�#��T�y<@�f=�B�� �[�f�Bx1y���1*QMe�)j^D�@����V'��N� � ��i�#L�X�k�xA`��퐻n0'��M�]J5���e�g�*�]���(�ҽ���h����Hs�<T�vX4X�Q����N[�^e	k�2��FI�]6�N2���CUT�G;�0�RY��j���]�j����<	�3jt: +,lr6�N��h��x%�AF��1�u�ݪ�ٯ�P��[k>"���KQs"S�B����)V�9*�:����Es�y��o{�ְ,���ǲ�%���D���{�a�&
[�A�������]?m��Y���V����=���bfW�a%W���U��kK�/�]��s���~���Q�KA�z�f6�ۛ�?,B�ئ������r�{���`Zqw?�����f[��y��B��ҟo6]��p�O���ʍ@�V�`иЬI��׈��h�E/�'�\�r�WZə����3s�}��}�^�ej+������Nə���sK/rٻ]��p\�w��aXÓ�!"Zow����X��8f}�_����%�Jw��/�{������Z+f_��N��j�|ٍډ���vV�~f���s��v�P�w��,���Z
R�V��B�W�A	
�<��h�W�~�� ����F���^�àC�ԀO.�w�^��&��p�~SG��L��-\뉧�-�|&7���޸�gtYJɉI�����ɒe�k��9�I���t&F�I����h�����)bxu.$4-��~�v3>TH1MCכ+4�	�7,������i��0�C���>'�䶋�#�#q�����T՛:m���)׃���w��t�! ���<���W ���4%!`|y7H)|�i×�r�I�SF~��I������� b�n\ H�)�wY�9m�|7���<�ꠢ+�;q�O�ұ��{WV�Q�2�-�{�� n�RQ,,c���>����fQ����Q(��j��a8��tS��%z���tH+�7�7]%�r�_�_�T�m���)�:x��h��a[؛.Y�H�R�Y� �coQ;Q�8ܞ��^!+<�c�(�AV(���!2�L?JF�<N�͒h�H(�I:Ͼe�z���L-EH^@H��b|l�⢳I�ۖ"hl�@��ޔ35�bVȃ������nP{���34(�:G�pL��+����FULxOu��(�7e���<2e�L|���OA�"����_ЋT������%{�����G_3K�R��P��i
�:��z ���:�@MD�q[�NǅY���6D;�v�0�<!������^�C�����P�8�)�\?V����XH�d�C5�u� =��G��)Q��4,"9��5?�>�'�P�2g2y�҂iC]�%))r#|"n�|�ڼ�^^�(dZD���Tp�k
<��Q��Gze5T��[Ծ6�;@��
�ӣ'�#{N�}���"Q@�Z�q�N4�,�8��1�:#z�p�l���P51��E�`�j#kj򕞖��<�	GL�y�EJ��YG{@����@ruM��m=��+�}Gl�E=��F�~���)B���9��ԈD;b$�A$��ʱ Wa�דIf��֬9e���������'���?;��'��|���k��^��l{�Թ�� �Y���A5�̿�ePE�!U`:���u1�i�xV˩�k�e	�װ���I���(=�m���jh�}s�)���x̅i���j��0\�1�Ϳ�FרɅ�	nx�0������z~��/�+	/�IL;/�������`��U�oPdW�?|[x�>�<�M��dIUH �4S+V}f�]�?��9mx�Qb^�-��Yk
����}=����"�un�Ȥ���������	k��8�d��)��1�o9w����ǆ/z,ٽ���gv�Yj�ϕ[?� �e#{� Z˳ئ,!�$KMc���̱1���Y����]}�sʍ����'��J|.�����ᲄ�嵩��z95e�Qq�^V,���[��f���ER0��洬���u�d%=�7�61�\��b�pGh�y��ŕф�V��^�N����r,ޝ)Ȫk�P��E4��6����i�<�ꄕ��#� !��s�VԺ8���]��0��/����$K��U����p7��4A\
���JW@s��7W�sg�H��(Kd�""l>s�Ɇ�\�6����`١� K�����PN��GASb�E?�}1��ȸ_��?�!rQR�����.���8&��sq���f���D4Ql�pp����Ƚ���ԁ��;L�����X{���w�#��j�*{9������\��$2���,�7��Z3e��4uI��8��"��1<M�|@�_���Y�&l�N�����܃����i��ų�>#��6�]�ǿY2�.|�f����`�M�������[3�x�~*|~=����i��ĭa+�c�%�xUD�J�Ͱ����;<D�}�����4�?E���\�����dw9
'�>�\<�$�!��Aj
�ed9P{1ϥ�IJ�֎�ɐZU,��.Ow��O5�䑋��"���zd~��vm��G��"�o�Z #�e�.z|Q���R ��a�ޜ���}Z8]�z��+��\�V��Td�LZ~�|�lʒ��:��
{K���O����!-�;�;uрK����� P)X��g�7��͜�s��S �M:DT�_ƲDU�xz��|�y�����]K�WNA�b�DҾma&v�Vb�{��Xp���nQs���ɾa��T%s3Y$4����vU;�T��1,/
�Jw�ym���JWo��%ܴ�??�ȃ0�� �vG12�����׾z]�~��H)ΡX�W&������P��I�EC
��\B?�]���gFzu��W ���W~}��o�-��D�X�̀��nwu[ih���Ff�Q/�r bv�\WJ�lM4�����Xvd��}k�k�L���u�A(�6�5��Bot]���Zp�uIК��í��HĐ����o�|a9������aYp�C�4d4b ˞݊���٨�Tv�B�]�E뮠�3�]z����Ua�֯�ʨ�܎�@DŅ�B�r��Hvf��R��D�pL�z���_X�?{g/�?�G�����B�`D���_+Y�媄��B�%ߟFw�e_]�7W4 �o�6'�78(���wn��c�/���ڋt�A"Y�wW���5e���B l���ɸAke���և�lY�!4zZ�Ȑs�G��wh�?�R�k�Cn>��_f�n�.�M��N����\	����o�����%�g�g3I���<��5=8�Y�Ҍ��x
6���E�q��C�o�F��!IqQ}���"s1��pU��=����>\N!h�R�7q��4Kˮ&���Y� �놞�+��B���Oƽ���Ϧ2�pW�Z��2��D�uu
���'�.����X�h>"=�k�K�3Z��	�q��������`����1C�Ӫ��:�4�����D�*�$,kb�]2��1�ด���>R[i�r$���Ű�Nb�#�r:�|�1�H��]E-Q�3�@���?f�E�� 1%V	�7\(��܈)A�&E�0p�3�³8�)m?�X��"��[֛����(^4�(-�IP�	�A]�}r�8���"v����
�j=%�*�K���Y0F��A,EV�8����l��)����o��
\ӵ=�M[�_�!PI9:l�H>��"6���9�>1�_k����[i� T@��0���!�+�"����?�%��HC�-���C��j�.KyR̻�����EB[�E���'�Z	�e��	4��*孓�Y�D	�l/:����O�螁�x�gO�ʙ���+�v;�El���=�^@;���L/�fR��������� ��-+Q╠���&�l��4�]s��5>��aƒ�Bj�QSf�?��]��ʭz�_���U��j�%�7v� 7ćk��k��}}���4e;+t%% ��@��QB�����at���M�H��έBr䤴��9�x����B�<=S(���$$�Q��_4(݊���݊�+�_Z��.���$4�EL
��9�=�&���/m��4X)Nn�2�l�^�	E�b��D|���//�v��b^�H�{��w���. �R>#�T�b[5��L�`b�&�󖺎��y4�ׂ���I�.��^ׅ��*�b���SYB��S"ld���t��e�%9Mj�x��`��W�ʹ�l�Su��M�
{g���*)��xJ���R�"C���
=��վU�j�(+DO��
����$�O����Ӗ���#��ܑ��6bKrU�5�0�UYP_�vB*q�ٜU��f?�+Sk�̏��.%�Y�|��b�2�i��j>��tR�����������\༟u�Fx���nÌS��L�� �%,�/ѴM�3���O �|<_#��8"�X��l(e.�����:��6x(u1��ʵuU��:�������^!~A�)
��'5�O��Sԭ"|�](���0�#�9�����C�x�ǻƭ�S�dж4$���$!R*29)3@
6�p&�/rǸ���NCe�f��?7���r�$}����?y� <���G22�����՟��
�u��N�Zy �pcg(&��!�o8�(8ט�.Z�aT/���Ѳ"*��5���O�m��*W:m$\+�^
���3�։�dp�+���t68B뮿Z]n|�?����đ��zEBoO$k��Ǭ�·�.�	ü��JM����R��x� 7�۷d��!<��4��&�IظL���	�ao;.�z���?]7�uS�F�l���/��\hw��)�����F�zK��-C(&� ���	  q�����y��S��J񊌭��W�kV��?ˆ���i�g�j?G�Ɔѧv�f}Qجx�_��
�ZB�f�Σw��=� �㦤�K�U1I�i�`��u�4���KHH2�^����̆�}Hq�c�[��]�ʩa�d"����HKr g�*I��wg�]Hv�'���vh�M߆~�����]k�A#[II��@+A������H<7J�)��� C.���uR�{�|�4{�8�Ed�J��T`��?�n���$�Gb�G�'����=<Q����(����K0�8�٩�^>B��d
"~��iB�ΖReO8S���l8������_�J�R���(Ϝn����œ��+�U�k�ɩ�en���� ��7-�{�������٪K��%��hC�Pp�y0���s���rdb��I��&�i�|l�1��Z����XcYj���.o:�w~?\{��z=���bBBm��3,��>6���W�(�Hc*}3�T�?ͥ��Ή�i~��cmL5CD�@J�����Q����	!���j4�ެOM��J=� ��/��:�~O�\0��d\��en��j��]+���Ɔ�8ߙ�V��p!ev��ԙS3��y����D�j1�2:�h"��R��0/]��W�����YR����~�X��빗�����X��]]���Cl���Y#�B(���g{���_=�a��*�[J�j�COD[I��A��p�)a����(�8~7?���Ye���|��Rx���5O=ab�|���qZ�H˲�����a
^s�:�[���q��6T��8ylZb��x.)�T��uB��8�W7���Ey��xqycA�m������Zx�W���U�5���x����d�Gr���X�ג��T�a���7U��o�p: /;�j�V�)�/��l�p��n��pd���"
�>�we��h+c񄶣�f_�sW#F��r�$���?^����j+�9:��3� Ga�-�2Z;�|z��Ŝ4؅m*��(��U�n�<��'�K��/�d�S�Qڳb��Q�� ����E �y1�ß�E�\�<w�FKl��,���\2�:���7S[�ۛ ��b���^�� 6��D�� �XoXBX��ou]�x����6����L���D�P=�=�Z�L�+��!�Cks���L������~8ad�/OhD
.�,��)}��F�i	m�T���0\�ņ̓$���ܻ�8K(��+ġOy0��4�����^A��r� ��ph"�G�B7+l@�� �S��TDkP,)���9�i�ǒ��*)H;)�b:�a�,�u�{���q c�*��S�8o'�=Bsϧ۝	����c?@L�'�"�<6A}{�Y��d"t���/oD��%r��ӋA�	FPĬ��S�>P&BU9���`�g0 k�&o�3�F�5?ÿ �B�!6��u��ų �/� �Z�A���,$O�i�S�57������4�?c'};��h���g�RB��b'�h��'ĳY?�%����ؐ�W�D�Obe�K�;jpp`��j �=گ��U$׏�;�S�A�o!�弨7��ofs0�f�J۸5�}���:n;C�Pz'��հ7��z:
�o��t&[es?K�8)��*�Kn�a;��������'.���噐TS��N�)Z��g6�{���rA�#�r�¥��^bGj��}}�ս`_�\��d�8��C{�n����K��e���� ���(��@$�ݰ��g������?Z����&���@7�	�#��n�{�����+��A�3����J��*�lg�u�k�IT&�<�b����߉H���8t\|OrE+����Gv#f��&��Ӡ��2y���wa.ʙ'g@!�:++{�#��XL�Ҿ]SzW��&Dh� I����6T*�_�Fw��/5X>��K��	$+,3OU�:�vN'`� 婿n>1trR(�>5�.�j��Za�N�����-�K ����+���|���+��Bb� �z�9!����e> �&�
�U��$zMN��~�cr��%��Յ��^����z(��d�a�[���rk��e�K�HZU���R��(F��2�tk9pY��薌�k Z)�߅�,zc(�/��w5�^1�iƴ��P�_>^���LM]��L´-��Ϗg�9��^R��5�0�џ�y����o��@���]��aH;^��mY`��Q<)���%Ci�� Z|ws(k��9�I��]f�	3��Ar;p�!��'+��|�{%&�ho����v��g�H�B� ��w:C21��D�$d�n>l��:8Kjx��FM "�����DE��M+\?��/��H��D�O��ĩgP���3Qu=����mj�/����!֟?��v�&M�ۃ�k�|����Q��NE"�w:f����R-#�O��� ��~m��&=����i�2\��'��%z���o����n�������𘊐��*[�$:����R$��뉃%[��ɘ�ǟ�ʙ��m:CÓׇ�|T�9:L$ԳL���yq�-�E�G%~l����>�/�\���{>t�~45 2�e��%�3Ű��J�����y
�d��j�a�t��6���= ���l���9q?��I"|��?&Ҟi�N������A��Dt��5���r�d��&V�
Y�U�?�����N��U��m�I��N?Hu�h��1�>�w���3��BǶL��̥��:1e���pW�� �ߥgioNM5�vGN�ؤZ��#���2���2VL6��16�Z��8�H�'j&�^��v(�>��r���J!�z�Q�ԭa��B/ZW��?��P��I#���4@"Nݵ�i�e�`�$� ����8Dt��z��"F	��Y-���5rh*6~�����\>!�t\��K�	���z�����$����gn������r�V/ [�i}�p�M,m��W�\�؁Puhq�o�/�l�~�Ȁ��>�ezT!nI1|y�A�E�aD���E��	�v����_'��jY����
���w����9��4�,�=�A�v{3�v������
�͜
�ެ��u�y����d%$��Q�)�<�a�ղ=I���:h@\�ɚM�%��ɅJ��u=7��5	�B(�~W�!x2a�� w�C��Q���;��AFVq�i�F�1�C��O��/3�W��>����f�U�挾��RF����f�Ś��ęI��k��ތ)..OĈYCV�inj��`s�SoG����XR�%[b������m�}�g@�;̡�	��p�]	B�b/��E$m�M������xLk핟\I��S�[|�b�g��j7�Q�P)T�w(�k� `W 'X���9�/6�q9AP�X�بLv͹�K]�|<��0�EF��a����i�|ê�_���6=c�򔬂2�(���X�CM}O�➮^�d�.}��FC"�^��NL��hC8z��b���R�x|C���1Y�h;��3i-�9�X�}�'��*�*D��8Ř씛 �Q}J1AQj�iÅ�.�V�".�*54���G'Y�"`D�.l���	g':Ѣt��/\������lڭ�@C4ֽ��w��4'd���Z�+XM#=\�~�Y�� 3�Ί�C����wȓҧ*3|�^B0�$>��Y]�8���jǋ�q�&PqN���)4�J�*�����S�),�'�q<\�� >�|���,i.����@�Ց-��j�ڨ���#n�������-�
 RZ�Eh������z��������O�2���_69Ž�/fA-)���"������wh��J\�֬O9�M�p�v@�(,��l�[��­U�x��L�ÚZ�����/��x7�nQ;�?�td��-�euY�*�(Ć� �����8��n��V<	�!�́3r@*J�8��"��O�-9-m�S^��!x�r��?�f�b��Oot�ч�;�;��Г���sT���u�+/��au�{qR8��5��y*��P���1��巏g�"�{Ҁ���;'8s�Tԭ��q����'�ϴ�5?�ԇ����\�gѮ���"�r�"�~W摗��!�J
�*F�FL&E�չ��_N}���y�k-��Z2^�H(�*:R�aH�����U�� $Y�`�:IS�<k�h���z�{mǜ^���?��u]�T�A+�]��;�D2_B���`%)���#���6�|%!�)h��@�C�On*"w��.s�:ԉ��;�'EN�����v�Ü���yd� 5�u��:�b|�TH�@�oŌl��y�)�R����ԣ�I4=�IYw�a��s4��לI|���Ӆ�<�,嗲��s�:���6;�w�yߏ��#��I%��-U��7? �=�8���s������@�=y 0�\¸B�	j������;)82�R 댁�V�y�b�z_�Ki�2�d	�<�f�[h���r�LB<��R�Ҍ��g7��z���
��4A�o��;v�B�n.'���D�N~v�x�A@
OP�)-�h}��GB��p�>9�.O�v�l5�-rr�5P�K��^;�o_ �~Iǥ]v<��Z@�Í)8#8mx�ǌ�u6���w+6�s��ԍ<���AE��EG�!hR`�@ �� ���y�*!��ϵ��z��BY��D~����r��P3�(V�	�Ƌj�u��_�%��КƦu���h���/i*h�4^W4GC��>u�Yr��A�SMӐ���&t(�'yqD+�7�]��~%���C���S�ˑ��yiP$+G���6�;�� �5�\�[��#�1�C�܈��٥L��	���)�,���񏈄q��|܈Wr�63�CM��_�3�*.���.7K�0����	��uc'�a�!s���j��#ģ���&=��Xٔ�p�^��a4�*��m���2��R.N���̏��D��A��:�Cީ���i�F�ĥ�h�b F�*�U�`��p@FW�m�bǂ|�2�_�2�9>9����]����%�$>e���\yJ�S��q�15�ɒ_g��%'4�S�Ǎ�$�\�٘��+8c0`Ѝ%��,��
ݑ-������<f,ܾ�#�V�A�[��:��;�ny�׉�̤�˨j#R���xݧ����Yϲ��#���:�݋0^6�	}Ozs�)"��%1���V޺�^���UQ:>��n�M�m"�"�6��{�"gz��3��GP�
�G��ն�j ��sN���s�Y"�u�!�s�tp1E�|���I��!��� Ɔ�����.�����|�&8��ݧ="3�f�B��&���U'G	H�7
k�J,`��	��IA�f��I��x�n�/�����C�=����]7�"�ۄ@�8�c�D��-��=V��1�$ƾ9���!�i���sA��U�A �׈"1��a{Yv�]�7۾��HAwmo�a�'P/���0�f="��S�EA��*E�.҇A�Knu�}�֓EJ'�Ϫ��ȿ��4U�`p:��25M��,��FŊ�
��ܗ����@ɫ\+��n�b�N��N�-S�L���\�4f)����$�^��?B�!Z�}�tǅ(#D/op��T�|�7:ۂ��6� ���A/���uB�u�0��v+@��d��N�f��!�̟����q<��}�z�b �z_��8����\�!c��J��9��c�'/B}�V]�J��5W�����0�Y/�{���zM{� ��I�Q �WL:�&�Q��ds�~�[��A^g#�I�	�<�L�$~�7I�9X�����粢���7iԁ�.��Ξ�wa����p�����כ�`��;�K�9�i�̘^NN��rhr3�m�G�N��Wa���Jͷ�ᖀb�`��.��	�n�D�\�:}�u�+�98O�ķ
/���&en�*�>�ìE%�(���#%�6!�y�����[��C�:��#g)��;@���TE~�������D򅗍$b�NѢ�,��Sxj�����(?VJ'�ɦ��+=�Q6lيi���n �TW�S�ϙ�W������67uK�dOT��Nź�"|���V�8�4��]fOZ�r��Uf��S ��o�`C׎�3��yW�����|Q�3�i����F�WG�����:����0�&h���}|�p�5
����R�v��#��K/��$qC��;ʽ�ܡ⼹R�� R���4��m��Ej�Q b���.f��d�S+X��:S3���1;��#�7���"k|����g�DQ�R]M:%ޅ-@�?��k��,-sw���c^��]�f��py�˅mFY~9� �����@���o
�������P����~٤�&S�p<i��y���^;e��˦cb���/�;�Bi{Yb�~��e���Qd��kp����%R�4OBt�̭1$>UŴz}٭�S,���ª�R0y����r���G{x��lB
�B�=�:ͮ��D0;�'da��py�=������Y���;�%�B/�QW��^�z�)Zvl�\+E�R�ra8�� ,���qt��y�Ǟ��a�m`\k��˴{�P��ϊɡ�u._Tԝ��P���ߚkwH�,�,v�$I�
�a���jX�RD}���A,��o�s'�nq�Z>l��q�+�� b�t<��01��K�̹v��u,���c��a� �-N��G����|W��9N��L?ڛ)k{U,s�>����ELaЪ�"�.7��K".ʸΚv���3�l�#��'d��#�PE�1xGW;�����B�a0���sa��{��aq����Giq�6�Ͽ���z=�~	���`�"����H1�{A�n)�#%�0�]DA<yD��R��ʚWp���y+�o�� �K����6-�W@~�(��WH6�����
-�S�� �(�-1Qs�{ �Ɯ��*�ld�utZl�|\��]���$�����aؼh������p��JGc�#��?�U�`JEW�`>9ɋ�F�{[��V,V�r�s�5���hĤn�2EߴH 	S��ac�����y�NA흅�嗒[� ��I}�h~\A�EOTJ=�&�t��W-5���Ff�D��<y��JՊzh����$�|��O�Pt"�'�.���E�����+���7.̏�7����Ob�|���:�0I3��!�T�FLܤJ}�EX�~�����)h�gR ���/�g�.J:�o�x`�q8�^ P{y��\m���Ð�w�m�*��r�:������򊜩��$�f�{��arF�E�A�$�$U_�chf�8q����E`�}!3O���פ�&�����7�U�f�WB4n}ЗA���R�eӖ���fV'�$���b�!��D�֤�Gi�6���ʥ� $����U�*�w{RH?��V�_��Yϴ�sc;͈��P�k!�up/�u)��upH+�3�(��}��a>Q�Ċ��|�R�������T����͆��W]:�?Fí� _��8x䠒-ڰ������_E�]��8ؼjxq�����\ ���4��W�yZ'���0&6b�Y�Z��5hy�ξ�!��f���]��Û�RQ#�{�z���L�z ��S�F�6$���L�@ W��8�=��yY�Q�A؂z����6@� 2����4;���!�ʍW�p��C�C-� �_A�ڸʰOU�T�t~��\e�y�=�˦��~b�Rn�c�e�N�-�"���K���K1�K&#f��B�r q�̦���:P�{�Ǫb&�?����j���F���1��.4�1Ȍ\�F2��Jy5���j��3^����.�vJ��Nu�����˾{���@�W��u�m��Ѩ��wƪEG��9�ވ�[1���Uܢ |E8\vVf�}��jg`�|�f)�Y,�_ 0`X �#&�-��TPrZʈƜ��vE��Y������V`TUE2o��J=_A �G}��E���F�o?d��	־�'(�>L��ӿcK�E۠�7��c�+��s&7�)�,A�P�U�Ƹ5�Ale.<gΕ�Y>�#b��ٹV`�y��d�H8ho1��Ð������g���Zu7�[�R��2J-�.���;�ɛ�H��qn����i���:e���U��S�V�k�jUJP�:�mZ�����7�)R]N�� �ˠcY+bq�t}y��׮�^�.3/�A��2��kV�,�-��� ^��S�/Z�D.鉭����M��_c'��������Q���c)XZ�p�0cI"5B?7�0ݨ��h P��md�P(�҉���.�ҥ��F��6���0���I�Fm2�S1N+�0��IK�z��G%��W�Kxu�PA��V���{ǖav�p?� �D {lP�TC>�xߴ�
P�Lz��S��C<݆ݸ�[�Ҥ�	�LW5Aml�����^���� �ν�ݘ���F3\SL�3�2&	�N����#�wΈ2~2��Fy��4N��^�4�KF~��D�B��ѷ�'�:?Q�kfk�.y���n�Q�v��#.1mg'��v��-��8&~ꊢ.bmH%�P��B,�8��Xt� �U�`(E��gn�n�I�_�L���F�<O?ײ~��R��7�(���ш(P��pN͈p`c��҃�����@ܩ!��}�f	�0�W:ͅIE&'+��L�C�v��O�7��#��S�Guz����]8��oY���������<A��}=�{�v�8:����j��X����(T�H�LMGΧ����*���V�ӫg��x�;3A�<��#�����Ckg�b\��Qhe���u ����O�Sժ��{m�����a9a/����т��$�f�_�s�_���B(�;s�A'�vc:�s�'�����Bs!�'4G����vM����_ыN���dܒ��4�ՠ5>p��O��u��H9%C>t�t2��F�@<M��n��[Ul�s����ޠ�^������Ě%#��2nZ���ȓ�$�������.�������NR8�6�Tw�M�I�{�e��ӣ�ۑ���i.d�g����'#Y�z۞];��e�˖N1r�?��{�fQc��Ӊ7��e�;\.��D."`Ya5ˤ���Z<�6޵1��^-H�5��� ��w��4�g1�l������DD��<G�oڭh=��p�T��3��QF ����~���F��x��� �=c�i��cYo�(<,=�ǎ�8xc7T�lЃ��yCr���T�	���.�H�)S5�&�
���xQvE�*5�d�`4�ى�:�4�'xck�p�������#,��(��jvE��H�0��Gr��ܚ,�Fϧ"O�>H��Kp�5����i$R��11��jl�|��-�-a�e�mȍw��nb��&�
��mo�^�,���qFu���L�9D���&����pON��n���Ĥ_CJ�\�ጦ�V�\`�Eg�xL�^�L�2W�>���r9r�]��8s��Y��V19O���b8�2m�Q�l-^�X����	W[�R�6���^���?��_�^�
���bA������?�F������J[x��/]��Y���j(�B� Gl�F�T7
V�Gt_sEA��V[k��g�m#� ݛZGB_0�+�b���F�s�:;�Z.Q\��,@��!��`Xoe�?�1��E`��{�֭9�D�u�7�(pN�~�	���q�Gb
o��&M��&��}�����u����;1~�P\�UPe�J�Cq��+f�g$]~O��*���u)�U�M}��C��8�l����^ޮ7QN7S�dO�|�4v/w�Ȣ��.�*=9�<t^B�\i�&��$d�w`9 �������wC����9��=9*���15o)���0�=�zߐD��k�]鞃o�H�3Z;�**�3=�����w9+r��N�\�|Mg����
���K�-�,�VV���q)�Qb�fƀ�u6�K~�ﻂ������n�Őm�(�$�^��)�ei0�x����0�`�c����B�JzGj����ф��~��<`b���z@������1�w���Wq>�,�&�U�� u�1^�:~Z����~�o?��c�/�ro逐4�����.Z�H�wl!,���VoԿ�V�X�y�X��i}��m� ��0ᩏ�\��b|�W!�J�!�5��ȼl`�*�}�Kj�rF�선>ՖX�[r0~N������=/|�5�lN���y�2�.��\�%gK<}z������7�@
s����3M/��������YÉ.?Q��7�����:��	5=�䑂ŋ�9����ª	q�.F�e�;;�������w����� ?#��pB�v���9�7�0n�$������P�覚ȋ�Ǎ
��I`��E{8�^g��vGJ� ��7��1�x4_�(�ʜ��г�	�S#}�J:��lJ}�`Њ��[kʧL9�=�E�9$���	"����ג�.��e�^�.�d�f��1*�" ˿Qd��S������GrTCJ�y�Xߨ�a�����VYfWR�)V�z�b�5�SK�.Ұ����^�yY]+���F2���)Җ������}$9�&�N+2�p}�X0�o�<_!���)�CI�AVg��K�pF�{���@E4�$�^��Z�c�n���s�����:��C����WU��DoO�q��e�
�x�к�\,>�h	'��C���ll�3��H��HQ�12=��v�fG&&
a}�i%��
=J̛Q�Q���W&]�K*�l���\��d�xľ��v:��fV�7jicK����g�f�f ��l��a�,�7��7��i;�C�m��Ѣ�]�6�.ؤ·q^��2��qPw��g7}��g����+�)ہ[��}��(�|>�d�q�1hѐ(k���MŢ4�eA�q�Mm�q��u�Ņ�Iŀ�w��X�O�gUB\�/�AaQ���"!�^�/����������R	�\¨��G����|'��4�e�+�g�3]4d��t� �(exd'�[�����K���S��mSoY/��$rz2:�"���#H�7-��B� %���w�يS�(�2��i�R�z̱����1���as����tи9�Lѷ�p<j��̓V6���zվr�SCnU.�'Pҹ;jpӧc)B�e�����K�D[��]�y[����Ud� �E������~�\G�����������qЙ��y��+ ]T6"c�A�?.c�8W�Q=��i��CY�7n���%`�����Z4�fީ2X�Će�>#��W�F.��]�PZ�Շ����پ{���ָ��.�O��v�{ >F�1˄��ܮ	�ѺS�R�	`h�`�u�e+פ��Eb�x��s�2���0
��!"*�e�V���}6&����D%	��}��3g�����L�F�ղ
�Tt�пL���r�f8�)�Tk�OSTv4��ޙ� l�acZ��Ʃ+��A)��3DE��(�c�>d�	a���AT!�������vՀ�f(e�9g�@�\�T��z;/��!4��<A�|<z  #u&@5�G�t�q_�ʈ�3��%P��eG(IO�N`�x9:J�r�0ҩKs�ӳ�pQ��+_�������7��>�X��rV�&�)������h�Ho��
��Y���T�$Xl6�W��R +�j�=����eP��AO�7$,Oٽ9��Gz:�I�1[Qn�?�%�u�YD��_��d���k�ʙ|��"���]�Y�y(�AG*v����=����׺��{󘽨��0p(�j1ڄ�-w6��+6ٮo�c�9�#��bΥ.0��)��c�V g�Zc'�n�NEuYxVT3X&p���*�X��׹#�xC���j~��<���$��z޸b�/d�bWR�1�"*M�wy@��Σ�%gc�F�M�����x2��[eS����߷_����վ��GɊT�kV�;�p�7i�^�<�1�h�ܠR=X�i$�ȏR�,x)�"�#-X���\բ�D�Gg�A~�����󐈸/bfA?��0-AF�)�dk��·����kT^r)q7grp�3�X���a%|�CoT�B��Pӥ�������ZZZ�6��
u��6��i�E� 1���d�穊�DQai�Au��IoRt��n�%f�9K_�c���"�����h:q��f����P�c����7D�67��=/b�I<��=$g�9��겋'��2�--��H�F��?�y�G?���CX�
�7�?��T��NFB��?��*����`���$ɡ^1��b��G3z��4������͑��~���<������X���R J�!�����~�;1��y4/[+���T���Pѐ�H����&���4��j�����G�S��b.^E綞�ݢ���1���&�X]�䞸�\�Ab���3��OV�B��}��tb6�TLml���톈b���T���3!��#�&�	j�2Q�f�����pV"?d���bgH��5��i鮥����Ȃ�+�@�O����e��P/ X�����~���ڨ�p?8��|M��� ���D���#�c�O��@�_#8v~�!�e�춀Ł���;��k�Z�U�N}����B����,���?@�u�^�|x�N1�����۫[ Z4u�k\���ߝ��Bά�r�CwH3�jY+ȡ^�|iw\��dsF�Kt� 8Q�s]7�O�B����hA>z�w����R�U�1�d1S�̘���aȚ=Ϭ����y�Y����5�voW�C���k�^� ��ዃ(��Q'�k��S|i��U��1��x��S�L��Z�ϻ�o2�t!�[����C��$�	�⑸f+֊>���a{����`R��cC�l�kd�Wl� `�/�$�9��K@�tݥ��xh$΁0���RF��{�'p ��vb�t5�,D��T�X���~o��sh/~��9����r���E�߅
��J����OY9�����6�9~`A؟O�;M_U���mJ��kt�~T��v �)C ��r|�������Y�F���W �;�fhؐ����&mo�T�Ё�,�!����ؙClm)\W�=����)4�$�nJ�Ș�w�#a(z���?ѱ�#��t�q��皒������+V����E|k&��y���,���d5�����l�C9��&$	���`~c�U%�Wɜ~*1�Ӡw�|�o�y*�5e�z�+_���I+̲��*.�L��tT�`4�	���?f����X�n�q�!Qk�qy� B��L�=W��g�V��5��~�d���d2}�{��]!R�t�O =����I9^�/��@!��%�̃E�Gx�Žю֩�`~=e�&(nN�g2_vc���`�r�3�c}���Ka���.��2�����«ѷ�!�9M��S�b7$����x��Y�`��7��`�5��`S.	�m���c)���`9�8�n�>��ɲ�nF�h�y�;f�s�qê�0��g�v��|�F6O؂�y6��J��O���_6�
�+��XX�>�;}�_[�;��-j�~��PK���>=�Z\\v��M�>6�HR�BBw1S��)Q��>���p�	��N�q���Yr�����F����,4�5vΫ�}DQ���0ح��6i���	[D�p������y5����y)�B��4D#`%X�H�����k@f8�?��}�x�C�,�x��@�����؜�˽n��Xg��-ۧ@j�\�^V�+�����P���x��\T��.?�+��I�wzOˮ�=iO]'%j>�Y����]� E�SpP��A���)6��\�]�D��.Z<]�G����^�3ncg4������|9}��"��+�;��~Ks O������͗?f"�`����ߠk]V��N���Î, r��	?F�x�]���[�ѫ�ׅǮ��$��h�w<y��7�Ga2(�<I��y*�L�i�S�ih�-"�L�S�y���nK�߂�c���c�0q��+�@$ÏDD�\,7�1ø��h�KA�S���\p,~�+]���i��ڶ��n�ܰ���u{s��X��e�y�c���a����T�?^��/s�J��g����"�ѿ�h���Y#��o�Z�֋���j��G��Y�ɲ��\���ƞ���x��(��l�vZ���.�I�����%"�	j����UGפN��}=���I}Y�$��(�?����	��u�K��>��HU�����Zt������)�j�ݬR�nY����)l�a�,�}�F�m*!���Vf�M���ﵷ��?k� Tw3�!�nrg`��o��R�\��+��u�-�Nx�����<Ye! '$;fk��ɷ��ԕݘ�s�׏�-ڶLh�Γ��-����OoQY�:Ç[��q�����-��d�#ʬ�9���r�zڤ �{�{������N����L�q����;u�6�� #�Z,�fwa�N�M�>؞ۇ�Ӕza39@e��'I˒d��/V�� �|�	�	�Ίy�fƬ�>8	qGl�Mpaɾ��OO��������	��as�7G߂�؜(��B�o��  �MDp��$��u$e������I8u{?eEb}o �e���R�<~�8�$��ZA������rB�����wu�u#�v�q����}Â����^m�A���S�[mk�9�i��Y��j��������]^�H
�u��D�����35_� ��&K��d��d�T/������z8�0��<��+�u�<�r^��
e	`����_YgCg4kk{��J~��z���~��)�9���9�xy����F�Y��i�<��M�Z|����y��Q�5�?�糷��R��<��� ��F/Vs'~ˋn�օ�ԯ�z��l �OE��-T�D!=sd�,vu�g/�v&�4 �:q���]�������\^��嗎�%�*Yy�w�l.�����X锄�2��C~�,g]�����<�+ˈˉ�Y'��ؔ�湹Jd���>��e��*ANR(��4*^TP��9ܱDT�!�Z��o��jW�9
|�
�Q�n�%P�o��Qo}n!�&dB�Oԉ>�-����0ȷ��bG��|?�^��O��=D�T
J�O�T����2�e��j;<M-�D�=�B����/�9�w1l/�
�C�CScIt� :���4Y����̍�f�M��疔1��ú���~�#`�ZV� �	aH��(.��'lK��S����О��|p��Tꂫ���A=�e�g�<���+��k�=����0Է8j^8~�<��P 9�~�X"��n���8� ��(��89h�<��dbRSs�|hp_�*�ܸ��[k�mђ�;~�c�0���,i��or��(�̫��Yŵ�����ǳ��e=eƱ�D���K�IF��w*���BkSb����)d7�ʜ�>����%�l��ԅzA���j�\/�9�k(/+��-�\��;��4g<�v�,g$?���!_VF�g�'��ï�UK�n[��JNn;g�K���c��a�ϯ�W�4��2T%�6��4�}�Z����!�$�
5m/���U4E����t�eC:�C)�����@8-�r�A��.�U�ۍ�P�lx��2��ܩ}R���?��P����뉕";
����9�a��������������"��4��TJ�l˰5Ӵ��9E}�:�y/�b�U�3D(�m�����_Z��xN�r�޽<�#��58�8J��V�ED!b`g���pIm�6y��S�Θ4,�B�:����׽�&b��ChV�,q�2�8#s�E7�S9RL<����!HWS�SN�2�U����R��l�@(8��IV�vݒݍ�S��_s��Ɲ����w��i( Z�-<�>u������q,�<5Ђ�6�������`�P��;��L�x�#��bf5��U&'�8����@���+�#���i�C~�ጕ������0-��l���Ɣlݵ*B����=�W�x*>��<G������8o�	f:vTlN]�Ey> ��ﯠj�'S�5+��/gU#�o��2+�]Z���qX/���`�[��%XW`M��=h5�
������L;2��쩛��̼{З)���Z�x��	'�%���Ӂn�z�q������x��}�����^��-��"��`{Z�)�U]V-5�\,���xBOHvMJK�v!M(X�$bL��xC3�@��:>.�������CΞ��\��]�U����][_���/���`,��hx��ut����$T+Bd8o����^�]�_�R�7����Y��'[.�����每��
��|I���9kY��P4�b\�)Db���WRT(j_~�zi�(����3�jV��=���8^�"O�!s�ͼ��c�K(��7uX0X��t���>����X�K�iϠ��>�р]��Ni'�����C&�A¨`�����?E�9Ȋ�@ ǿ0�	������i�2�v����Ny�B�4���������X��5.�fd �Ob�[�*^����^1�:�>h���l�ލ�5�r�}O	i�6��	$�Mi}/�E.�2�<�0Q�m�/��-_���?�D\8��[Π���}h1��4	OGB�@vi,��N7S�ƏK9	V;�z��H�{x���m|���H�mz߉O�Wv���(��{�B����F�� ]����Z�&h9)�Q�%�a�ƨ��;�,i�N�%mz}>�,C�C���V؋�)��k�)S���$�V�P\6��`�����P�y��G�l�S٘O!�!B~B"
��>t�k�C��T$!ɷ�O��)�2�񆃔�j� wBRD�~x�b� �q�^�zdf3�Y̐@�k�h¢�W���zJ`��+7L�!B)���zݎNd�U�M�"��@��1	�""�����ho�@��'<hw�Gfو�q����z����O��l=���H�BT��/=����d]���I���߯��)Q��T1�MY�3<�{�5�wA��?֭�Gυ�,�
Qo	?��:��v�;�6�+`xvZ��L�眣$��=�l��¥p�q�U:k����^�;W1j����)`O�k�i4u��ot"{9�K�9��@�g�O��tS�W@E��ʯ��T[��HV��_>��z���p��m���z��H�����jxYNgnws<�B���`�ʪU�P0�E��镣���%1�.�IG��|~9�y|�R�o��5/��?.�q�����A��Q�WQ˃����9���v[Y�iJ��8_t>Ǐt�
z�,@��sg���?y�ވ��-������6\i���dAm�U&�Þ����|]�(�t)�@;x���g���:�@���,@.�('G
�T���4"-�^ �P�����\���2A1&x6^��i�љ�|�����yp�Oj7��<؝�3Eu]A��h5���x����j���������i~����len��I����F�T�I��mj
j\1��VK�L��QR�<Y��P9����6�� �9�����w*����'���&x]�m^și�}�LU��ܴm�p<z�[�azP[�����uTS9şL,�dF����s�nF�t.�����3"\���귨AJ����;�ޢ�L�h�Z�)�Ms`t�p<9 ���N(��r嚦�n	�K°�p��r��きs^��{��;~��K��ojg߆=_���[�O���l$��@G=���!yepv��J�	t��Q�*�F����3;���2	@�Q�̟��A�Ӥ_$?���=���X:�i)Cl�rV�9@Oi%x+��ԇ������~C'��(�P���(��[@8ng�a����7������d��u(�o����}���8�����X��d<�J��{v��oF{����`A;</�I�U���p�:�wc��T�f�/��}����0�@n�ZPA�{��.Mً�̄�.b|B@�9��� ?:R��ݬо�L��y蜯�m�A�@�`��Z�3=�0N�f*��J�{"���xOQ"�D��۰�l�6�|( �k2�s{�f��N^e�0=�������iN�kk�*���;M���N,�2[����'kkj	6_�Ü~�PP��FI���ӟ����g���#��<J>N'M��~+h!i݅��vs�q+�q�����C	�J��㗘	�&?�LL����[Z�Ԏ�p+p-�SD�y� ��~+���fu���&P3&$�x� ���yr�~|TSΊ�S:�9�73`�D]�so�].({�!Oj���ju����|f�jV���h�|c\q��;cV��PWپ���J��D�wT�6�B|��/��w���܄�|�Yg���^$F��N3��i����El�d��/�4�?��ƴgN�
h���t�� �iZm�+!�x���{��!*̬��H#��{���ugxN���fk���O<�@(��5f۩3k���y�O��Y\�²��]iY9˄L�W�*3���H2��6��c����,-#����bn���Y�c��[�|��p)��B�S��`-	9&�ʡ���u����t��i�O�|�)��L�D�0j��|*�c0�jyXR�P΍�1�(-D"h/v9�,D*J#a�fD|��*2y�>i�8X*J�Jz�tfbs���W�m<}S�$eT����0UuL�2Qn/I�Fa���X��#`�J2�wX�B�ɺ���Tb�bA�tɺ�3��![V�����P��kmbg��~������Y/�'�n�����Ǒd��62tCz��u]����geܴ������{)�^�_�4�AX�]f��U)�H�!�f�\�����2� ��H�y�I)���od�K��7�4
�f��q����#p���/����u��56����Q��2���&ʓD�oT�vj-�ok��Q���N�j"LOd�HG��0Wl$�(ei�� � ���C�1��I/C����Y_'(*L��C1f�=�e��nЅ�
� _�u�#I?�Ϙ*����q�_!�]����M`�)�[C(��(;3�49Jy��5{z��tn[�e]:YE(w�E��ӄ=8�,'�V��S�*�O����5ۤ;�G6ک ���o����Fh��]*�D'g��y+�*�g��b��t�+��3K�@������{f+�*��V�� �dlh� 	���h,���?)歞/1%7,��;���W�s��j���!!x58d�9�Y�s���Y�+�M�P��&lZ��k��|��_� ����t�=m}�x�Z�~/B� R
8��Z 	/�Lif��&���$}T� ����I�	�>�h����]X�9���n'YnA1[�|2\�kx�NN[���1���P�k��O��TB��l���E�Z�	��^AA5�/�h���������PCŀ��P���#�v!�-YQ;jF�661�>�^7 ��s�BA0����)dہ�]�!�R�A��2]~!�2��=��	��VU��_�2�0.�'�s��fg�5�d�hXs ����&��a���0.N�i&�'>�#Vp�E�|���4[�	�5�*ci�h<l�!��r�дdgf��3��	Y�@n�[OK�͡��i���p�f�e��;�e�/=�r��F�ӝ����/]�gI�Ȯ�w&�Wl�C�(� �%�"�9���wT��YG��62����_��#��(�>R��e-+3`�ԙ?q�#-��R�j�w�`Ӹ��������0�Ajz73AO�XW�N˾m�y  �����d�g����E0�>�di��?q�e�j�ÿ�18*߅�
������	�o/q
w��v�?�mpf� �E�R��'�?e����l�xQ�w�3b
<U � �$��2Q�zY9d
[��X��,�l�b&~����Q@��HEb����+t��_��2ī�@5/���A4	����y�<��ȳ�k��%g �,�Xw�M�zş���nVo���6]�Yh�P0�hI��4t�w����֊��͛Ƹ���L�?��orO�,��HO�z���ɋV�j�L�ل��r�t�2D�q�]>s'M��GJ\��$^��xk*���Y��/��:�?���W!O�sMhX�W�[�����'����"+[~���j�S�]�E@���l,��f��(�r������@ȭ6� ��L�)�V���M��`d�W� h,��xB׺i�^;z���UѴ�s�5�r@����Q��.P�U��Ny|�8p�~"9�U��a�#�� CoE��� �Bv�:���[�ZHG�!���n�����)�m�Fk�!G�w��)��b�8��0�?;�?X:Ȫ��ݑh�:�}�PR���v.CdC+e�M�-�B:�%�l\��VM�v�_��M�Ɗ ��\@�c��BbUu6�,b�&IP=&���0S0��7{\Z�ΟC#�ǯ�}Mu1�"��(�Y@����#�0�Jzc��y�J;�ĥ:��f�@Hօ{U;�(:y֝̂�/�#Gǥ2GT����q@T0�4@�
���PM��2�q
��)z��

��61[4��V�et�G�Wmu���� Z��j����4^H��h2w>�� @c��1�aS�k���e;J���<?�3�	1r�4�%�-t"!�J��l��g�uBn��a'ݫm��AkY��K�,�@p��m��dN��6g�s&�f�]��[�O�m�C+��aƾZ���g�ſ�\���p�p�Q��4����s|[�L�)}6W �?4���I|B.����}���d�
[Z�9��j��m�fQ����Xo�'h5|�Z�x�\�X4�d��K����VŜۼ��P��fH�e=�sҳ�0�k��A�p�d,U�
~�"²��p��c[(Hf���iՓv�l��Q��7��[�07�#��:\�K�-�W���
��\aZ|3zC��55zZ����N�W �K����3� 8�c��o,#�=V�d�OmVl__=�n���d�
r}t�h�X8������8U���.`/̡ �X�v�\6<t����br���#(N�%�����V�Yy���ݵW�=vNSͶ��֩����	ȳ9a]U�h� jv��C�W#�u@Z�.�Ϟ����x��ڦf\{g�=��1�f/�39S���Y�((��P���TJ%����h��3��n�W�4�����N��U�Q�xa1�&0���?r��j����W9s��"i��kW��W:�)M������FQ�>}�Xh��"߉���O�S��5l����۝\  ��os��"t�B�#B45�Ƨ$t�Y��~���	^�%��螀�7z���)_�[���}"�o�,��=��S�\�����3�_����h�� ({������'�nM:w�����9�f���@��C�X�$钪8q�X�d���)���;����_��K������WH�}�(q�B�K�̋f��U�z�,�:�}��`,�ڐsᮻA樁p�EH�5G>�-�=�\A�n�I�x-�xT+�X��\ֹ{����g���H��~��V��cе'��j� 32L��N5W]�����F~�Si3�{�+s݊���f� 8N����i�Í����c)`�J���/^�J�tvZ3�b�M#�7�,�.lU�|��"ؗ���Ѿ0�L����K������a�J�f��Υ%؀����W8pCl:Kǻ>!�S#H���}�BC�c�ܲ�U��(A �o�p��(5�1Q��]y�S�>A�(y`Lj���w5�Dk=`���h���q�K�1���(�$�T�v��뒢�͛3��~�f��e��Ǻ/�`&��U��F߀8$��1��,��pHS��)ڌ��41b\#%I�4����Gn��(���\��2<1��g�iL�P��Zni��H��J1F�'�R V��xu{�R�����%J?�����95׷�Q齣Ϻ�R��]���Ơ8 ����m�����;"%����G�[��La�͙/r�+�ׂ-��A��[j����!��Z��BdKQ�������p
'�+*�q߀A�rl��g� �b��~-�8R�;�q�b�7��9%��b(3~o#�>˦���
�W�X*�}�ږ�w�m(_�
4[
sV\�:��2y���4{&�b:(5roT�B@�;twkV��|��N��&QyB��5�����Be�2-bHՙ�{�&�s�Xq�]:���ŧ���%�f'Sޤ��8�(���I<���t}�?U���W-�T|D|���d�<�6�Q<_�H`�tu)��W�$���U�^B�c���r�0�}��$�mYX�~�<�↲l2�Y^5oo	a���]�6���a�e�N�o����6�.c}I�г�D�N���?r�����/�t!E�`Q�v%��zD�_l�;^)HS�7e���i؁�2r��7��ӊ}���I*e"ο9�)�\sܟ�C �S1�(���f�-�wʉ@��By�Չ�hh�wt6H[��
�d-��ý��>���z��a��^�}�����f�!Ff&�Lw�]��c:��c!��`�B��FI�U���|�27�|�Q8��j�i�~kPT1���<�lח\�ܭ*���u7�l�7�=��I��W�n����Ɔe1�:C�0������f'�Nyb@@˺��f��.���o>u-;|Ǧf���DA���
� W�?3�|	@���ۃL�*�"@~�6J-_�!u��6��H�=��DB�,�&��f)��A�_��-�6�%mU ��0�|r��^�?rxJ��K�W������Ǧ�.^?�jᔺ	�ӌާX�<���d�}/� �K�ރ��B����� �iq�Lo�n�=H��#@Y��#;~��u����Y8�Q�c��N �Xz�x�$�V$�Ƕ^��������|���t:�1d�1��H̮�;b�d�ߚJ��q�"���Yl.ܠ���6�I���Й	]�+�k��P��ou�� ��xY`^������QA�l�u�a��`�YOI��T��y��<A�b��t�@���q�Q�]�ǫ$��m���C�	4��$u!	��z��st�F�g�H�k�/�&����IP ��
ԛA)�h��jb���3`>� ��0a��Bv���|�g�z���2�i��#��v���Ţ��d %1�:�gC��L��cc�"���*[j9�� �u=���6; z�����՗-|��M�ǌ(j�=��]�����V3P�(��9�jT��ģȣ6�"���^�UEP����FT��/ͱvt��I�����n�(�SN�W$�М�'��Z��5�M�:�>�Ì�J'ܐ�@\�0"��6]l�RE^t8C�y$�:�� ��r����G�ó`ootȂ�%-�܃d��(	hN�����E��$Z��9"O��; _�Ʈe��YF�Ao0J�+���������mJ6�AD�G�ΐ�B}�AI�ݏ��s��4v4��5�����<pl�Ӿ=�f����т��+�8FM<-{�>�|�>b9rI!gKAֈ�s{�����3���(�������(����nm\�sGT�'d ����gB����I\���|뢇�?�oYW���p�$��O�8��E'�%ɍqI2�sQ3�.T&~4�ȳ2�A���{���Ԁge�EA�#0��(M��y4����|���,��G�
��_)���P:�E�A鈶IQ�= };q��,�84s$��O3�4�e	� ��	(�~��:����ܜdZ�g�/��j����C-�XE��������no�H��'��M�e��q��3����C,�`I�0+r��� [Y3AF��g�z�,��:d7Y��]U6�i� ��~ԷA
>�pF�\;��j��;�c�����:O�q�]��M�1�4��29��wZ��Z,䆠��S�7,�r�ډvn]�35��hE?r���2!��~��D�����A�>�nOƕ�>}�����Ҩ%%G�1߿�� /{����p���)a]�P�߲�ґ㖶��Kʹ�ƩW%ܨ;%�L�P��ͫ\���xCP���t<"��o2�~~$^���m$�1V
�6��r1�jOy�Y���u u���'��|�}�9��chU+�����خ���GH�����C�����~�,���Wˢ����<�!!���[]��!����:)���Jʱ�<������<Әwk�6h��x1�*��"���T��mO�X��-G;z-�g�4���?��Qk	.	F��Y���_�-7��}����#�il��M����~����"�mƻ�<(:u�o��=�	�fCpM���Ԝ���ǈ\�g@�cǺ�4�JG����_�PA���&���%�a�`,��M�qj��$.w�}�i�����i�V�ծ��.�p�Scڳ]?p��p4H�sџG���VY�4�nm��Ti��[�ty�cL���1V���=}^�{���!l�w�]�#������HRό�����ISq��	t@�D��9p�E�9Y�����S�3�m�&9�{�Q�D6�IȆ�4t��������-�f�Y{��]1�%9l���}����mm����¼�"u��ϧz}2F[��<4�����Ok�rm��~)�2Si���~��["o�m�����܁�s7��S�k�ٕ��nk5i^��5��y�[��%ҳa
ܮ��hT�]��v�L�?R��7U�@����̊	��S�!��y�1��`�=��F�����6zQSl2��U�58��L�'�8�x9��Q.aX�����!�
c�C��J]z��U/�$�@�ok���ș6�
Va{3� b�Ï���d��`0�R�K��Q�����`��z�ؿGii�ʚI�|���T?S��[�� :��B�h��m��zeMa	\�c�uf)����m4ȧ����B�"��1K"�;� �w����,�������K���b���/wR��u �Ȝ=��J���I���!��k����r�
� Sm��,�l�@���ϙJ1U�N����QT����8�+[��mu�N�X�	Ƚ��(6j�vLK+��%�����l���c�u@0ߌL!@�B��4�܀�C�efjR騋	m&����\�Qgׁ����D\�(��x�iCm�#�|�O႒�κ2 ���l��[� �K^�M��W/��+7o���Ūn�X�����"Hꢪ8@���'�w6���&�ɈR0������ˠ_��}��4��L@H9O-��2�ꗭ��
��(k��1�[1�Cӷ[a#P8^���
�U]j�e��/����tv穖p�6��3#�qS��%]y�
1���G�BgI@��Xs�qP_c�'���iK�L��*� 6��#b�?�2d���8f���G���Ab��n�`�!��[�r[�Qg]{u�������w�1���Ԃ{�� odt���r)Ց5��OmD���{94�}�м���f+[�
|?"'�hCZu������Ֆڨ��t�j}����� �ɡ���o��V{ �Fl��Z�U*y_O�{tŁ�?��V�N�}�9i���W�R��E���oHNX�߬�G��5M�(������M/�ԒI�_u��u; ��>�q\��X�'��4���u
�H��FSI���^�Q'�����~T"ʅ���'���-"N#ѽ��Շ�'�:Tz��ahs�xv��N���:�������A��9��1���KU[�J�6��7$��ۋz�����й�`�R��ƿ�y#׷�?��|��F�)�*P����s�jw�a5LR�UƦ^�"zyrӃuUTY������ǖvHC9����0��)��C�U��K�Sa�>�X�Hop�j�U�����i%m���L��J�/UK�ɩ��\��V�dΎ�ˁ�{��<)|�FCfDjcXmSrm�T2�*��T�z�x��b�$�i��̎d����?$����)�OR��ݎ��n�� !FM5���>D�r�����\��[�W��(t��H��?%�Z����|�_����VA;��eH�QX����-h�<�y�;����Zp���rٚ�[�T_#^p���,���4a�L�ީ����6#W�f�G����ô�'e�>Okѩ���֐z�߰�hl*����������5UD�<߂��C��ȚS�N�{�ǜ"]�8�ͪ��Z�tz	����p�!����$Y���MsH�w���YȖk����/W�jOC6璍»����PO3�Q���]P�1�1�팖p�yK����o�O�w��n�~��n�"�Y�O�F$@zd��y��kO�_��^M�В<�C��ӏ��r֋q��'*vP$`�� �� ������B�su�J����ҿ��;��Α%/)��?Qɟ��QM�~K1�.D��a�:�t��5��I�����L����e�mO���N�@��B~�v.�d�T<�Rԛ�V�pA���Y��t,At5s�k0*�_��1��2�`I����*�B4�ҩF�������*�sZy�ʷ��.�p��Fx��U6+K�x��\)�$׿�����؁����ۍ!+~��lr�ySn��˽2���]k�s��>��BeU�iD7��H��%W��H8x�W����苾'��{���x&���.��m�S�
H����}0�_�ɄlH���tǾ��q{���%�(�%��뢆��;�v�u�Gm�@�h�����,�j�%
`�6�5��g"���e6�>�&2�Z{��#�eC�ꝯΟ���h�Ч����U猔�0߮���~�>�a@=Z�%�}z7���z��A#�ۚf�Ə��@(�0�
|]����l��{��l��1i3�E��j�L�'�l�o�Q�?1iz�Z��Dg��0Ć4��W	��m+��C,�S�郁;-(2=_�D�5���	
+����AO���4�n7w)y&�S�3�7Ze�Vm�h�.�kpq�K�A�R���߬ӹM`���[|A��P�R�;f
c���yẼپ� 0���B�5�8�/1]���F�7�h@�� x�{��Tk��@&�X.����ߵ�Q�!	N��U1��ǚ�� �(Rc�P�~|�Q'��۶D�����R<��|P��/r;���)�^���'�3�f/T3������Zװ�-4A�ϻY4v6�!H3Y�:ҷ�A�Ks~��yt��n��:�0��U9@K�d��ZŖ�\�Z���8)*�`V,Ԣax@7��g�͔�f�I��ƅ�q��������v�d�I��1U�Zէ�&Y��1 1���i%+��Y��a�ӌ�9��BQłGQ�֎�,�om��9��"�u<����)y �r0uK�vz�e=���_��k�>��v �D����6?������y�U�A����ź����v�>|�
��ᮓJSܞ#|��߬���Tg�|뒉/�I^�J0��<����KR"XK�+ڬ��	s�*r��c�)������s�Om�9�D���2���j�R!d93�\����N��7q;��dC�=ށ�~;��� :y�G@P�X]"�&u G���ȝţ �X��Mc�%D��Ŀ>��B�(�*�B���N� �kRd�ͲB*�V���ԛad���AD{d2��SR]S4�~V�K���w���$�^�h�WH��x<l�V��_�QY��J܅�����~���s�Sξ_�����Nz��)��=�|���_�~��H���xMp�O���|$�KJG�=��.d�[��2d��^��\P�?-�@�P�o��'k�u��7�pSpo�1��4f�c�Pc��Ɛ5�Ʋ�;��r���k�>�2�d�=F��1�{���=.�fnf =�ҏ��yW��t�u]?
��"@ͩM����4O`!m�ꐼѺ.)�	_�9��K'� ��oδ�����qU�<N���-x7�&�o&΄� ����Y?/џ&�x���M�И�lq0�heg�.s+�7#C��|�hV�v�`>��9}��l
��y��$+���۹zW;ԋHy�FޣO&a���= ��:���C{N�Y�E���@g]�El� ��c$N;�\ 
)z
�U"��Vҝ�$Y�M�d�~V�Z56jim�TNz�̝����y�1�i֠���~�BM�r��?�ZgG@��fH���@R�*��<��vy	2c��@+.��y&�H
b%_o5���d�&Ƌ{*�׮���
�*��z+&��0����q^��A���!C�$��x󱼐��.m�,�SԚ_A�;b�鷲���	Ӹ����Ч�2lg:�2�礜@V��{:����?ǌ]�&?nWߨdnq�-)��8qE�=��.j"�S݄�V��so:����O��x�zF�~�R�};մ�1;�L(��>�������C$D�@t�Rƴ��S� ӬӄFd N����y'�J�'u)2��%=D�'ڋ��&��������0�{E��3��N\�j�,d��/�5�;��<:vM��ϫrE"]��I���uo��u��O�\!z&�� �2�N-�jD���u �\ύʸ�Q�:Q�S*����1��P6-1Z�w���Sb�!�k�R!���au:�����1��(��G��G�3��/�x�C�H,c"����IW�سI-������:�w�.��<sу�Gܼw�^7����Y4��q>����QGvi�_~פ�W6f[���w,3��m-�jg���]�h�c�ZX��d��#�-N8���X
�jV I�X������o�S���6U�y[��0$�����1-����<�����q�S��s��SAIμ����|���"|�<s���8�P�/���H.�\�xf��T��6��l���_�I&&r��u�s}N0�LH=k�U�(%󐷴�_���xp��4�ҿ(��	�[�U+J{ヾJ�|ah��� ��*��X�ӓ���1��]��q��!_���O�D���~�فhP�
��\��j�)<&.�MӼ�Nf��[V�鑦�J��*PN��b��qYx�>s�ʠi�c3}>����z�߲6w�����y��s�3�O�2�N���$�kU��+9�N����!i��bAU6>1�.�Xy�4yO���=8&�l�]QJ��p�oIާW�@U�D�Բe[ښ�T��Ԍ����3BP���,�r�%��ZWZh�����* ��J�p[`�LRe{݂�jen|�`H�[�q�!e���+�'�@9��w*5JR�ɑ1��w��RY��������ɵ!����oD�򯲆���/�׾�Lִ��4q3�[)�|k�=���� ���Ae�c��m�C�݀y i�d�
'��%K��5�.� <0�~��Y=#{ƮYe3@�q��j�[.2�j��N�s/�k@��du&�ꘑ�hՒYd�_����8���xY'�		�4zϟvF�sAA\o�ᢛ� i��tKX6h��2�hsI\��>�I?����ܶ~�7��<�c��\K�ë!5�
F짹�y�\�Un'ۧ��rI���\n��+���l��{�3�d�1Q�J���O�G�M�5�6�ǐ<Z9N+)zs�܋QM��)h�U�,�"���s�:[����`��,h���hZ��%b�ϓ�+�KNf�R\9���Y˺P.)���Q�Nǣ�v�2 �sU[��������Z�nA�0����Yh1GqEX�ĝ�g�"G	��D3dT��pqX�i�������^��V	�=B���ǣci����T{�F0 l�R��d��C D��p8Kcf�����f���Q�c��p�� Vn{���i�����M�P
�Z�K�c�ʩC��s���#�]��z�}Q&�3E��p���-�Y	?�ڳ������凊ޔ���K�y׹��4�zIy�?�5�M|#bh]������VT��o�.�9�HfM�̗M;����`g�f,-]G���IC�M03:5[]XX�����Bz�h��3�Ɩ$���RW���<�&�a�M�ٟڇY��-G��*g�}�w j��m��x�S]�ˢy�VO�
v�Sg}D.���U��L�c$Bs�������/�%-q)��,�EV8��Wd5S'M�ee�O{�%Ohy��\��v���2�ޫSZ�ѡ��C)�	��d�m����`�C��S{��h9+�]��7��B�zgG>Yl7�>��eqK��$����ї5�,������+����iM�e�0�n�O�|Qa��<mB���If�A�B��	�:��@��{����P�˸��ϔ�Y�s��|���8�9g�4��F��M����>�9l��}�i��o%p$A�C�˔S�_��ȻƼĮ�)�ۍ�����Ȅ��Ccq��
��F$��EyS^�1�4}��8==`j�|q�N�U�s.VK(��Lm��O�@yy�1MG��;g0��)�m\����
+���iE}|�/���lO���h�|(��q��`��$&&��e�K�=�^M�!C�;v	=Ա)�1�K 3:��O��qSC�%
��
' :5}��▇^�*�NT
}����R#� �����\����O/rM�<�h3���Eu�w�k���C`�54��9��Z�ÖGO�.��R=z��U�41v�� �5�is���[������~g��BQ��Nߜ&:�)�_eԯִͤ�I:W�+�ʦ�.�)����W��	�m��R���'%�R���d]��C_;O������X��+�W��2hn��n�?�g>QF &�9�[��;��e�E�(��2%�L�-�Ŷд'��h�JƂf�>Aư�#�.�=�[��cR�݈�]r���2��&�.���@hjr�s�`���aP��&�"�y�sn("5ZSiT"*(}�Pl���y����Jz�#i�
���P���&W�
�eC�ǡ � qա���ɪ �r*~47/��{";�>��n�x��U�B��og��O=�h�
�R`QD���b�/��#H.��Y�,��z�����I(\����a1R� �n�iC�L����A�^x��������@ ��:<49DP=tlLf/�7z�́<���^������z���/�����5�K���@:�V�=����5K��?�6M�O���ʂ�|H�jn�����T���B~oL�(������$Mt`M[J t�h��v�y�g�A�+�]B� �����=~�P&(2R�U��T'n�Z�	��5�7�B���^�wVv��ZԋR����
O.~��lv$�7���q?#2�����/Fk@�]R��Z�ŵ_��y��,}��ax�n  r�0$}�C�tu21A��w�.z󏓺yX�s��G��N=Q�z=_�Y;!�V�V�G؅�^V<5���Sǉj�f�_��qaAR�Ѩ�E���z��̫	6� ��Zp4\LK�q�Y�vt;�MD����&�[#s�s�lg�M|����"Z�s�F�����[���aZMJ���9,\�T�`(����$�f,��8u��&�IVag��S�`�@�iCx�\?��Pa�t�ڦ�KjP�3�'�z;�3�}*��љ���Nm)�a>ߛ�FEnЩc�S� Е���#N��¯JC��o��1w�8�?�2��T�%��+u�d�� �Hbˆ��&F�e��� �e�n������im�v�bTr��I��uܓ��;ǡ�s��zƲ�.�.���	p_�˘M���COH��t�8��t��!���~h��qm��r�9{Q�N���vÔ��Ù�q��(Ρ���pj�;�$�m��K�8j�����Gn�TNGXr��]?���S|�W5Z*�pN�B$�.�qk{��\�m	ڊ�!ѷ��3]����v@9���zVZ��WZ��� ��jU�fQi��&-.��P54k�`�X +Z���vy�I�?Ɂ,�]��˼�,�f֫
H�q����uT�+���q�A�)5޹7K$ܲ�,�8�f�f�-����b���E�t2Q\O��H�T�;LE:����8��s@��苮�/$��5�]���֢/tv![0����P���[�t;Zo����2@C�D"b��'6�<�Q�[� #���禛���ʘe���7	�yL�R\�kG���H���G&"6Bab鋭y����X͏c���p%���!;s�/۫	�p��b%�M��!rQ;	2y����VA{*�3��,KWDDd!�/i��G�'��5,8a	4������ ��5��؈�-�%���RW$O-A���5�� ��W�<���9��vȯ�q��K����t8X��ri�ͳ��)�`��Y�D}Q�������v��#ܒG�bF�.S�W�+.�����TK7���I����C��~�5S�}av��b��[-����6�KPLgv���DX{8�OjP}c�i��z�
�����l
����m�[�	W�fB�������>��y�B�, 9 &{��Ã�>�n���vj��a�n�j[�*UR�x��	,D���L�����H����&��`Î�i�b_՝�+�]���cf���u��:���u(�͈��*�:��5y�_�3f�Lf�<խ�l��c5���c	os�E�C�_�r�t^UY�0�f5qy%p���֞��9�YV����H�^����a rw���M�y/�P0�^2R-NZ%�:^ '�2��z3�VO��11�)0]:�!)2q��ho�!x�,%�z�8f�b#_炘�D���c:�.�?^�_;����,Y2�xf<|�Y�N��"�
��;�Z��ٴ��;dH�d��5I�R�*T������^Q����D��%e ��mh��V��س�t[r4��ݷr���	f��^$�طD���s|7��|�*} �VUA�-��h +��Q���Ns��\pˉ�
(h�Ĥk�V=�����~�*�5��	��\�k�ߙ�(����)�N��~�ǞogɶO���ľ�C��['Ӎ�^ �W�&�qd���p��Z;C����o;�0�����ҍ�ܝ�X��E\�,DP2�4�*)Uė7?{�Ŗ�^;d���^jΡ/�?�9�;����� �e3X�����ё9蠺���dYm�B8�ϭI*B�3�~ڼ+�������	�A.z�T9��#Q����y=V�}�9JrkC�G��1���R�����fu�%[W�q����,)�iK0=�1[��+�k�f���DH��Q�_��lO۞e֥`]/�t��Qp�4����d�<6R`��F�ZYyƵ�3o����H�y��������{�I<"7
�ˁ�S�3���#]]��>H	�k3>�P�o�N�e�h���"�VJ��n	��2r�iD�j�P��*F�x`=FP�1����[�8�8X�├"38ƽZ,���H�&���䏻�"NtM�K����0v��g���s�/_6o��!��	z&�� o�+�t�'�^2��I��+�YK���Lݱ��@;c�mW��̵����ԓLe[���J
.=���u�D6��<�p6�O],���s�D���)���<��r4-k��Ih�oJ���M��Rk�o�S�*`/F�
����#���X~�.�N����Cj�?T������׏h�&��<�9'o��l%��N0U=�O9?�	3��v$=?��5���M�38�S�Ec�����B��t*E��g�D>t�!��Ӗ�ؐX55�BPɣ+,�����Jvp�=��}1�� ŖG�8�0�ߜ��֥I>s]�D��\�}H��wF�ڞϓy�4�؎�]ӛ������B��*������A�ņ�zt(dyo)�j�2^J ���P��������g�l�#�`�\�v�Yn�)�|ѡ�(���D̆p�MGVb���FGa��횰t�i�nGJ�k���ڄ��\o���܁��{�馅�=9e����H&1g�N�t�$�0��=t� �LZg�}�wr��b&��feĽ�7غ��\����D^��2�a�+h*��d�4��9�����,\)���ơg��*֕I~��H-Kٗ�3xި%��A�`9*�.�:���/0<�.�*>�؛�X?�����1�SO������ø3�V��h\|���ts�_�0�7��P<�ְs�å�p��߀�8���6����p�;�t��d���̽�H	So9��$��+'��[eYŷ?Ǿ�lU��B$��b�qIQ��z�g��:��f+��4����P�E���Ó)I��g��	��ܯ��(��.pw����m��jB��Z7\�׋^g�dncn+�̫ a�8
�(-��+�P�������Դ��]:�+ʻ�+_C<w�Q��S4�w~��}����K����s��7�c�0��~Y�j%FO3���H����d���v�n���j��Y�E{i
Δ�=��M\��C�u�,T��,^*[� ���	V'm�
�����#&hH|�'ؽ�'�޵w^l��!����6��	���@��Ƚ-�K:�cՠ�H?
�{M�-��9��4ړ�����R��_��nHݭYA]j�
0p&�'�Pj:������E�U�$\�%D�ʃ���z���EʄTi i3�[q-�T��
c
�'�)Y���xoO�3���}"����+�`I@��5�I{-&�����r��Ȝ�
7w��ӹ�=����6('ث���8-S�QYA��X>��uk�o����������|� Q����x�,�*X�u�N�q;#�tq����n
C�沶��l�,U����{�8�y�m��CJ�����F�N=B���)���Z����
Tj�E�&��o2��f�6A���4%޽������	�'���8a���cɖ(�9k �r}%pIt���
H���ձK���Uy��aHL.�KO c��ZVi��r;>l�]����)"�	�����ţ��Li���5C̊� #��	tJ\O���>F#��S�U����9�g���,��{�2C���_��Lp�6���? �ʆ�໩����� �Gŷ|�@���J�y�J��j���.���K/Nbȓ�ܡ�L��w��2}�z�v�5�_���O��i��ǒň�q��ʯ_%��s��hR��_ԘN���P��(�3��s�հf�4�0Aw��*�R��
Q6ᷳ����kn���m�,n�=�RN$6��"mmv�`�@�ֶtΟC� C�ǟ���H�>L�=N�&�/KU���&��(pV 5���a�[�>��D6�
�����Y૙���7q���~�[�;,��x��K���1��0���7
W�l/z�	�D�r:�4Fr�,
�`gAoც��Jw�w�)>Ѷ��yQ��{�@w��>r�����C(.Z�}�,$�G	2��?GW�T�����L�l�._\��o��k�Bu°"hx�i"�X=���7#U�a�7��Y/5 F���Yw��]:n��[�#ߝ���_M*�q��ގP����y���{$Q��X� #rw�+���w��C��/�wX~Z��Q3��H�8F�k��}��.E$"׼X�گ?�$��u�d�(~�m��
�K�l��G�2�*��kʱk:�WAn��#:
H4U4��|jj�; �@�
J��Hz'\��i�:���!2N≠e��\(�w�Җ	#)ziw.���M}���o^m�d��F~4�G�~/�8�	'Ч�9
�ه=$�x��!.���>��̔M"mn����J����?%GH�+��}�]#=���g�K�Hb�I�{;�t?#K����U9;�Q,�\��Z͎�G�#r^���Kp��w+D�А�9,�"ۊ�*e���"�b!2C� �4;���3g�^{��I1�('eY�F�lC6���Ii%��w,y�m�9{M����Qm��g]�"�(����j?M��w��N�@޹_hB�&z�Ph5�|s��uD�ݔD�!{k\6��v a�'{��g6G	��@�k9o��7�!
��o@i0�(mΊF)	~S��M]�fK��S���%�����b��tT^=�Ӳ����ڇ;���
�=t�*�.փ�xt�xG�D��>��Tm�����8..O?����΢:��diE�K�9ɭ���d*c��e���@� ��O1ɮ�ڞ�2��Ϣ�Z.gq4���1�ޑ�|��|�4b5?P�sJ'W��,s[�~���%j�`�ԥtb��4�3��� �NpJݷ7�eu��J[�~���Wj+�҉$��Z�Î�];M1MV���=|c�q�Ƿ�F�_���r��n��r5��lPI� ����.{Cj�3��L��eT
1��s�Hm� ]�@ �Iv��)͘�0��ga���9���zCp���C6���J�����"m�w;�)�F��+�%�s��w �0������hG�H[wB����uũ��M:Z�t��;�%�pC�T7*y�ķ�\Ɗ��
r��>~��
`�܊Y�`��G�8��Zo2������������% �s�g�>!���	p)���N��+���YmG�����N����k��E�=2�[��"դo��8v�O:(�ܭh�p�p��8n�Gr��F�*�=7���]���kx��O�X�����V�`!ŭ�����JQ��+�b�������V�yi�!�uL�i�Lt��w�I0����g���	)_��a���`��T�g��o�m�-�SP�R��"�ߓJ�a�'��r�0f��y�`P���?�3z�l��d "y_uli�f�&�4����X$��Җ��dXg�܈��}G�jK� ��� ��'�륧i���<OK]���sS�}�˘�˓=�egᅾ딮��Q����UE�9]��7�T��O\sPM)�7��N[Q��w����J�~�Ԇ��r�S�$r��y5H�'�����޵��:,��J����i��}6� �� �n'�)h��q#�(�!���г����������ϩ�Ir�����T�o@�~���$�����8�6�T�$6;|I��!3��W��L.��@>�qK4�&�)����63�3F2�IkR�w�cWH��$���_�������fc'fӟAH����j �oY��,X/C�r��,���k]�_I����O[aZ�Y��c�#��P�`�" ��q ��ô���b�R�%Pn�+w�J9\$�w�o�υuF��"��H���`��􈉠R���O�!�H�&�|qm�3�O�R܉vio4ӀcqpʗC�5�ª�������j3�hz@�uI~�&�%��(��I����D��4��H�6,4�ܯAא�}�+d�����M����Pݣm��<0 ��_{�)�ȉ�Cc�g�o�� "����?X����a�s� /�j1��;c"z��?�ivń	��,JB݀����'�)��}��eL3�~d�W��ށ����r8vU��bUb�{v~DǗo�3�31��@pD�X��t�a�w	��	N�_�����جb��[Oy_����Bn��F�:���W�P��|�?���Q�H�}�lȑ�5�-�K�$�zcӯ��\B*8�ʈ���F~q,�ē>�8�ߨ���GYz>j�#��v��WA<s�2C��%���~�E,!_z�b�A& �	d_�q >��]Ԏ�&��,$�[@�?��Q�!M<M^=Fe�vrҍ�-�H�TK�/�"�GL�F�aH���Q[�D/N����i�bhrH[��������p�>`���O�%qTS$ٖ��֥"�e��A|xS	�0��Y��p��YBJM'D�&XC2�ai.���5{NY��8���o�2�s7�D~������7���s�
`���8�t�,���Bif����^�3ǠD?4k��ަO�7�\����a�VA-|�Q�ji�-�x)F�cOSRT�`�A��P�hY��y�.L_���"(���Sh�����"��Qe&��m=o��N_Đm��5�阍���t]v�C7�GĜ1�ՓL���Ƀ�)����nf�*������?�+�X�a�ټ��NF�@!F��T�:�܋�4���j�����t0Vܝ��v��I%tsFѥ�l(p^ߏl����d�%��p�t�G�B1*� �0�3�˹�Ft������-�>�Wh�G��9a��l5�Ty��n�?X� ��qG�3��f]�����ل�Mr6�Q�<� ߜ�4&�"G�G��P밻���h�>���Z�h+$w�A�������c���kqI6�^_!zw
��*Ձ�m���n�?�!CQVv�POA�G{���lfAC��_�!@��DVe�W.(g���G�.D]�HC�hP�|�JDy9F,���1{�`�m�	pET��e=���_��Ku�?���鐷��;�۹◷7ޔ���O9�I�g�$��ыo�f���8�<��O�B+�uZ�Cn�T�6^�A�5\&��6�ޕ*9l��`F���y��	6�m�C,~;$;�y_�>���.ή����+�C�R愳�V�V>�r��<��jm��{�Ãe�j��P��'�^}�+�+b�B���Q��.3�^4������%���6�ļ-�NK�����9L�πje����q��Zw��� �&�?T2�)jG[{��x�3 �cs\=�	����`�m��y7�I>X;C?·���U�����K�p��\�c�����A�-�5Z1�JU����J�B��&�cl�'
7!����L!�Bi�xj�s Q�L�-���K R�P�v�+�5��`�>���埊Zt�m� ������߼�?�}��܎�/�K=�B�_�Q��?�Y@���$Rp�Y��Bv�4���ɯ1gj2���gU�j�p�GC������p��/���̎�Y'K����; �*i�؛��~6[J�1��ъxȶ��Bz��g-������7�t#9~8�q�q����HRm�x���io�c��,�%~�̍��`HW�pRj�Ə�2�D�aT�^4V�Ơi�6�D韣�ȋ�b甍(U��S]5Ԝ�_J�?�T3>G�@�ÒS�4�!�i�-I�U�"��II�~Gv�pW2s�V����N%�ԅs:�0н�z��K=�,~)q��Vi�7\6��eH@Cw�n��m@)�ʊb L�T�㽐6�8tZW��J��[�#�G71�x�Y��~1�q�Hs� �IDSD"����[��rd��� ܵ�Υ-��Fv�'�3�v.�f�l)8�����B�ul�"	�K�e'�]�]�5Rs�Wh�Q9d�����^�I���h����ơ�,�h�����G�G~�kx���HN�IՐ^�R���!=Uj!�w�[��e�Qn(h4r�;Y~�E �2QS�o��˯���e����!��ퟌ�W���VېP�n�JM�ѱg#�,yc�Us�:x�Zgu�X&��I��/��C�7FvU�>���P�'�謃�@�5�챭��y��P6��ۚ�
�v����%�#�$��и_T_=0�L��s���L�@MW��q���bp��5��]���3�yW����r �O�]�@���*K������~d	�.�_o�=zk`�e<=�W������nE��t[k[C���K���3��#��R��#Y�w��,��s��w�ɆR����3qJ���ǚBN�����o����"��s�6�I��:��o	��'�%3}��}�I񗦅��1����<���܈��6ʂ����=�P�Ĝ�W�~N���]v��췬2v��k�	R6�����O$Ȏ�iU��h8�0R�G��h\�p9�|-C˗��bS����C�%؄�6�ރ�ʙz�����e#��R�P�04)D�hh���|�"��+{_�����{+ְ�M�4��dl^చO�����P�[柚A�iKX\���iU����Ϊ+����'"BX0f��������L3��r�F�����/���4��B�X�n6�s�:����3�p���(�He��2{q� O),�*u����ri��2��J�Gbi���A�وdP�X��Mz��e��4:J�rF�I*���������r$�Y������ތy#��N���1���!����zѫ0��-*�V����6@?HT�&TuOZM�u�7�#�Mdm&	��t�0�nR�榋D!'FA2ًpn�>�ⷷT��.�����Ȓ�=$D�m a3���ͨ�c�9����*e��ԏpY0�z������{]�3W��0a�=���gxt�b���\����OӲ3u�A�v4KM1ҲƯ�%wM�8_j���U �p�9��m�8?6�eb�@o�ZRm����lRy���"��CT6�Y��LiHE�sS�'y��i����B?]�Y�n+�h=�}�O)�Z�5��!ƌ{�%��'v�L�3x^VZ]2��T�=]���ښ6�����&�w�jkؙ)%�;MϘ�T\=q�]U�
�ѻ/�r�uw�W�#O�son��-JT}JP�R��Qa$���u+><���>��e�pU��n�y��?RR<��<��!p?�A��˦e1w�3����N�km_:E6��M��O =C#��^�fq!K*?��z�7.]�.�s�;G�_��!3#@U(�AxW+\����b����j� �)�`�h��O�gp��o>�!��,���O�m]/1��1[+;��Y�t�]I@s{�vI�ij<$�_���{�;Cٻ���9�/�����+�D�$G�3��:Ѳ�i	_���À�	����u����i�1)h6�ͣ����
ۆ��4TaY�<���M�얨]�JI~�mO|�V�? ��_�K���m�
_�Wgr��S�w_�&\�*�����L);�aE-��Fpϝ���4y���b;�OǗ���&꜔΍^P�@G�S��<ȣ��1�#}4Y�OOL�2�����C�_����K��\_�,�� 
:���A}� �m���;��J�*��n����D�9�Y��IL�輝d�rt�u^WN�Κ!�c|Dk�񘅠��'�f��C�T#�r�+�1�D�	���
�}��C*�4��X
T��~ojq&o7���U{�LBk��p����z��E�GH���+4�W�Y��yA��%#i��	2$�(	� PQ�w��'�Q�hB��D��#Z�R-�!�S5sƉ�xM$�}$a��5U��{�+1�Q�`r����ʪ�w1�
�?E�+�;;V�S��o ���������[�Y\e=e/�Ջ
	"��$��R����̧=��,��Ӂ��S��j����%23(5��,O�r�Z��$\��V��Zn��f�0|g�`?+�qu?���
\����oaQ���.z/���q�b��F?���Ã���K��tֹ���\����O�>���,틹[Ѣ���k�Ėf��L����)���r�d�����ь�d;�wb����P��Y�?��,ٜ�Bl��;f����'��"m�&k���ƙ&� ���F�8�;�bd(��-������%)���6���2��)�Ԧ��A��=�vUT��:��V���xA,RQ"�]�\���.�����)-�35�{C�t�f���;���y�nD��
���3��
��~�}ew�9�ڊ����+J��M�����t?ʎ ���;�D�F��D.a��C��p��^+*
����"���3f���e!y�̔�lm����k�o��IN"�C$z�a�tx�YP�#���6]*�1�Se�Rn�M����T=�
��]�>��S��h��	��Π����&�~d�r:Fn��q(Gv���2w����{:�;��ifz�n2�޿�K�GZЦ�� �-ݯ��8�O&�%1��p�&=|���|���e5��xn��#z��d>bw��Ʀ����lr��.S���F/���q�a|O�R��*�[�6�[^��i��"Ɲ[0�������;���)��+�5�6q�������>�A��ItK�:�*�68F�jl�d��8��w3J��]X�DI����]�;`��Z�$4�h�}ʋ0�Z7�#8���59�=���ؙ������7�R��X�+Vp+�M�K!H6F�<m�}�?e�ZY�5�]�6_�������>�0]$_��a�.��\Ot��gH>n������p#���<W�H�����*n���v�Nڼ��G%e�H�A����@���������R��;><6z�K�u�g�Gu�vG~6�+!>wҴ�&�3s�ŶCV����d�/��O�V��'������j����\�4���`j�`Ըe1y���-/�_�>_�6Lu��K�A��[+|[���"�2��XR���+�6�5w�
��ĭ�7)�`պT�f+W.:j��. ��.���UV.��b���/H��pr���v���e�`V#.ehg.���K��D{$��~�E����q Kxa��2NH��w��y-��"5H0VbgA���OAb�[�}6��/&�u�d�eo��v`�0�����Ũ*0U�(�ox�y�%����� ����9U&,!��-[��� -��Q�=Gv�79nO�7)x@�`�Я�4�`[�c�G�r��A3�A��X��r�]�BI�3;؊�)���y��
�Jg�X�̓�>��ơ<u�u-"2���9u
4�ѥ��k������*j�����"�c)���|l/��ױR� Q�O/���ANJ��Ag8��U�iG:/E����Y=�� hT^�:��~o&̊�c���� ���з�a�]�D��f�/��=ܚ��X8��(Fi�~���?��;�UlnA�W�s!���ֿ��..��7�U��'��U�ؔ�+T=���tiD�s� ���RC^*vlh�b���������b�#Ni�省S�4N��%0+�_�4��'O!z c>�eJ1l9.Ч� `�W�l���g3͖��+���!�����8�	���+�ar�*����ܭ�#�U���������d��� ���@�R����Fv�g_!~�s�p' A2ևK��������?�O�o��/���Y�q[���̯�0�X܅�@���ɡ�z�F+mN6��y93�q���|r@����8,0$�+Z.o��f��Ϩ,?w����(�F�TZZ���
��9qW)� �C"��C=L�ouĹ�x�E&܏����2�Q�K���*H�Nv#�;�g�qD���e��?t�����ř6�n���S�r���u��)��/M��d�i�x��P��C��cF���T�ffi�;�� �l��G��F�Z��VL��{g�ҩ�ǘS)r#�%�^��ޢ�Z؎w7��5\�Vۺ+�}D�I2��2�}�3O+֖�{>C)
�vrd;���0wtW,��E:���h�����cjv�Ȉ�E�WE唺h!ݻ�3�bUm���B6fc�>xB~��z�Cڽ 5�Ch�H
�|�G�͑�[@�HG7�њ;oу�XuИ
~�I�z�*Oq>�̄���tnH�Gt���pdtN�XNq��Ɛ;����t�=3F�����5k���p#������Ñ�_4^��� ��UC�9� l�q�7�<KҍL�VoėO3�'����bS7Y�W��j�5|�����\ʢ�Ev1�&��vI"5v-��*�K����R���Kҧ�  ��Ku�xy!m�G�i(�'��@�����������]����C�݊�g\��H��o@I��䓵hl;�CA��-NTV�!H{��;�['�o�*|��z9+d�\udO��=9���ʚǅO�W�J�9:�=�&�'�w�Ab�9�|��D�투�Z�N@���S~/�D�X�S\��-tL�d����D��q��)��*�}]�xm�~~��ܬ�^g����k0wS'Ь�֟����G��:�_9��e��N���w�()��s�8�yC��˩c���n�V/����ɑ�4��3��.��k���3jt|	���k�Wo3�a�b�G�BY��½���2~���?C�2�.?���	2H�Ț2�2׼�lqc^��=��T��mV�zH��^n}�Q4_����Z�&�cIE�X1�,W��+ͳ�<�.��X��t_��IO���>�6y�*�C�f]v�N���4�gg��c�9X7TC8�X�G<�:I;���-6�If&?�%hk�	Xt��.�E^�I�\��!��6N�Vn�Ui�V
*|���g���k�M�Lf��JT�" �d3��v���zB���^�N�j2j��cc��l)ȇ������O��i0��Om*
U�Zwv�A�C6�{����(���>v��k��۩��x���*�<��D�|����3n��Nލ	ǰ��4�R����&X�-t�0�9�ʨ�v�s
p�����*����n��zn}h�-��pxZ7�.��b��p؈��$3�'(<6�-O���f��AJ����0ƵM���/:6�I�dIX,_:��O�%]&ms�V��-���2�BC�_B�]�Z�GӤ�ԕ��T�~��������hc<*���1�ougB�H�}�no�K�hO.�t�V$�HLF��ztDRG����+�"��z�y��}��J7t�80�p�[��[:W|қ%di�4��ӝL�Jn�>(Y������uq�}�g�4�& �a�*��s��nJ;�L&�P` ����X}�J��3\cdtY!f�-��f������vR�h��5Y7���80d�X��>�Q�D!ΨT���`^��3��n�Z|��ؾ+♧���ͯ��kg4%�����ɝ��tul�J)!�_4�/nq���AM���2�{�?`�����ž� ��z'H.����	2���)�z�P�}���(���շ&�sJ\��q�Fn�=0gY����\��5	�k*�EL��J�Ή,��J|o"���
��Ml"�WkP&���G����8+n���<+�l����)�hS�ީ�[�,_yY#��a�Q6E�҄���ͯ��&�����T���o��%��E�-j`�dԻ��X�>����Kb�]+�����A��]��K�95i<�؂JX�V�%ih��Gt����x/�3!�ѤFiD��W�AG͘1���\Sb�����yӰp�ȅ�qA�<��l}����ן[)<48��5Պ���@��}���i������Z�N�����ȃ���s۞����҉����Y�07�&9�ԠX&Ҕ��J ф��(���"w�J���/m���2��m\��2�y��A_~fF�S�����3 ��8`uW�sC���T�?��6U$�5"�\#����l�;mf��q
	�'H�	<E�I'���kt��M�rd�h�y�f#�O%%-�usx���)�v5ӅvMZ��Ƀιu���o���e��B��ǟZ�D�S@6R+2��oe`���{����[vM�뒈X,�)·�k�57�#e�ѯK�S�W>�3�f�(+ޥl�:"�D��q�H����ړ�A�F�?}���0B��z_R�� Q\�e�?��j<��ܧ�ox�(F�F6��.�*�[�|�K�%gZ����5.���]I-$i_ ��*bɋ��Y���{���Z)���5�%(���dy�7#��:Ӑ�k�	z����k��.������{⯿��@�k�d�<��k �<
�s���%Q�_Yhz�	A� �@����^/��\Ґ���
�vP��P]!�����<oG �h|��)�p~n�{��G�� /��^���__�i���y�N5��,��$�3���p7b���%j�k�~�I��LF@��*��	��t7�M��n�I���l��������#=�eɨ�����~f�y�|;�s����O�R�j���X�J������bD�����@��|�sj����r��K�Q.�MW
, �D�b�I�:��4�
�M�9�"닄�q�z�T�U</�!���n[�	O�� /M�����S���3\�Y���h����t�� �:�7�դ2��ҿ�~��[{'�d-�@��Q�:'V�,Նݭ|�( ��E�I��ʥ��R��\&��S0�m�s��ȉ��/��zR�k{�mjL�m�E�-DȴA�0�r�z_��b^}�A1�2=N��"��r�fKȼ'��U���n-a�a|��a�@�e�"A��GO�̷��p��jA��_u������_�뒹d	�fJ���8L{^�w<�0'�E����E�C���:چ׭@�g����=d��ˊWF߮��2j���_b����D?�����˝-�"N(/fϳ���j�$������^�#����=�C^�{!�q>�X�t����uڰ%s��$��Q����j!<n՚��H�(��0��	x����s�6�Z{��Xܳ���r\���Q����f����ش�W�E��mJ;sJJV����|dX��Jd�݂�G?( �H�4�t%�����}���� aD�^mI
��O�i)f^G
gX��T�s��U�˼�TH�:��M�<Z�lK+�
䌿�!�:�i������G�(��w>!�{��S�TQK�6�_��<:p�:����r:_�T8{��R�d��,����\B0}����ɚ	�Ɨ�Fx'Y wմ�P[��"ʈZ��s�(*YT��uo�	�7~��4�I� a������G +f8Q#�g\|'��m�I��@C�%��K��`��K�?��bL8r�MI�34�ӭ�e���c�Ͽ�Ht!���mv�g3UU]ߠolU�F�V ��<�v��̮~��kZ�G;ꇲ,!�]��O
ޑЄuڭ��~E����Qob4U�u��;\�(������[c!d�xļ��O�So��;ЍnX>H���bh����])�r���y�,ˈ;��7��%�~)�6%�I6Q�a{1��Ys�
s����;ܸI��M�\4BYHm�D�d��cv-�T������P��0���/��[��`�X�k��bQ'���o U8�PI1�D�⛉�6����7��s���ĝI�
�u����~�P\���|uˬ�ҳT�TGq�4b.筍�G��y=�60�#�Qm1�n���p�8���[��B���{E��$:``��-�^�����&n��g�ɖ{0����<�ޟ���P��0̥�����.1Xaf�{'�Ȥ�boO���x6y����w�H=,<@}��:����0bo0�c,�wI'��۹�/��(#*bm�Z�a�J!�'a	4i�;�A8�c���y��q&��u����P�O����:���+��
Y����{�Oq��)�S*��M�o�8ߡ�wXنB�ҷ�XӬKh��IxU���@*�ɽQeb���c�e�;��������%�?������2�g����ܶҰS�Y�m�i�U5O
���:�A�E� ��Ab�BVIv���C}�������"6�}��g�a|7y'��O��W��]>�,����wG�YL�d�����/�ܚ�`	��8��������9R`��e��e]���Ɏ�Te;��w7��?t����S�����j�-����������f�\�-P���%I� .�Z�f�|t�Y�Y��k��P���E^���ó��˶i3+7i�C*U_λjQ�;���fN�AѶ�� 	.T��� <7"
"a#\���6�+���_ܴx|�+�#b��a�L�Z�;����.=WlJ�y�VEp�Q�Ĩ�7�
�-M]y�4�u*\�"�k����1�2���_�o�Lm(�252�Ԉ|��SqqC������/�{k%����O�P��Y����ys1���W0�T\��m�{�2Kg_j��b
k:�@�<���>��1{¡м��61�y��B��YQ�TX��|p�J�)�����i@RB��jF��B߆�`Bp��x���WF���F�ڄ�7[�F���Q>����\��q�/�l��%��}���������R�E�;$I	h��\t����ՒC/toI�]A�R7�B.��|�} ���.W�!��������ͩ"�bs=�Ӈ�>`�՟��S���WshP����vZÕ1�L�B��[����T���W^C.�A���/=_����l-3�����2a�tC}�/�/��NoB̙tf���ٳe�7��62�C�6Q\t�\S�5����O  r�n` �șK���K��K��u��v2�qT���/㍍G�u��-��P����Y�_HL��~[:z!�������,�HmS�,4�MU>�n��M��ʾ�.�^~ʰ��#�Ѫ5�D~���_�5�=��:S�+m8'u��ў�޹h�QPk)��޻ �v����Ӎo�6�"� DĬ����m`�q����Ā��X��:�&._r{��]��1��Д�'�4��R�Q�N�Aߘ��D�5���((�0�<�D���[d�#D%��e���<Lm	�w��B��t��5���8i$�[��>���vc��8ɏ���%��2W�>�|@�,����`�i0!��������|��F�Q������+2�����;�֋:C�G_���p/}����cz�[r�ޯ��S��יhE�)]B[܊�܀�?C�rb8�ͬkPKbn��)1�r�qa2�g�H��p����L�y߯�7&KSl>�Tv������	O�7;�g�oK"7{��S���؍.X��7�l0�;��ԤL��p�v�=�d�H_�&�>~;�i򄾮cΔ-#��n���ֈ�o���d��U]�s0��+*ɧ�Ŷ�Wp���L��*�e���æ&{I?�
هYǟ�"��4V̓�n���3.��h�S�&�&f�fC�edc�?�w�#�>B�ڭ��O�V�w:[m�[�B�*k�Y&$^o���!q��j�ȯ/8p����1��G�� ��)Z9��SK�=�X6�Tz�LKsd�]�D��Y�����K�`o=��lG[�-��-�)�]��5��=g�-�h�Q1�|�O�6��s�~�q�����B�6u��"�ȧ�m�6�+i�4���Z��=d_�6��}�Ȇ�/d�<�<�k&صw|@�F�
,��Ƶ9k���X<�"���+D�w�Ly!y@��d4����3��eȐ��At�C�R�L��}����=�=�_�cuG�y'h�L���UyQ?g 0(ՄQV���~\[J�ݽy��o밧�|,�SL����X�H�ޣR��a��+>������>ɏs:Ej�C.��8�����?���!-���n�;��0�K	y��h�Ϥ�0&\��&�(��	�b��o�i����mE�)�b@i����[I�|��-}�CO�/D����RM�l�[n�U��N�R���)�<�[ 6y�����F��k~��Z�m�����=hO�/�*Y۟0�6u�WZ	W!
HópB[��T/�N�αM����ŧ�Bd��,���Cx��:���o�9�/6.�%���:ʼ�s]D���F���jO2��- �o� D����K����Ԭͽ�f��42�x1�<枔K�
Z&M��vڔ(g#G�Mx�쀹�ǆ����%õ�T�s�I�X�v�u�eX�����TGFc!u�� ��ԓ%f��*�_|ª�d����'��ő^R�}���y�9���+�>A���i���h4TFg��Wh���X֟!ƭƟ�oXQWh۪�m�Q��������g��Z�׭� �Pڽj�%��PDn��;�La��j[E>x Y�s�VZ�&R!��[���M�02� �~�X�D��AR8{�s�$A�*dׁ�:|Y�^�v�0H�[��F��)���F��BqgT�����*�Dڴ�w����؅��K*�'�dld��s�-��-�
�r7z�����ʳ�q��	)m��&٘l6+���S���+�v�%�(�`<I-�#W��у���Q���M���Ɓ�p�Z���b�N��$������m�E6�<5��l\��Ǌ�г�P��j�(�<���[Q��5�P��ɦMhҼO��s�)ׁq@�!Ml��l�#��z���Б̽��d�&_}
r���W���#}TLDɓQ'��1���]"n!�����n;�le �m����&�S�|�u�o�9�I�p�!M��x��)>��%Ν���7���R;�����tb�E# hpq�����#��Bn��+)~�#i�F�l*~��n�P)O���"��{	U�;Fȼ8.�R	"�j��`Mł��%��6�抢����E�&)��5��A.'	�Q�C��+3����Tf�B�yi9�I%�7�B�b�[fJf�Fނ��aUƌ^o;�~�[��KӁW��b���x�q�Dg�<XY�oK�	�W]ZY�������xM 7A�9���R�h��L�$���Ʃ�&,�E#��Ȼ�g�c��Q9sxc0U=EMb`Ė���/�ħ�C$@��J�����W�8�j���O�]�痖~`�������7*�	p�Ä��J�M�Q�����:�[4�.0������G�ov�-ʣ3#�Cǁ���l���8)���b7�2� OJ���X�F��[h3Y���&�Ss�NP��=����4bA7����2p�&*�TY���1S	A\��Y��	��zHtMd��{~���@�C)���]?ǣg�"��Ju���kM���Ov���E���ߣ[q`�Ë��g.�蒇�%�:u'vl\| 2.�Y����=�ҩS�>>$Q������z�M��X0��a�� ��s�^#�tc�C�ō�C��w�1x��P#�� ���Da�,��Wc�@���G@G�t�NV���!1�H���E�9t}I�liUgH/D	�@�����Z%�*��^`���i�(��(�����6���}1K��Оq���lN\ZZަ$�uNSI���N<��䷰2�����D�Ζۉ�zR�`}��[�	�?��Tm+*t�I�H�^E�ݝQ�x�炋��穳j��%�Eq�ٓ�w����G@�)�)�5p����CO����J���dA�:e��O>UE�����(3R�LC'�?H�|�7
`a�!�����͵Cy_�F�Ė)tY!���i
�>0� d)�9�0� �x�����T$��p����^~� ؑR���ٷ̳���KwA/"�0����kO�St���>�C_ec�Ʀ��o�J�3jڭ�@�Ro�Y2�j���so��� �S.�a�~�!�[4���*��6����P�M�##n2%��JY LF"ғaZU}?}w��p��'���DyT![][�5���.l�7�<��k�^d�7y̻|�{��A�I!�tQ�)0�g�)3�ev�YGi3����`IЂ�<{�������R�$����g�0�)�@3����
{q6�+R��d�4�7��F�`Y���-�|��W���>ؽ�y�I��@l����O�󒛈۾e�����	������;�B���n\	�JF���yA��0b��f�ж�o���Ato5��Cн�|�(t�
��6��<p�E�3(4�C4p�� d��yu�9\B�J��� *�: �.�>w��鸜3���>Z7���%���բϹ�f��j
��V�w�!�f��]�(��0�V��$�% &�wQ��+��q�h�?��q]��g�І�O���p3^�,x�c����Ƹ��)��<���7��\D�&�^"��v������@p��I5c�Yؒ�Ud��6a\t~��VR�N��tG̈́�V�(!.x�M��y|	`��Rf2�xQ/$i��$5͓;g���r0З��{p�n����bx�I=;��=��g�t���Eމ��$rx�rc=��P�*�At��1�Px�]C�e��^���SЪ�v˸v�1�Qe��
��dʪxTjO���5��Ob9��B�++弹�A���aX��C��Wuj�h8��� ���/k��lb}L�m�L���'������"F_�w�TZ���
��Z���hɟ�r>_�$��?ܼ���b�W�,�mT�Z3�}Z� H2k�}�Uuz=Vo7��H���hOx�x�e��Q�cIN?'�BK�ޠe�2>cNt়�s�%��`(x<�hz��C �g�j��EA#���n[2�x��P��?�D}��#����p�~�[��M����h�;,�-a�}$z���K��Hb-GTЃV4�:Un��^UW�H�AJ�Z[4Qk"�ʃ��6���Bd�O��c��-v͛t��NO��w������Q5�Q���[8���i�D��$Qc�o/��x:u&�=�Y$_5�Z'����N;�8���U��D�v]ހe�q}��ҢL�02�Z��ڤ�L"G��Z�By����}-d��=6�H���ع0���msn�C,͝P�B�|	%p��~���bex����c��猒�e䔫���L#{D�Mx��n�=�D��~��]Ӣc�5����E���{�~g���,�b���q��u��fts	�j 3髼������Nļ�j?p�vсX:��@cCCqy�Ϣd�d�5��c��޻����p_�#���l���v��(�
��q��q�\�MV@�(�~a�ބ^/uZ���]t�AyjD�;!"�y�bw�Gcc7����߹�	DD�y��p����~p
k��_�e7݌��{��Il;�"5���O� &�}�[� bG�ب�v�!���h��T���O�2W��j��8���D��
�,�S�5I�M/�S�G�8�6�~��n�2^�]���wE���ϒa�`�4�tl�w )#�1�S;Ko�.�u�-�.#��m�������X�,�5�:k���~qyW?�⓸�ðs�FdVP\��f:�*>[��H��"2X����� A�>��"9&L��C�*ܖ���h����>�l_>	y9��`
�����:Ń]������L����,�>��h�fi�i�V��o�&���mq"�l���,���SCU^��m�s�tcK���tId��!]�7.��9@���}}Co^��*�l�a`Ag'Px��E�l���ް(-~�t}�A��ۙ��,I0?�Άބɬ�B���6�Te#2�W�,��I���q1����jNڣ��M�2��npʂ3yx�6�I���ڙ�<�c�^A;�(�YD��c�׸8d���8}�0�����{>�X�q��/e��_*�R��� Q]��|nz	��6����F.RN��z�x]���G����t\(V����O0יə�d@12̛����蔾(��g1�<g��Q�Q�n���m����3V��(�sQ�𲢺��N�|��q�b�B�NT4~�>|Z��-�Z��K1��YԵ���$��c�j��:B��,E�#�;�C3�E<u��|ͱ�r������ѝ����p�`���J���$ �E�ijN��X�eIL�ӅTޤ`�����i�dF*SWLKM��6�_�y���;%�
Ũ���߃C����X�i1���~�7������l��b\d`.��B��ЂѰLCy�綂�JixIqdR�)^���3����/�D]��Q�U��������s�����)�Q�C��^�>Xt�'T��������L�.���e#��m5��x͟K,v&HCP$�Z��S�P7ZBV���c]qܣ�@���K�sϮۣ�bL�N�����1J5׹�
�x�2�P�j�X�:�%B� �h�S)�(��:���5��u�����k�Z�.�6��e�.��{CD�}с�y�Rl�K|f���g'4+��\��r��*D�O4ѭ���~j��6�_@��Xߺ�����΢�[�"��"�c��0�l�Ie�=i����#��8#�b�N��(q�K9Ob1�m��R�� �P��К�>�v��Wl����q���׀�jj�
D�<溢���"W��iE�g��5�t���NJ
�4C2�9-�%U�� �f����u�b]X�2�PesY$�\��U9�Ul+�OD/*(n�N�����+#5 �+�7<��4�v��:%�Z�W��D����������e�ʤ��,�8c�\}I/f�xW���;<�+t�P��X����3n�BպSߋ�jM��_ғD*؃y�����΂ 31��p�q��8�{�6l:��Y�'�(�BC��9q��J�b/��T*֩8E���z*�3)��-�H�#W�i��!�q�b�?c0�%�xm]X�ZW�pC~/q�n���<�空��+�f u��y��1t�(���E7���6`�t���e7�����t}�PlHWHm���W`�J��,��T�r��U m m�A�����ÓT��f�1f�h[>�k�f}��52����a�%Ba�}q�ԩоޘ1d��G�躵�7�hN�)J�VY�Ø���J����FQ���WuK�,-
�T��l?��=�R��n���.RHo8�{�Yd�Fv����6�b0��l�=+3/�`I�˙P��A��z7e���NP���5XV�MN�j�b�����kWf"Kn��l�複!ߢ��F/�ϒ�Yr'�qf���5%���)+��Y��3��o��@�soٿ����_)�x34�!@E�M��f����q|�eW�w��Jŧ���Hu�����"-���W�J>�r|��ab3dq�T*������ۄ{c���0MR%���]K��(:���Km4|6҉���벾x�? ���o��u�<�D�nͱQ�%�\:\�Ԙ~�m�M(A��-�2�An���r�I���+C��}b�,#m	�qCLx��tCԔl�޳\�n�d��F��y`G�>4�%�����"��k 3��Om�r�L�*�����E��S�;l�o���='�w@X��с�;�K�7*4�`�$ڱ�����Mߗ�ì1�Jf�M�F�����(t�^h��].Np��ٲ�_�9������%X�
$_�pq	��)o]ؔ"�	����!����n����X���~F�cGK(d��b��O3'f3���+w��B�Zd{HYE���*�fӅ�'E�wO'Y���e�r}��V>�yH#n� ͚BO��� ��ľ}���/.m��,���p�-���2��r�X�)g!؋�f.;�P�T�F����ҫ7eI�<����*-�XHX(�͢o�ބ��2�#:Gw�p��i�l��N�T��l'~R?�(��b^��Ͱ����([�*ن`��˫�ߎ��;�L�6e��+`|��;�gA�����&��7w�7۫��)�X�п=+���l��7)��>'��ɋN�Z��7�6^�3m`t��1���,b�� �F��!�] ���h��ǌ�vF���z=O����Z-�.�b���19��M@���7]�RV8Q�JL��/iҗ�A���U����L!{�e�f`I��I����Tz3"�`,�r߶[נׄ
{�D��I�W�]KX���X�N�-�O0uxn�R��^��"#��д/��=�\��k�k�.�F��Nb@�O�^a��m�S��S(�d���.�_�B�tpt	�0g�Iۊ��NlL���I��� )����&/���0�n��eV��
������^ �x�� kQ�=�C����A+�������x�o'�,"��/�g��*V�O@�	a�>l�.g��:�bCa^)�л�N��ܸ��%��nÖO�T�����+�	%����:	)��nO�-W0�j�[��Rpw� �&�$��R��pARZ(��$#:寨^��.�At��w�00�Q(m��զ���Fчb�*Ma���Z�/�:];�J���{�����[�N:б������C��s?��u�U��C9�X�R�ޒgl8̎��ro�u)��Vo��W�jz�n���l�o�4C�_����(��H��]�GoE]-���:Ԗ/C����]�g�����N#��E�4�4��ǲ�ϙ�zm��e�� b�0�^m0�ƃH���������+P����Xr�uvd�����M�p���ɇ[H��-���T��ʁ��Pl�� �%Q��������#~����� �I��T��SQ��#A�f����t̩�!K�Tv
�:��:l��T}:���	w�)��-��/4y����"p�%%�WB�NG,�B�M�m������x��ͪ�?��ឣ�N�s/,XO2�9���%��G̮�b�s�7����^�;��N?է�i
ы 2��7�宪��̿�O��RZ��g���q��)��S^*m�� ^6/��;�Z�B�!���Q"#IŨ����	���
�s|���k����XtC]����t���œ�� @�*��.���U��w��V�2�#7;,DZ��
�'ɍ6���x�
�<q��:'
���嫱Gmq����G�b��Xi���{B���%��m�-��R�n���Il���A
V�EWC�.i�=��c��x06�OC�(����u��/2[6�m��7
� ����@�k_�����-�B�f�����+)�d�<�1cB8c���B#����g)͇���C[*X�6�������o�y��z�D���9M=z��D�9������q������U��U|��3�۸��_�|���wtv5�A]c,i׊e�8��#�f��*������(��Ӕ榸�\`Oz4��J�r��7�i�>��D�f6�$�l�����"�(�tXϸ�0��Y_|Q`��
wE��q�;;��D�^�0?r���ٮوiW��vJ�ČX�{��3��
�BZ��.0�a�R��K9sƑz�ѿ=� ��;6��>ǔS#�������Q!C�.G�Shw>��ȗChn�+��$X�J�W	���C=)�������H �ۄ��f���E{��*N'M�i��/~�Y��Y?]I9ͳr�D0
�u��w����2Ѱ�A]c��P`Q��x��잜����P���`Q��jX��+o�׼J|O
���f8��w�o���>I��B-�A�C�^Jc���J�S��i����%����d�}�ɱ��$�bTFB�trK��:㶅�c�*�gI
ت@��$��ɋ�|�շ'�EE�X*r��[���R��Ol�%�j�Mz_ٝc?���ue�e��u�;�X3��rt�]���o77.���v�u$�y`Ƥ�wۛ\�E������ō"<-Ľ5��ZYj��պ"�s����h�|�W��/�%��+��B�QĄ��玚�z�+�N(���lI�c>jz����B5��H����};ubk���$=���-�Cr���)i��_G��P����ޭ8+��2=c}�_��=���/H��8u{k ��E��c� (�(_���~�;��I~6go3�(����K����F��IU$V��wRbT��̖�Z>��go�G�b�yR�Pu�l����Z�mA�e���.��`#U�'���jT��[�4^�EX,L�y�G��v6(�@qgF�� ʳzTM�A�:�!�T2�@+�%��[%Y���DS3�;����}��,�Dh�Ԟ��%�������׍��'�u�CC1(�<%!�u���*6V%B��#��$�ɕɸTN6��Z~kii�ꦁ�j�gL�l������[Ɍ�/-o@��$p
�=�嗫�����K�!��:mY�{v�E��{PW�'�p9Jr�5�20u�k�\��=�����9�x0�M�#헩ݡ&���D:X8J�����F˱.������<s���b]�`aO(v��	c�F�`���l��G2�0�j�A�kƆ�'�M�1{S)˽��Ǔ��ǖ{�K? )">�هMR=!ULph�K��7,�t�xi�9C�L��W!�BD���Ym�#��9������>HV�G��s-b.�6�b�Ɗ(��UFH���4^(	ea�K��s��T�)�A7x��-�
h�<���Z���E�]��̟�P��-�z 
*� ��Ԣ�n�'�D��YO��.i�9);���H֒����A�Ok�M0��ш��Xϫ��L!�C�+O�@��yQ�UNMh��Jw��P+���g�a�x�W�*=��Y�
����6�Z7r�ٚ�e	_*��Vr����>B�6�Q�|,fl��'�_����\�r8�����8�Љ���Xo�SA��.����B�y~
��g�Z���p^�5p���,�$�z�>�HDs.�Ϲȫw��� ֚��)\E�\H[C�P�-��!���(hLR����9����X�0�Um��;�#�	�<�p��|�/���z�����C[�P�[P�o+V'��=|��	)�mݼ�	p������ʝ�2;G3%�ľAW���%N��K�ת�m���\�WeF�+E����
N�>�9�آܐ��p�qj�8���L���ޗ�V.�{�)B�z� ���L�Y�-\<��Q�ܸ��s@�{�V.�T��`�aQ�J�t^Sd�J	o��4���k��Sq���	�/Թ���Ȓ�s0��H�_��u#i�ȭN_�S[��|�q��{�B;V0]�K)��5�(��V`��D�m��Ď�f�L+Ǵ�]�.c��i�o�#��Ô�w���Fp@�E�kق·�&�p��T�k�ʼ��l�L�=`O�ȴ���"�36�i��r1� tO4e/S!lt�g�"�Bv87�cSt��6�#�eAj)���t>-v�%���[v�˥�p8xN`Ù�.�M�0�~+������	��a)����W6�D\�M@���L&e�E[��:���� -�l��|[�,�d����Z%�7޳�.�S�(�� �����U�u��4V�F�����'��	�Aw��S�Z򘮊z��N��a����v-�(��9w����\�9R5;�%?	��*c���L��z������?�fG�m����z-�9u@kf������e��*wH#7b\C�sCY�4�u�8I*��h1�Po����+�eezO��v۷�*��̃Ld�:���Tm'f�v��AX�,=Q��Tr�a����D��+��H�q�d�m����CC�����̖x5d9�U>��)f�,7<�_uR�-��H(b�����%|S�W	���Q�����5u$��m�;D��iuΡ��p��9�"�V0\�(���W�ۃ�^D����p,���|'�Q�@�"top&%����8���\3 ٚk3��&�����*�o�w4V�6�(�ُ��Gm0C/�;��E�Dѷ���6���G�E�9Y��:D]�oAڗJ��5T$6}8Uq��;���%�Ȧ�П]�7�c,Zi?"�8�C���J���߉ڧ�Q�S?h�8��0C.ĉ n����-
���r<�i��o0О�3}6��Z�z�e'+�������7�A�,�DH�3�Z�i�����-yz����ޗ]R�֋��i��پ.��*�OwI�(!�jωt��$�K�.�]�B�:d����Օ���ҧ��/�S"9#��Ii&�ƽv,�y�N������I�,�|�:R�����n6�XsX�A��D`�9r�z1�O��z�@>�+^f� �x�I��	}b�;��dD �=;��ĭ֚y��˗ӡ�ɿM�W���P�ī�	���ic1��m0YRe,o鸱=�,��Z�����H��1�;�f� 7A��(W���ˁ3�����I�1�
<�w�A�ɦ��`�?1:b�i�>7U�7h�n"��vG��o#Ù����>ak"��er�XO��:vJO-�s�W���'5a��\IB���(�ct�1}�a��Yp���;�A��q���:�7��Þ#5�������	��5���/S䷻�T;g��OV�'�d�bcZռ4��<���񅢆!38�Q?�6��l�N�[�j.M�,;~�I���E�����הN���	_H�11�Y��dv�H��G\���i�wzʲ,Eh��Y$��A))��=p]��6L�Y�a�?���T����Yܬ�>{h�3��e�o�3��(��@Օ�����?����\Y�]�Bش���f�A��_ۏ���;$>�}����M�}�C�1��;�J*���.3��� �ht��@��	���'欒��܋}r!��i�7lX4�g�ݼ�4��\�D3�g�N�M�"�;"-��/���Έ_�w?z�����4K�Q���yK���h�Kb7�#�~���x�8g���*��B�ҳ�/�J�Ah�vN��EZXf�����4�j�]y2_��s�1׀��W"i;vVBW_9�S�Z&|�t}�ݡ����T���9&��^�sՅm��}D4��
B�gS�����Q���XG��qʧ�A?�A�O�O�7��Xe���#2_�Q1[�/���Q��{�sù.�}�4gJ�U��l�a�?'Ͷ'�:^	"t`����ս �zO�&�}�,O��zXRBt���z�o�%���A�l�6���*��������~�^9��@i�-Xg������c�G��kw��Mά�#�޺���D�:�<|�(�$�@Ђs$�yKy`ȖǕ���U������&�|Ś�
JE�P�y��#��3�S�/'����Tpo٬.����uV}���d�]���͂�b�:D�tNb1��
�1�	:V�y����D/�]�G�I�X+��+��c�e�X�e��_e�p�����x��#=ُ3������-��&��se!��;��6�ʹ|9)�o0*U����+o���9�=�ߡa#d�w��Xb�sB�r�)���d�t���ax�-O�17��ԭ덵��RP	)�y^��u����Ԉq�֦r����r�ule��=w$u�m.�,�Y̗�&v���t��LK�FCy�`I�V�dXɺ���B�~IV�q���x��������h��^r
<�P��4�?������Sճ����;��ɲL}Q�H��h��j��ޜa/�Z�,U>��ww�vח�S��ad>A�Kw�w����8��Z5������ L:�q�0K2���/DP6���/�hlGv�tw�����otu���*Yw�a�\���=A-�&�ݛ��s�C)���ظ��0z�pn�F�T5�41J҈S�a��f�j�oC�q4��ѕ��9��L@����f��'�85w��[���^[�� �ZcӅ����<@�,�ۯ�ǃ���8d��t��G���)�s~�C\���|	�v�ò��n������_��w���f^��-ܰu�����+�S�:��=/O6�����H//7R/����8~��I�2Ym�(Ͻ�y�t�����o�џk�V��JmE�֨����H�wz?�Vy2BcGX�vA[��T	��C4�aM�e�McN��2Rxw�`�1nq~���-/�oۏ�M�����3U`��ՠ���ظ�D�ȭ�����I#A��h���4	���]xYk$QiI��Ħ�Eb�4�Z�cw���_)�ݔ�=&�B�+����e���'�ǳ�����^Yp�	�{:�u���%��+�Sw�e�~���3�""��S��M�\Ȣ~Y	sװ��e1����C���r��/�{A8Xvf�:>�#���cQ�d�rՠה�9�Z�ʁk��%l06�AЫ"cY���qa0 A[�/!ܬ���{�Ӗ�=��>�e���K�7rg�p MȐr�.y��BB� !��5so���B���-��řA�;��o��M�]��VI�Al��Br|�5H��1E'�֗�������Vq�D8��_�����*]q�y�������s�ӑh�S߾�d��O��b����Ս����S�V,�M9�ڴ�i�;��kf;*����w'Z��,��`�O.�c�T�9Q2�F�{��lFiK�=Czq��+�Tk�n������y8ŗ��qjoCB`��s<\ �s��������QM/���2���M�47��s���'C��d�������Q|�>��L�iH��ݜy?.������%#n�E:'�� 9�}�����{�Q�Ҕ�v&�$��1Yk����`P~�fX	�\�7�L/ؓ�WmX���l��B����؞�G�O��A@�<�Ś�х�)PP�=�����bM!�כ2�3J
z��'_��o�S����&[4�?�Pb����`m�e[�M��ߔGΘ <Tn|o�|��4uw�	|��u��HѺ[�9�ύ;;Sf	o�=�+�$m���T|I�4Gw����{9;�G~��_h��o����*�n�쬞���U�I�n]�i|4��J՗�^��~������	�-'�F�x[�3�3s� j	��+��P>=�B����;=�!:�O�%WDq�P�2ʓ��F�OS����ը����\�Ϟ���ᷮ��w����&R��Y��ѻ>	YC������ў��	=Z��x�⒧��~b��12��uMm b����	��sp�jR!e���'}�0ϻg���P��Y��z(?�9���ZW#�N�m#՜��=%�+6�%�@,���\��ryЮ�zG�o��V_�TC�'�Fg�ؿ���]8�	?�R�R�M�/e\x)�|u��72��� !��\+�a�z&JD�l���0��麑�1__�f��e��U'񬫵e�4+Tΰieמۗ�U|��\+)��T�\�.�j��{G�� ��^�Aj}Wӊ��6��w"�/�Ǯ����T^kL�z�>?���m%���I�{��x�0�{�5��{�O$�r�uyJU*
��k_7�oj��M�1��=`�Ĥ�b4ɤ�"�a�/R�=��N�����V!a3����q166���-~W��`�e�9R�����aY'c�; �ᵊOio���:�9���S��5oh�=4��x)�����L���tr�A�N�#�"n����+�ў�rp��m`6�W�w*����%�(4���.(=E*M�p��,�QF�I[���QJ/�O�"�Uhn��?ۤ^���+����^��.�s8Ԯ,*[�`4��ǿ�.����u�^F��R�0}���.�P���$ˣ�I�OB����+�:��p�� ����d5����Lz�y�!��I�	T�0j��X��4r�`�E�����uA�H�	�� �aۉjm�Y8#ڣbN��I,����'���-��^���⠗�Th)�О�jX���XO�n~�V��mڽ�D�$�4�1Ӯ�:aȝP3�?�m?�қZ�4�;����ۍ(~C�[y�q��Èob�j�UA>�ZJ^D��]�ee�>&��>7�nB'�(J�B&?N��3�Su��ϲR�r���qG��.������>��G
>L���ˁ���Zk��2K����� �BP"����PUM`���3��g�w&�VD��Ej����&c�<B3^�|�s<�絶+0��+Az�W�n $霎��n�|���m�X�z���vPB5�����d^��K�X$��B�^��D/X���e���N�4�8yԖ�I�^E�~\�p��̹]���87z�#��10w����#�F��z�-�팁�Z���o� 2�� _�����;z���LЗIc�� P�Fּd�nW&̈́P�� �ch�e�ڌM�k/zQ�(;��C���In�RR֧{+����+�ES��ms?X�>���Z=���3`���4���Y�����a��;3�[s�_m 4�M��p?��b���թ[:��e8\}d���d��ΆN8�H�@b�;�B�u�w��̔k����_Og��1�k����kO�[t���w+GS�@���RD��y,by&��{��k�Ho�/�uP�A|_�6�������������8�7���b�Iv���E���������-g5�o�!�Je�*"��/L���ȲC��[���:��8�J�c~zI�/��k�Po5cl�tq�K�K�i.7���Ɔ�슬Y��To�j;�cݭZi���*��鶝t��,amt�?���Q�(Z�����9�g�o�{_Y���6{x��Q�b��G��8_�����z�%b	U��f���_�3{��H���Q:�]W.�A�%a]��}"��ܓ���03���<�(!�/��I�~��H��:�h�B���0~Ƭ[O�p����7���# ��j.����]pE��3��$�*����F��R�5�E�@R�F�[���J���!�����bІе��E,�ay�v���~V�B�6c�m�"Áp���eW����8��eT߆�OR��d���0�[�Bd:C���/�W_�`q��17@����Ց$��ޢ�E���t�����mҌ_ �=u�Wx	�w��o��j��x z���r�� �8\\�HO��3:�|�x�}d�Q�'ȧ�A���3�n�N�����puPq`��c�w�cG(�)��L�
Fl-�
O/%`��s�`���k�M���gu�A6J>��7 � �p1�[�2n	�0_ �6OpwIa�dc��C�N��}�"_\I�~��{v ��R�T��8�	DhWcSoQE��g�J�e#���l� NH�⁙5�=ק-����M�/�Ւ��/�!���~��Ӝ"^G"��Cߞ�F*��D�;X�h	�3��s�0�4��`�O�w+c�Y_V���f��Z�$��~ =���y�����|Y���W��Lk<�� '��n��ߧ��I��°4�����2N�d�'�f�v�S:F��°�C�V��?��ZgY�I�1�*�EJ`���~9�Ǘjg���m��zu���b��5ĳ��]i6?.����3/�r��GY���4�CT����7D_Ӻ����&�	��A�?��UL���Zt�zU�J���!eM���5f� ��j}���^�Ze��[�ܣ�D>�|�SᘮiJ�N��P-R�r�����uP9/��(����P�*'>����)r7Ӟpb|g�>��}�}�TIҕc@q��j�[� �羍�:��:!�x� �=P(W+�|���-y]��^V�d�1���鳿H���\��)��nK��M���[5��^���L�AolH�'�Ǘ�
G�������;g�;���=�E�t����&"x��{���i��cI��2�Ț�;U����!�
 �.� H���4a3�)Tq��]��b��I�9f���|I��F	O�݄�Z��/>��UM�� �Q�l�������g�cO�˶e� D���	�,qB�@��Y���4<]�A�� s�@�s"mNV�o�s�k8��� Ỳrd�BLށ���/w0(OXцإp\x¯�*�$qr�!/>!#�J��NFZ�&SC��L��XSC��;q%���������m���Fy��7�r�+����h[nF(���&��1��~�b��Mn���6#�śR�{g���;���C��ŵ�z���ҿ8�(#���pI��
0�İ·{$S\�g��+�?�TƷf1��i���50>4b��L�xy�v�fW��7Rzw��k��o6�5N�-���8�s�t�ƭ?��m77��='r:@�3`��{zȂ�GWG��.���Y�lg7}hu��5�C���z	n0-��s	qA��i�o�7�C�����=uVe�}���A�9�"k:갴>{��oH�v�|�Eצa��!�܊�-�j܈��KGO�#+L{��0v�kI{!,�I�5t61�p����v޷B�����oғףs�ά�
<�u�����[T��J�����D������ER�#��m�
��5g֥]8��0���w���Ġx����=�V���'����_c֤�+ N70�{���qhl�DK�(Q_�ë�Z�|Z���[*�#R3^�b*��+��6�IN��S~F.���ա"FkvL�QJe �Dz�w��˚�p9�i��3�̇ϊ���t>�<���=WPKv@��������*��Ed��Lx�dF
QW��Z�3�w4��WE'7jg�����V{ne��3D��"��"�-SrM��e�6�NT�t����k���0{��b|�&_q���L^!
'��P�p�+y"˟���{�>Z�1��R/��u��Q5��t�������@}����
�������ְ��W���7c�xE�|�2�}R4�Ɯ�����_)��ԥ@�d����83Pd1��� 5���?�4�e�v=j�ϺRqL}�D|"�fUo7�o8\%����'`a�ȥ���T$�i/J
$��&60�����s�1�RD0��<`L��)��*����K=��L���������{�څD��㖃���j������7�\�e���O���=ݱ���j�Q�MMY�6р�h��-����S�H�{	�7���t�:�؏�eG�X[ףo-�E�K���� ~�p(��ےU�ϟ7E�E�$ej�,h��3c?�A�NP캷J(?�U)�ݤ�a~fz�SH)Oץ����{	Q�K�~�V��+��R�Fi��lĞ���u}ʽ���IL�O^�!���ϛ��ױ�%�c��*�����<I�9Є��iL�4[�ZUNN�+8?$O����LK/��A�{���������Q��*�ųO�*��YRx���4���͏���w������:^g'�7tu��rV��yF���-��u?&`�U�& �Y��t���ߑAS0�c��s0��#Un�sۿ�/��7���I�O@�?����O�8�#ۑ.rYt�a�M$���S�1�C	�g_[�ߎ؅4hn/HE}�>�q3M'���uϔgI�n+D�`�U�ah�I{��R9��;��s��z��
���1�d��$?s5Z��=s��b��l�wC�jI� �+V9�c�.�s4@����+���}��y�w�a�,>��]C,�^�o�d�k���X]{>BNwQ�[ʹ��Vl�1�!��7Y�mQ�g��G�����F�Y�u�a01���}���)X0��&��x�d�]	=�\��F��owO�d�0Ә �l�Bʨ�Ou][�g�y[Xs9	���7�G�a���a'��M���,T?���4����a�/�@mQ9��g� ~���Ӿޭ��(��)b����πm,/�٬����^=�c�����J5�+��i5°��е{O���|�d�
o���'	���pDb�M��F�p�+�B�T���JO������eG���g>����ذF+3��sp΋X����	_����b�Z�z����K�b�������-�e>�������ŬqDV�Źа��G��Vŝ2���C��m�'�tn�EV�D�*4��|b��Ufa��̥��|VD�Y��6P�8�̀�	�U{�^E��r������
��S
�ґZ6�!_O�������\��#�|u�-��^%Μ�qV��/�9YJ��Af��H,����<9C��fr�_|f"�(.�F[�Q	Z��H��]��.�a�0�FTuȉ�>%�d�A59���?�1'�tR1��K��,��L���M�nI�c4ybi�6�E��oA;�7��n��)_)�f�8U5�6��l+������D�c�>$v��ƻ�,Y�-ũ�o�琏�ҕ�u��ʄn��@�x�+���ۋ�$��m
L�R��5�̙|��@q�f����\�HLMx�x��kcv�����ް�-P\K�~���%)"�1�:�c���f�	7^Fˈ�*{����7㣷7V�,��L��(�u���
L9døx�@*���U7u�PmJ]/�������jo�9�躺�v����NS+��X��F�w;��iN;���?�b�c���]��V~RArQ������K�:�ҿ\ �r��koM^���èi�����M��h��s�7P#��{�&�A���������'�:<�G�$���a��ͺ�~��k&�9�������	��|8�i�������S�=+� CZ솗4U4wK����k=*}wh>�.e�VL%����b��q�h������ ��X�H��?�Yq�o'�R��W�ܪ��G>�������S��2a�_%��M��V&7%�U5w��Gn̘�g<|u}���t�{��j�P�nu�+a\��!a��Zʯ��)���S�D~93k�Ёvߵ>o��KI��|Kv&M���y��m5� ���f��i=�Jv� �����D��!����k����)ˑ����u�%ʹ�V/;���FMbi΂��#}��T���S�*w�B�xpd��]ǜ��[FC=`�e��E�y;?�@�L�?:�S�̳T�e�4ߡ�-n}��np���9����i7�P��7���9q��@&0�-��c�w������yY�d���Iw��^�?��c�A&|�s��&�P�'	^�T�
c�e�t|�M����=��3�C�����-c�;��3P�����XG	�ڑ8ݴ�+��CСq��q�L�����O�-���t��	7R�ʗ��tWMg��o���Ɯ�V�DFJ��'��VЉFlm��~=ƌ)R�XN��;���ܲ��-�ی�%���s�:�U��A�#'����Mg`�~��JC���#nx
�.*(�x Eh�&fMrߞZ{7گL�[x:��ɉ�R`��*!$#�1Kl�)�#��A �u��3&-b��^%g�Ά��D}�q2����+�y�|�R_JJ�O���^�4��i�B�"�bǎ�����cr�N�q��eb�A�sI���7�r��y�F�9?�9��F̮�(�>Ӗ؊�WC��3��kx�}�+�\��ፕZi(6h�'��\?������h �c7����F��M��8:�����/]1}I�;eӹ��)ȴ� ~P�a�_Y�8\_�)k�95�|��?�w��
W�U��yFN���J��4�$�~�h���C\,P��`z��F~@T�@���Zt�V�Iᬽ�z������L��78��w��8��B=��c1?�\��L�(F�)j�<�-��K� ݊���&�{��w/��X�t]�J���|���s���{$�z���#�V�	��o��xo����,�VJ���F��*mΛw��78��犍q�FZ���<�ϰ�	�є�,~���X�AS�i���@cJe]n��bQ�q(p,57��G=�^;�V9T����Re���^��^���A��c��(㩜K�T.�q���������F�ԄE�hvg�]�OsJ&�<�6��S�%U@k�l%G�$�
��h�!��$��(����y�Hq��x�XWic���6ްB"�'�ʜDY���TO$�ݸ�˘c�	 >�(��9O$���MM`�q_	g�(�ۋs�`1c~$k�xRtNN����'�0r��wNw\���%�<�R8�I$i �b2I�,��	�TgN|@��m�ݹG�Lj��K�I�lj�Ɖ����Ԝ���kt��] ٓ�P��Oc e����������\�<'������n��e	���dp7�d�"��/��\���H��}�G�w�sܯ�	�͚X�`F�u�xiD���Pc�!2������U�kz�)}KLi'��y�C����}�r����~o���_.w6�$4�˦XYڮ1!�}
P�4֘�,=�k�v����Nb[�v®�	@Яt�{���M���E���]�� �Ĉ���py�$H��8B�7>^�Q����!!��2��˛O�Qh�.��K�'j��Di*����hY�����Z���o,�f������M��i�R�g��G��f�c1*�S`�Tmo-�������� �=�����\�WY����n�[�y���s����x���^�
���T����WH'��ea%۽7����~���(o�����U���mm�n�Xy?�LJ�/n#�Ą>pݶU��1����Mx����@���!3�81Ժ�&/���q@������ϲ��C��C>�;"�ϕ�X<e%`�v`����
\e��~��70E bM;�'�Ι��0���Pf�fF��i����������f�}Ɯ�$-$I�Nv)�������I�h@���0�I��#���p�}��EZg>/���efy9XA�E�8(�J_��k�%h5�R7d���KP
i�Mk�����+�T�R�A���Q[g͒,.�Y_��n'	'�`�Ԯ�zKŝ��,K?���dA�-��Z�9�aL`3rڵy�����M�c�J����Hy�ܪ��P�&�:��'�/���/�׀|6z-�8x�����l���[��C܇u��M��.�ѷ����w
i���������Z.U9Fcm鄀x�ˡ5C�1Ѹ���D���`\O��X/ 4n���x����.1h���	��V�.����]�zEu+5�� ғ�?TJL���3Hu�\&���
�3�<}�4�k{��%���}��tM��w�a���>kY
c7�n�q�D0
�qƫ��W�^�{�9�>	0�Z�P��E�;�9�rQ]|x�N�����ِ�б�F��<���3<х�K���W��<x��n�����Z�y������ے���c�'��qB�e�RN}�<���^c�t"Py�[&���n��,��2����\� ��5�S��ܬ��v�[��"�m۠�?��s�S�Ұc����JiS��s.��'��M�8QO�j;����{!���a�U�?Ex���u�<%�š?�8��Q>l`�BT��!#͑��ԐhjҨ���^BG���� ���$�WQȹwS~�Ӽ�Qj�h��B+���H�C��#�2��p�ݥz�x�-~L14DH�
Rf�.9`��Ò��3rd� hA�C���wfQ����MSf��M]S�o[8VQ8�/ЋͤGJZ�~D�9�5"��+��=r=�-=���d�"�)���J�����X��*������t4FWt�Kq����k�6�IE-L�:V��Lѹ���x�Ox��ٳ���K�ɷ?R9�HZhZ��x��ߑ�Cٽ�H�|鲣>�����4�'뵨��dlKr]�hSe�8��I��;L����S���*R1�¥*�G��B4�qy� g�K�#܅>e�d�� �^��������ݏ���0�_)��~�g������̽'���R�]Q�M�V�?��)�?FEq��1��~�T�ĽL�_h�V �_	��>fuS�\QE,�K�������|�-b�'m��f"�)1���?���������繵9SBsv�����B�������;k��QY&rb���1���3@'^m�}E��@�QG�'�a���7Ϳ>ҪE�n��E�;Ϣ��v����-GO��\����~��)�lKgz��.�ݰa��h�3|+��N��7��A��^�->cB��Ȧ���m��3ȥ��#O���mi����v(��U�!^�6�f��N֘ >�#������p\������&|�L��x�8=�*}�!/�\11i����[���"�*�a{���B&��*U�
���O]�Ӆ�6t�tΑ�J��ku?,z�I��|S[]�`U8�n�������K�23� ��ӧ 12{E����g P6,��5��-aWZY=�n-�]'TU[�Ӭ"�}��V���D���R���\��?� ��-�Q��n>��8l�v���}�@���ۈ}�a�����/F/�X���f�,�ਜu�fm�c7��M^�U�$�M��)�|H�D�%s=��2���Y�����q�8gB'Ъ�T [�`�O�bߡs�ڧ��)ʂ�W���E37��3^`�+2��j�Z��q1�'T�'|_��r���I�ׅ2٩��uk�Q@/&:f���-(^�_�XqM�����
�Σo�����H����\>�`�V�2�$~��g��0���xgE�_��;�;��.d�V�� ʄʚ����`ƥ2��ז�����
��5���R-�1�F\�Y��O"G`42����r�xP��c��s�E�$�=��h�g�.oU����3��D�q�e��Ne����ͱ�ӄ�#QO���w���� ��Oӿ��m����ʡșv�rX6�T�m}�Ȇ���0�9�d���0�w��b�C��j�KIpHy]�=Y�z#3�Rv���m��`�3���\�]���=z�A����v>�;�6��X.��-y��iA��Y`�7�-�ר^^�Xim�C�c���R��AgM��Z�Ʉ�1��]n�d�[�&��o�-T~������ZfUyg�/�=������C�s���T]5�ZOL����+'B��؉�ɌQ�!�a)�7��u��{
9���� ��v���� ϒ�/��LV�Ū/w}��7�9� ��_T��<������\�]9/��`�D�q��$�xO�k��g���oܤU���S��e�f����~�.�08���j�W��E}�Yy�k�ݑ �U]��79=^e��^����8���	�,ho�a�BD���HBV�{nʴ��L#�j�X�����YM�\���M�l�ЉgU�'�ܹ��� H��i�Y����,���9��#�z���	;�E U��жp��|���S(�E��<���d\���e�<�N��U;*cMq�i���ںNݽ�����v��M�Fc��_�x�����+� qS�������]������<�;(�산>�z�x���P�ǞΗ���,ۙw˨���g��S2 ����zʹFŏ�S��Vo!���o�喔��ʻ�h�
s�1%\R�3�M����	�e��Z��2��$z���ڢv�2�'Eo֙�'O~�y�'ݽ�f��A���[�4%!t%���2O�7-�U��EX?�4w~��=޿�4W�u��h=خ�t 8��o���"�g.nq�s�	�|< �62U��vJ�"rCS��sguh�1�:�ބ��8E���=HI֢�x���儫�����+�~Epjq��i\���ߛg��J��Rq���qB�\�������v�Ǯ,��
p@���m�S���LR��C5�֡��ӡ�yJ�w4��ۙ$!	��!(u�A{Z?9��"��-���[���U����p��H��´�4&3"C�X���~�!��x�H@���?�c�1�H^;��"Zts�	[*�S=v{�
/}U�S��������_�M�R���rˎ���فr�˸ ғ�ib&�TaҶ���Ֆ��M7������OE,sl*�G-��G�*�V+$��0�Q�I@�B��*"�o�^�Ӝ�~!�ղ��YeB�ݶXj�VqH![\A)j�i�Ip��%VS<�exJ3=4zR��&);�v�<��p>ЀIR��1�n�X/�mieg�ǇC�HP]U�2"Q�R�_lO��1kЦ6���r�>f0������	��L��P�#��4�
�y�_���]���,�/z�q�G/-!:���z�"�/?���8oF3Jf"⍔�"��;����}�k*L-��`������V�sk�!l`�z�uqꍇ�iI���7@g�tf�R>B��F���{�#�q��<�f�Ђ�������Ol|�R�ԑ�_��c|Ҹ!O�&ڹ���9h�ʤ��E�h��N%��|؎$k^�Y*&�RΟ�<��ͩ���A����ej�Ʌ�la��h��Ѿ��Vh������K��u8�O9�Ю�z�����:F%..�jk��A��ub�h�gi�:?R#��8��ǭ� h�:q}�'�N)��=&ϖ8D]�
��2� �����~��`c�/2>�I�!&����J��Լ��gX�^��S��}]�r1 {�����P���/\G�a���,Og�<b`R#ȿ���� ���S2���o-�p�a5�d�`.c=�R;o:��n��@C���֛����&r_����!hx_�XF�{ԏ�xm+`�!ق&��Z��Mh��={7=�W�:��i�-&KhL�x<��gA�ɠ��G���3�����J�5+e�
[GfXM�鴳�pAz�_x����\�[�96�q��9Lt%��`�$	DPj�
8DRYg�D����nܖ'��$x�*+�	�c�O��E�r4��~uC��L�Pp����B@._6szI��J��O�B�99H%^H�ֶܚ�_���Z�o"���&& <�~����jŗU=BO�hS
�Tf��n�:�h⍬��
����ؑ�dL��F����� D�ɹ�XJ0�����i3U���s�8P�K��yw��B tF7"�3k?��7�#�+ʣwd�>������-��^@�+�2O%�{�J�,�L��:�P�ncp�[�q8 �nvI��lp*��Y=W�JX�qV#J��?���~�QJ�H�)�G����Φ/�B$��O��lh���U��Zg��RsAt,%T7@���2k�)�F6���������g`��l+��5��͢P3]�0^��Z�� 3=��y0,
�Ir�E��?��+�P�n/�Y2��1Q+�ߺH�c'�--�辢a4|�u��i��yF`;���Y�7iY�n8D��cf���0��7'���񷃑@���j�����Jp��V��a}�!~n�����]��(%�B-�o�g9}ʓ5Dvji�Sb���i��ͷ!i�;`���*�\���3|G#�r�_ӗ�1���)ס��J��D�
dsf�\��������J����I!���L9��b���>��q�}�*=���x�ٮs�l�އ��dTsٱj�ف��MYO�G+�\����c�|w�iJ%o¥o�f�4؍�]'*c��voWj��B�"0�g����!�������R�����^���$"��}�b�W:�J�8�����Ί���G� ����]Pa'��2wg�Na��������;�C��Cok�Ti�H���5�ɢ�oj������<Pɬ�MޤC���Y��w��Q�
\? �H ε`�֏�Z�<~��W�Q�<�)8T�+<�����C�Ad#�s���ww6��כ�G�U�qf|;GB'����΅7��'N�4|��}6m��-�"�1�%�e	KN&1;�Q�j���T�t�z�2�c��~�1���=�\˴��imj(��"��
]�ar��a���fC���VО�s��w���p�ٔ֏�J����Z�?����Pť9��ʡ�/��=t�'6���wq���0�/����(��r����J5TY�,M�9�6w��e�X��i��e��_��������&e�&hъfo`vMl��ޯ�
I���0=�9��>�'��<������b�8�@ qqO���4۶���؂��H�g����AF<�t80什֪���<}XvC|l�x�S���7�}WQs��\�(t��G7l��MFN�&��Ǎ�S���H���#_��߷{'#K����H��.�1�G�мY3�>���Z�� ��<�:�ޒ��w}�=��+7�߄6�v��mR��T�8κ���A�G�!�k5��ߍ��ut�H^����-F����}�^G����'Eno���4/�U�o��4C7�-����2��Om0I���	xSj'Sa�E��}�r�rr��Ϗ�Hϐ/{���ٮ�x�$m�q�p�.����l����]c��������t�oǋ�Ĳm͠��g*kݔ�BKP�Α��R�L�%�C�-y��2��=����o ��vI�|{.�W��b�I���(PD�s2�9��o����B�/`ۑf!��%��E�����$���6�>9���ͧ��u/�6�Qܮ�cn@��`�����O�����8g����]��`���:�L�H������ۘ(H3*=n��B`�=�+b����lM���.ҝT�R����q �N��6'�N+�e��`����ZdtZ�TJ���( �,4
s��.GJwPs����|jsB���9.��˫��BZ�\G�|�N2��Rg~yD���B�uh7E:��q�댍��u���I!�;�������m��o�J�H
R ��^͢bh��[�EIQ��8"6����>�����ָD��ťP�E�󸢼�b.�e|nϓ������]�~E�����;IRhM�*��B�4���ޕ�Ƀ_/�#f�_�4�R�_����	�p�GD�61-��F�K�-_�0�����:B���Ёġh>�E+�渽9B4j��Lg���Q�p!"F����"�f���v��
-?��x3�sz^2�F����=c�59������2�{0Z�#��W��0|�̖d�c�JTw�5���3�ƶ����T�\�b���A��Hl;�%�؍H��U�M^qEP��$��LN^-�X�o��'�+�"[�6���F���'_������� %��h��c�$q��By˪,3GH�{��EHԠ��7,"��$�=�D(�1�b*�"�-���|2o�#{�;�"�@>�����϶�t��kX�.�F̱#:=jq�b��ZW�X�뻊�h�����'�*��;�ǃ�����-�$K�msfB�D'5��Zr���@�~1�~;�ׁjV��ᵌ�Fje�I��2���լ�f� �X���E���"���X���ݭ�'���P�ʂ���n�ݰc�_˶���t3 p���7��I�ڤ|��6dwq�~���.�0I��dktab�c {F�_̉?��<�9w)�,+.L��BU����(��D�_p�ސ,��T�6�R?�ȍ��Ȉ!>�=����g�\VN�n^�ƀ��F�G��'ഄ�����$h���*�� �O�V�ϕ0�KP6�M@]|�N�i0��hϦ
��*�n4)����C���q���Po����y���[A{OBKɊs��c�۴����qB��9��@��V�/ o�kH�wq_c� �1�,y��Jq[#c���/����������Q,m��M��uX�\uu>��O)�؄ĉ��g�ΦG%��8�\aɐ��\��3��(���EL8��uP8��M�=�����K	��y٭��x?� ��?ˍ�b����|�΢��o������7(wׯ+V_��X�K�q ��v��=�B�4���V��ϓ*��穣��Ŷ}7���Iu�]�M����g^��j��]T��A�9�MM	�%"��_u�B��k�O��K��7�����ӎ6U�JY�?S5S7��MV�C��ʵe��ţ���{a�Ɠ�BrIvs�}o�V�"���Ώ��b:7���.�	��/C"b����9nNx�S�4��v=��J��H�Ԭ���!_�.A�":��z?��g��A~�|j	�d���uƛaE���Ɵ�w�ZaE?�M3,6M.��/�Տ?9�o��sZV"a
!�!}펚}�ؗz��Zlwl�im)M��>�9�y�<�G�H���
?O�8u��|�7A2ֲ���i�0z�j�{nB�c�G[#d��pE �T}�q'����Bq�~�M���&�J=e�|H��%F�{�R�q�)�����"QK�|o�!�C��g��d0a���Պ-���-J<�,�v-'�����9$6!�gߖ[�W� �����r"����2���{����&	�$�ZR�Dn�y�$�d��d� u���P�C��~����(��OX�T���s�I��D׾ʞ"d�=�1ɀ���7���~t1["X�UVM|�mN���sR2.�x�����J6��Xe��z,�A��CO�qT`J���LË�4Ԣ�}�n1��o����U<����QwF�\IT�&+�u
�C�QG1탾 +Ƃ�1��6I�-��Q�Z<?�p"�c�����Z��ﱝ����L�lk~� "�T�H=�|�v5o|�6�v��	�a�	��*(6�V*��[�y�	������#VX"ۤ��I��#�����W�L^�O;,�H�w�(����*�$����=�X�"�ȁP��Ka~���w��rs51Y��m|��4Ĵ�o�56�~���q��-��B�a����ifB�)�����N��W,�s$q� ��k����;:ա���(E�ѷ@�]�����������Ԛ7���uPZ�$���TWz��H���kӾ�
�Tݽ�|��-i�Ey��ٔ!u��^wa�	A���V��v;y�o�5������9lA�M��럚e���l�>^�\���z6��P�##]![�=$3H
�bԐ؉O,��b^۴�q�RD��#<�zHoAb������t�9]�	b@'�g'+c9^�6	��9����At~�F�b|��g���� ��K�����!���V�i���,`1���n�4��kz��P��p�\PW?�m�4��b�Iץ�Of�j��e�k�7Aي�?	���ך���q.Q������=���O$���o߃i��
���j:Z��ВK�t㺈�R�9��Q�6�-7񕙱e5�1�7^%��w��D���Zxo�JZc��/b���WΩ��7=߶��d�xuE�$�!�3��d��"�X��v*������@gU�x뾄�㼉��4�kS���O��i�.���P/�&ԗIQ?���J�;���4��j2A2�zZV[�II*]ARq���O��8�`��)/ %�ܰ�Ϗ�e��#��X�� !�;b�Ձ���_n`@�8{1���F~FI����۠z�-�t�f���k����lőD5�թ)�?�Xr�?qBb;6A&4yy�'Pu��:bګ�5������O3�Lx�ma�k���睓�F�Z��@պ=)�!	F� �w��&�b>����&�2ϊ&��R䏵���`I�����Xb�#�5fTӁF}��Zx�j�����
I�N=R2�6�*R��U�^*�|��f�!�՛[ ����|KˇPV|���Xh��%=}]P�7Ŷ�Z�*i�4��A�]�4�������a:�����@�S_�hTГ�b¾zC�W�X�^���Wl��_7NZ'htlD��F�l^/����@nN�Ҙ�m1��mSǒ�Ӵ�1u&{"��$P4+-.Ӷ�̉�#���}���=��^%�`cQ8�[C}t���(<�<ſq���6̰�&՚�x;�ͭ
�h#�v��r������Cd���
Mծ���JG� �� z�"�D�������"r���:�H��·���;�*��:�+T���x�ຆ��Tp*����w��N���b�0�B��7Zlr�����g%��l�mu�i��W{Q2�SD6� k1D�ۿ�u;4��*����+O�]e������$���Q����GI逃���'2JCz�7�X	z7�W����4�~�_z��/�ѓ�I9�
b�o�����p'>ǎ+z���o؛��\������Cgt��GG��䲆VCG���'����:�H
��4t���fkz�ՕJl[ٻ�c��\/�u�Ձ!ZKI"�І�,�F��;}�W��<W߆G�E���65Q~��D��y�mg���Zkѥ��[�����)���T\jT�JZVʓ��&�ʨ@ne�D"��̵��+�-9d$r0�Jf��ƴ�~�<8�����_f-��yLN�J:!}�O�|��K��]*k�N���=�!��9E���B������%(@���kˁyKjN�����d�	���J���y+�(�ѓY��ȫ������ގ�*�[`���68�v�����g�WvV�ո������� �tI4�w��yϦ�UAeۉbN&�FxR��������S;��qؕ2����)���i@�sϏa�v�gl*+��U��P襩��5��35��Ld�V=l��a$x&�zq�6LW�(jݚ��B@�ѐ��-a�!�K>�%S��y7�hNϛMC���ָkH��%`6�H���-�s��'0I� �E6hE� ���$(q�]�5[��͎�Q��gOo�!�����k�`�]afx+�Du�2��]{�h
��Dd��]�RW	-�ە�#C�u[�L �!�����I_
7ث��U#:�������j(���<!�m�IR�y�$8�햑J���1�!�ϕ�W2���Yn��׺Bb} %|g�P��W�8��c���&��z\3�H�;,���Ԣw�ņu^�Η��W^�qΡR�a���Yӂ3x߷���?��'-hA֛HI@,�i`�m�:��ƷpA�ϾsA�Y��R	?��H���^��vdz�^kǠ�9
���Y����>�z�`���<4V�(^���Kr�($A�"����٩c�*r�TH� N�]�S%}'��z��Q�)^Y������M��8C����p�A��p����y�3#�k	���0��'�d�2a+|,�R֮6i�a��퐒�O���_�t.+��ߌx��n�f��#Uf���s�7y�f� Cv,����7�"�e���ՠ�fO( ���H������*�+�k����2e���Vh�� ��&(�J�֪�ܛ;��<�;�	��Nq	k.��:5|��o��3�F�<wN�\̅ɭ�	�K�b�.��<��V��v����Y�b���7!=�oC��\#iۺ�2|����R5i��$���NO�*2c�
q7�}�����L��my�ۜ���_�Y�0{�թ��ǎ�r�Q��Fs��֟Ϗ?8�WDKg�jG�\�驤��>��)E�>'�<���`M%�j���9�N�9�ϑy�1�%���!!�) �d_� R���%��:���O�/	#�=G@o�b�ă�"��Z�ܬk����	��^i��2�c�X��b[�:�?���u9Fc������ĤF���BwA<��]��]�,2|�Xu�\Y�l��t�8�wB�B-�K�gPi�gd3��37h>�i��q����Xh�0	d�ב��xͽ"�	��1[�t��@�g#s%�KnFz�5v
��V��H��6�+6^�;s���Pܥ�H�0�E��xh��S̐��م��~M���YigH~���;H� |���q����w����Kc�c�'�����ʈ�sE�2�Z��1�$𣔌%����?5��f�S�Xң���߮�3����b�M�](�3�^��
��J巟ڝ���O�(�i+����D ����y��PGU�޳	������&��K�vL�i��Sbč�O���s^%���I�����mh�7CL⤳��Ͻ��s����L��P����A����k@�7�q?W3�gr��^�lI�8�ϗ����x?���*�=Wr'�_�	_OݨgS������#"�3���'vv`%�z��.�4�^
�y�D/r<��l�:��k�nh!&������B�B$���/��r��a%����p�C����� ���iV�x�JZ]���i�e��o�Kc]ES�Tn'��ͻ�k��0��w�;�V�ߡ�]�ǎ[ �1szKo��Fq��z�8�	���q	p��U  >52X�9�3������d'�&�V���~	s�N�;vE�Y%|�s��J1*��E�u��Z�}0��A����/Uı�lO��rвq��(y|���N6O�r}9��;����p=2%ï��·ݱ�������w��38oQ�D��V�o ЮPN[3��]��& =�8��퍺�`�F���N�oh�j�[�H�P(���d=h~� ��k_~N���D|63�X�Z%޽1��8�U�]3���k!\�tȨ�g�#�NZ�8�'|_�M+�n���A,Y!65�����J�'_U�+x��ؓ'�j@"�4�םA�!\����߉���۷�<�pd�rN��\��2}����I�l<I�cb|���9��cZ�3o�b�v�<�X��*������F�,DF>1�L�T~*��xΙ�
ǥ)����'�S�_�۱)T6�)D�vwW����@ʏ��)T��{�]�1������郶Wt�mNH�3�#�r ]��p�07i���:]"�t�)j�B�� �\5�R�fo4$,�����a��m�hy�D��Qek�l����h_y�����|K���ӻ�L����7�+��=r 8KD5���:����;jD�c�R�N%��6o�W�x����.��a;�aV�W��膇,6·�!��\ӥ3e��wf����h��X^sb_j���z�gg��6�\���P�OC@Ǿ�J������+m�փ�༅�J��č篢�b)��m{a5
˹i�\)�jp���\:Ľb��|nD��/⿛�L��$�����.i����ܳv�v�����c6�KOq�p|h���J�Tp��P3�l��{��x��N]Yz��M��.�[�-��R�9�GH�V|������ɓ9J�_�/��J��N*��h��Ov���ʒϿ|B���;�u)��ژߑ�Z/I	w�:��F3�Ϗ��(��Ӎ �c��	�X���Zk�O�%�� 6����Q��~R)�6���0Ic9�A��`��	xR��"��_D(*�����G����V����]�@f%�N��a�DY+�j�譔�s�-y�=�ђ/�QW�VD1Gp���Yi�To���W-�{�?��e�N���K�;�!�Eťq�r-�b�G�6_���-��ɏ��G����l5�v5�c�� �bĴ�	K�~I>������
���������q4	aש�I�Kv�Nʢ��%��7�ن���� a�����J���.��͌E�P(�}���}C˞��HA��Q��y��)�8�I�=+��޻��K���+tH1��88�oY+�6D/��:���
�����0����t�r����y^��e��)?���t�U-e�9�^eUY��,)0�M�b�Z��r#aZ�LP[���?Ǆ�czkТ~-I�5D8��:#	���G�����O�tGH�'�o3���ӅW\�\&�g2������:�RK{�>-6�fuz/�T<��Q8�Tfd�>�[�b��)m+�b.�֪B�/�p0.9#����b�|��U6�غK ���/��p�=A#U�4�ȗK��G�v����c��������������&Ú[d�1�p*~��� ���!�S�p��E�:�.4����?�=<,�#6�\�� xՄ8��(ɂ̲ĂJ/PQ���d��b��6�])r#xh��k2�cP�Wh�*�
�P��	
���J�����O �L��ܺݚ�|r��?x�'ú�±{��lk�����F/��l\k��n�����E�d����t�J��y��}�e�[s��^�x@/�E1V����p�4���E��?'�5e)�J��h���`���n����Ă��ʮ�$�ȧ��w'�	N��N t?� qS�,���h���|�܉�o��J�l�o���ņ?h]r��3FI55�f�v��]��#~���z~��SO'���]�Q�:u�)~.(p��TQV�-��Y�ύ�`ϤA3�t@���̂�<�h�Y'MxxA����mFW8 f�J��H�6���xF��>"�nB-hBa�G	��CF!�N��
_�+YT�M����o�<��'�L'J��{�I��4V�rc���&-�Վ�s���^|����q#�NAǜ����g�S��O)����׫��I1�MW?����&�_�B�#aX|��:%G`nƜ~tUҚD"�؊��'ᑚN�RE�e��sц�BՒd��uuYVU�����7��5�Ud�k��̮gƉ�ZF"���8��q��f,zg3gFi�{��W�~͂!ǻ�%Ӟx~z�t<��v�J[4�&r\(�����r�Wc�j��zɳGʜ�o\�٢\[Csy�8�\�M�B{����>F�c��Z���TO	qϏӾ0"��T�5�QID_}��$RW�]j���	�	T�t�*D=)L=�'꿥��/,B� @�)@�f�vq�FSйgpa�~Fa��8�ɼ�P�����I"3Uz�ϙ{`a�8U��b�(���V͍�W�զlr���>}���D�7��u��D�@��Ր1�ӹ�<l����7�@���b7:��W��(��09���p�9��k���r.$E�Ń],������  ..�y�B[̷�5j���d� u���̄;�s5rf�/6������Vx�
�v��S.�Sļ��8:�������@�h�\U$��a�=�OX�n���1kN�m]�p�_��lrq�5��PC��D���@��Cb�T�#ޥ�|k���ْ���d�g}�2�m|���i_F��gրgE�������͸�aA�s)G�j��eb�ek��,p;�R���m���#M�X�������5�V$8���F^��>��Ͼ5�c��o��,�vJ~�f�Y	jW���l&D`S��0���.=��������r�PC���3tPJ�>s��o�=	&.���l�@��ATe���{�ŎC�dw���盿+�����ݴ�D]�_j+�+t��ѩf%~�(��;� ��ߥ�k�?���^��g���E�.Xή���1u'ٗ����5�����PC	K�'�:�k�&��!Ӭ~���N{�J6�A�j��)?�;u�5uBR}]���#-����w;73�����~�WN�7�
	�+(��
R�b��d9�=$-ŅҍW�&���s�Z$�5V��O�BK��4V��#�]>Wr�E
��W/��3������-w4�@q%���gj��[�[�w+�KE�u��v�=�d�S��R����o��=O���:�/�?&,LdǶ�@��v̀�G�Z���_d+���������=��¬rG�)iKRn�`p�1ܕ��F�V�w�؆�A����8�����Nt���)�y�K����D�c�[Bw��ZG[�Z
����*k\"G�����E�ZUEE�G�j&�g���LŀT��YM{|��-��zR��y˓�n�<��Wl��k����n��ćϨH=�C�0hvGu_�v9�w��+�՘�Z�,`.�����$�tLSx��X"���:����M��^8��S"�bDz�c�H��h/|*�	����lt� z�T����l�E-�=��54Z�.�5<t)���a�5Y��|S�ʳ�{� ��⨊�]�<'��{&�u�í���l󻂻�3cM������ų���hㆺ���WW����i"*9tN�Cݪ�h�6��I)j���@�%,�n�p~v����!A����Qr �j���4��*N>#���z>�������H<)���m�̱��u�k���\4�7@^�w���k���򏾣�l6�S`���sF�-�Pӱ�F�T A]��n98u�����7U ����j
s�z&�� ȑ�@s�YT�,A�;4��6bN�u�
6~�cH(/U�#y�m媻�mi���!|}����x��4���3@���T0 II��5��I*�2�v��͛]�}�c�7ߦ����I�MXu���ͯ(�{����!k�>�||S��~�|a>�x�%ڀ�B3�pt�L���<����9�2�"� pp�DY�%Wj�J�}�-�"�j���7�i暢�*;����uU���0���F��Ҡ.��zS��V1eP�u^�����wj'�4=�"҃^�LLA����/��R���<�؎>�,k�=C�ʥ�{�i�fB����+����mDV�B�%���@��-8�f�.�� �}TqJ7�����zC6xGfb�0݈
hX&r>a���-s~�������S+Pk5L����.�ĵ�ל��X{sȯ�ɏ0��}��%g@Q-]�09N-gd�݊m 4����Eu?P=��x��or�#�8�ӡH ��h��}e�����{�PER7�n�0�*��-Y���*w���AU��.&��:���������L�<��1!�;���k������>�$8�֥�R�^n�:��=G�	?i	2�5�.ˑ���Rxk�][L���|0T�0�8�5�ՙƺ��Z���<�V}�E�_�HX��� Abp���R�q1z�!�'�!�x�3.	�gM�sӠ�g�pr��L��S��Y\����<I'�58����u1)�'*�KN4�.y�����ܑ.���q�t(&'(X�ѡ�ќ�3��4�f�-垻 �4a	]��R��?#�j��հ��K��ӖLP�a*�t+�|���C�y)��Y�t��]Dy/��)�jy�7��{� ��:�v7W�/G���(�i.�DeQ��<�nHyX�E��d�:��v�;P�Ow�pG{=���A��L
�)�a�c�i5�R	%eީ�4#��-�� w) �S8��|��N^7��4j�6>���S�S+H�~?�;��&WzV�rfɋ7�;�C/�P��<o�P�"p��xy9�p垧g�B�B<�[ƭ��T��ɖ���Yi���W쏶;�,L�2�#-;������������o��!-bnL�էࢥAI�V�gm��_@dJ�&�Y��j����	7���Y=p,+�ҝ>a�@�R�c�UG"��D��7={V6�@�lr;
�ɥ�.�tY	��k"�����egߔ�θ��mM�F�8���9���o�ܸF����syzW��Ep�*����g���C ����~�%���HL`����I[���B&'w�]�
Oܲ��h�.X��6���O��R�$�$BD�zx >=�D�#����TK�:���u�m�ϊ):L#zb�p��(��]usTb��2�>i������խ_J���.�B^�)6��IH�+�yVi!��|�U��]nѕJFq������곞�gm�x��}f|�Hc �忨�֕�o�kCv�q�w�ё��'ҸS�o,1Q��՟�-�*v��_^/�b�H��-1�g~��҉U�yX�s����#�2u7�F�ѰSW9(���dE��nT�o�iN֖`}�����]bd.���Cu�5����,��6�FP��,�c��c�q�|�ԛV��@�(�"����ɽ��nϰ�L��	��ϗg	�~2N�T=�z��F���N~h��	��;�W �Jf�h��K&_)[V.ت_*ev�0o�w�ҽI5XO�?��L ����#����;dU/	�d8s�ϤEz��v��:?RR�E�!�h�!�"��2��f7�\XG�J���#��\O1��4�)&�.I��#I�R|Xt>�������z��Y[J���``Y��w�ʻF	�Io��qˊoz��C4������I��0~`j|����Ii�ݸ���`;j�l����:��NSkhbv:dW�V�9����2�"|��&/F�����p���n�i����ʐ�萄����s�(+��j�sb�rG��)N�7���?�f��'@�KQ�� ڿ�G��=+h���+�:ש.��H���>�]K�3�5���V� �o��ru?�����)�ȵ��,D�=Oʖ
D!0���#�`n�q�N��0G��-*��i�����v6E�!d��C��H�[�*7���D���{�#��6~Q9/m�jK�~kښ}��`�e�P�?4��2k��-;�a��F��[tu!��~ڙ�����c����S��c�ʻ�:�760�2cvJ�L���Nv�����K����"jR��z�y�V�[zl�\���U^iͥ	W(����x'@��A�L\Hm�S�B��|���v5p�B�ntr�T�j����#�e:z�PR�?�N��&��i��O�`O���s1Z���oE�8�c�Ȱ������"�~;|���&�4�~�W�� 0�K��:�j��x���������$�6�T�T�R�[��˳��c���m��"�м<��,��V��`?�W<V@#ʬ���mRV���K^d��~���w�b(-�������h� ���<Q��+$}�a��7d[����*��&����OܮD�p�+��;�����!�;���u
"�Z^Z�H`?I��K��₌�|}�5��`�L����{9��k��j�?Vhj	�X��KMC`�1�3$��t"8��ﳿ&�V�Y��[x�Jj�;=���ЖL�s�jR�{�_H`��w����g#;!Ԩ%�X�n�i�Ԕ�MHj3�t��ws�e�U�a��3V+k�">�2�	i�t�&�@�{�$��P���m���c
�r�� �^`��yd��'����o�;��3̔�y#-���j4o��>�U���p�e�0��Au���.jΘx�4|2��d}�,v�4�;P���>��dEE��T�֢,�2�^�@�,���C@��RD[�l9S�\�4�1�H�����=(,	������%��NtO?!�1��z�$��FF��`��ڇ�����YQ��ǻt��0�R�c��xm򁫆�U��M.ڏ(���Zp�aF.ZD�D]����r[�X�y��R�:�Sp�H���Y���#oyW�Xۍ錓pn��'0�S��C��T_ ����j|χ���Q�⨔<��-�VQݻ��ȏ|pZns���rV������p�p��!b�iǒH$��7��苝�-��}o|)�'�(#" *�kM����X���R�<�q�?Z$8�K�C>�d_T�%^5�+(oxH��k�n�Q��h��m ��3�q�������2��k�=��Űq:�x鱂�Z�Q��B� 
g�H��~�K�}dVVeE���x�1�]�[���T@FY��w�Ȫ�4���������Ҿx_�(b�w�'Q(Y�����V��(se��]��e |'���U�\�������t����^����T*�r��O>�`Y��;�f�o��5�n���_��]�5��`�}Z�l0��<@���C�gCK�mx���Y�����D�6ͷB]�F#�:���Հ)�LE����~f���1�a��%�l�������O���uO	8�`i�!�Fb��yc�Q�/E__�cc!��
�O��&y��D+VJc9����E�-��5����ǅ;�vߪ��R�����M=�.��Vr&�J�'��K�>�1�T~k�J����P�������%���灯-h���q���킳����\���cs�̿缼�F9SkAޒ+���e��7�S�Ν8�S�YEMB���}����;B'/�j��~��$�r`��p2���(֗��03*��p�N��(7d�8�LSa���T�G*���-��/˭�L]$`Y�b����/�37�4��M���d�h�dЯv�Ҕ7�Tt��Mw2�x0��J
&w^�Кi�^��"?1��-@{Aa�)z6���{i]lԌ^���a��DI�c� �z ]f�����r��o9���K5Jle$�!!'j�ͼ���DАZi>�gk�"���]4��JN#k��Kǔ���<�O�^�:��pQ�wyI��f0`{�����Fj@]�)K��3b��\S:�.��8���
lL��u��5ej�OH�J�&�anXn&�h�������G�~^/fo���f���S@-�E;���$�M�)�5XΟZ5M�}N>Y�'�8�Vf�5��kN��xB�d��Y�!ig����ͱI�\�\�G���F��z�z&�^�>��d�jy����3h~Q�~	��Y��p}�&	��s��>j�����s�AlC�h��!�����$54�Jh8P�-ѡkFOB���|�浣����L4��-�����qC�������V)ZV$E]�`��ݡD��	���e|��oXk���,U�n���"��f��S���q����>1���!,�v�n7Z*�;&Ѡ$ŠYk�#__V�W񸽷���5��5��m�l�(����C��pBx��c�� h<�2P+1�����[^+ʗ�T�2t�]����j�� n,0Fԓ�7�"F�aΚo�",���0�#�E�d��I���u]*�
��Hc�3fW�}�B
�~�����i'��3�bۭs�5~��ֹ�sH�׻�:�uFL'�<�3���T��m�St����Z�,CA|��I3�9��9����NC�޸����C����������vs�.�{H4,�Y�9e���e�Q��jA���H}�#� W��o�ExH�=6�c�!;�!�Ϭ<�o�U�#r�V��7�fd�% xYj+�!�Õ���_m��Z�-Aig�Dy�hv�_Fu�{��BN�R�%uVڂ��m��ҁ�'�匦��˪� '�;% �7��Yۙ/��Y&?P��.Y=�0�Ě����M���B���LT�A��^�V��䆟��4��x��$�\��k%K{�n�㴃7�u��i��vfB�GQ�~��ϝ����.�����W[T�U���-ߩȄ!0BB8��OX5���[��sd'��o��)�*f�I:Zf��VlCJ���b�)�&f��rĹ�.R��(La1_���p��r�1P/Du���6�u%���լ�x���$��t̿vV����&@����'BN ;�\}V�t9W���@�1�]/+�e.g���0��N�`�,�U�"�m�].�&h��6��ǩkO�n�4	!�/�q���C؛��iO4n�bD���u����B�!KVֻ��in!Wܿ����
F�U�>o�Ѥk���l��]]J�wE�H�E���J/I�@ζ�Ÿ.�ş�lm�}[}���Qd�.K�0���f���t����`p'�gj<"� ZV�^٢[�js|[�
-e3? L�c��\��|۔��i]Vnp.��61{��j�;>�H�Q�	y|�>Z��� T����5U�s�9t�˧�[��VbH�z���B�I�%�Sc�ԯ�6�S��套6 �8hAd�{�K�����?���е��u�Xރ�*�ךaV�d(+D��~+�7�t�m5J�8�!|�®�*�����dv���������:'���~\r��A^����T�$���9�%QŨ�K��~��,+��^|��NВer����z��r��Հ��ߗ8�C��z\�YI����ƒ�ez�L�b�6�K)-B�XN���Q,VQ���F��P����M��^�,t~�N�ּ��ڴ᧽&�oi"i�$̰��b.��֎=1�R�	apZzK�iXW�8+L,�_I���;X��6K7��)����N��������7$� aBj��]��^8I�	�ه&*�������IZ�4��]�����~j<��v�*�.��ݣN���gG0x��i" j{�:�X[���Z���,g
�e\����Ն8"��v7�ߪ� f"w�dY�G�����|L��M��p&�J�P����S�&;��pN]���?rcD ?ҕNB�*�+������㇍d��������\B�ȗ�_s0����K�"-������Z�$�wO���+��E��=h1M���͸zH��8��<�W�w��i�9S��ّ�3`�/�&�us���}K�҇)�i�1��B�X���p��-
\�#��[�e���J"�^�>��M�3Ɇ΀���c�&p�	�h���!Y��-lB����a&fnw�,��y��#X0�.x����g���ĝ�p�L��.��.��ٹ��6�L&A�'��2�Z��=*x2�`npE�c5���l��k����3	���SX�o�_͌��~ʢ���n�Q�\������x�9-�;1��\��N����5m�	(��z�꡿�}��n�8m�vX�rOU�����(�5�-�wdj�	qa���7
M�_L�M��<���
6���5�T�ł��R:xR���k.����%2���,��'�\���O�r��oջ9-b/��$��}�ee�� Iq�V��ʑ�K���	vS�<+I\R�Dq%�#27ͳ�s}���{<��t��+�Dٵa7����3��ð���1��j|h ּ��|I=�B\<��yTK��f�Fn�����$������51��U��&qX�P�$�b7���i$���PjwQ2��-h@����p�B����S`�?ī�tc�q��y�>EX��<S���>aS�5
�`��u����K���[�m;r�\�G�_�:R�M���a��/���s7�^I���R_�f�H��9��
����Wb�Ƀ�$���
�^-�z6�[��5�
��Y���_����wԎ��I�m�5�ImP�g"r�\c֌�N�!v ����1�l����K��A�D�^�ϯV�Ϲ%�S7]�@��1�� ��!d�i>jR1�5���q9�m�m�][Wx'�<�,�����l�_F��h�m�W��">]cW��V>RM�{�	�ɟ�&2��Z�z�Q�B1�G��$:�0��ꇺ��<�뫫ؼ�M�>R�l�І2oŘ{��Y,�-���w���oSX,p�"W-WH�9-i��iI!R����	_QA�g�3��q�q�-��I�K�]�~���L�.9�	�QnS?kJl�.94	��j>�2n�0Ś0���V0�ǻe!���$��ԃ%D~E�M��⶧���hhٌf=����t�u�^$��}yIOC�4}���W;���q����C���l�����6�,l�P�֕Ere*qN��+�B��	ҝ&�x��}�?|� ��$/�ԁ�߁�4��.x���2�����^�H|Kǡ�χ�� tu6 q��7�s�m!Pa-m_N	y�(�LKh��]���m-��}U����������RV*x��2b���	#�Ϝ�j��
���k�r��7�)���psh�R��2| !��%�xO�3�I栗^,�{�0�T�U�s ���k�8�ڋ���9E����\,���΂Z+P�~YR���3��.���3*��QۜO�|j����2�5ވ��jΕ��g�ͯHm}��W����HFi�O�5p+5�&���SR��[]�ˤ�$��T���kLe�!(��UA7dH�pA� F2Ս��q�ܝ�M����$��Ӏ& ]��
q��V�������a{fm灋��u��ŉ��T�z5oI�}�����-�Q«d0]��˳z����t�/�J-Y'�hk�W�*��ϼ�cV<<.�(����z�MXEy�8�ۢ�iՔM��/�����2�KΩ�8s.���1,������"�����]����Q����v������U���O�F���Cn}���J��c�~au9G�2 ́� �L�~c�A�s�`�J�;p�i!¹B!�E�'W:��������X�k8ۍ` e�VB�BJ��u܏ҡ�±Ě�:h�����K�?�~-2f5n�Y&mK�S�=���fm~����l(uJۓY"����*�ݹET�x!rY��>g�F��t��o�BNt�]�s
�~䂒f�/���֢*iZ��YEh_����ͻV�l0��Go�?��&ÿ�����D�Ք����[��a�:9ˌ����_��= ���5�?�V��g۸���Y��)bi��Icpb���:���c����o\[��u[)�$�EA���Z8�#l�~������G��8;�:��~T���ؾR����gh�`	���'B��\t
e��u�̧�Qš)�Q��� g���=w�l�:�zVe�k�HZU�.�S����#���r�|Y�fƍ�0�� L�A�Ɗ�
i0��I:���t�:f�+M8�� ���Q���FǴ2�.��ݭA6u�d�P%�֡��X��&��K�	��͎��(3ɮ�N���?s<�G_3R�>C�.������Csn�,�ER�'Ӟ���AP�y���F#b��Tߗ�g^9���ˊ�lN�UpR���d��ȿ��#�����/����na�U��c���p��w]>�&@@��ƆG���ts="�X�'c;�����a���&d�����a/�VH�]&K��9�/z�x���0RK&�G�@��OK%�q����&���S��Ǖ�޸wK�6�lŦ���m<̭�w�z[-�՗���bp�1�"��:kf��{���g�cW����;��dQC������B]���;p����H��~�32��VW͕J[�:���t�F-p��ֳ.��dY&� l��#�ʎ��?Q��/<Y)�����59|M&%JM�f�='*4.d��L\0z�x�s�W�����Ns|��,�>(Ƈ�|�U����XF���}mA�_+�I�@��o!Ǎ)eo���}.d%ݸ�}jdO��Y�L���RhJ�_�(¤���	�3��l,��}�Q�aW�4�q1�"B��������x��uǫ�d������,1f��]�a��cn��TRr\�F�D���w��1� �I� ���H�o��:���D ��Ι{�`�<��L������ٗ����h�{ﺆ�q~����R�y��]�-	�t���3i�Ï�Ī��\����Ӫܷb������_�T����_\)�њ?����c)݉Z?��R5�:-䷁��q�thC��Eb�4�\���ba����q�m� 	�-�T���N��|���<j�$)n���(
�3X����U���M��fIF��t�o������m:�ET� g�Ũn�dU�BW�_���&�eV�����!���	�����o�N��ϙ+�A \���R��������"V��s{��y`�Z�-T�Z���o�0�	U�C̎�ח�Z�%��\��	7��lYC1T�!:��vPY�qŵ�Hء��(V��Ut�0j\��8T�i~����iZ�Ⱦ&5��d\�F���W�@�9�B���|�Īc|��|TZg���=zh~�o��B�X���FJ�34q"����&.���77dw����^g�8�:+2~tʂ9~2I����Y��BV�ߤ�`�@l�|��K�ħ��&
Q0�[�����**&a\ς �4tg�!S����
�WL���"�d��m>�݀�+�|����h��,u4�D�7�sNL�s��֙	%� �����8���π�[�߃�I�[xGL%r��L1d�p.��Zg!ހ�w�l+��AP�E_@0�}�9mMMj9�V+��F�8�8�"Dtױ�2ŝ�"�w�Ow��?}���֍�o� �K}���9x�i��b��äL[_���%�@4ӚE���A���Z)��p��^j�d֋󅿱��xO7�?=��<5�Տ��`5�;��PlB$~��� (��:���
��/f�\ʷ��5�z�n������q$emkZL�O{�>��g���Ӛ��2R���7]��N>9�Eu��*V�,H�sĽ������Ӳ�=ēX7�G�W ���x������B��]n�e���Ԉ���=�|2A�d�,�GF�~~�w�hnsv�IV]d�4������\)PL��ml��Ź�<�PUq��B1<�Z�S�IΣ�~�ݞ[0K�t�����2�Mw�iE�I�Ao`/Bi���Xp�Ԕ�-b :��R��+َ�1	m�0cS�n��>�@�/��L<J0l�����|�~�y�b���oVpNy�y�bP���� d$r�e�|�Uq��hqO��,��l`b�����2g��і�_��IE����'[�8���W�u"}nmT�
�of�i*%�K0�Qڇ|��{��@�'^��K[��l]�v�{�P,����"�����D7�	w 2^��ܬ6>$��J}Z	�U�s{W���[�m�Sd�C�׋����$zvF��ҝ|C��@IB]1D�k��4�m�� ��#3�z.��g�1\�8���m��"ϿB�1P��{F�v�*�+�J~@uujj]<L�3�� ��z��dq(t�=�B��-!�b}Yx�߲��N܎U)P�G�1&��&��e˒W��~D�d����K��~-1�(��S�ok��a2����S�v?W���}��<����)b�1�P��}���-1�[N��T{{_n�5��6���Pߴ6h�6�m p������'\.�_���rR�,���1��c�&��v-�(>���@�fN���![��R�H����N������"�4�C�*�©d2Y�N+��US�j�Eڏ��d�lL�/����D�
�P�n�A�jw$�o��+}uu��(uO�����]m�b;{т�f]�[�G����[�#@����y	�Ak�nә��w;g���x��A ����bRe���̞�	�&)m��o3_�Ok��[�I>�K���i�,RG�4�^UF�n6�a��	s��k���뗇ݒ*�ԯV�;�y�6_接w�G���2�ES��\�	�0ɰJ�����b�� �O�;�@�
�^i��MR&O��Egb��Yr?_I*�8�o����$>�ӆl��y�PG�L�Ԩ��+o�]`NL>�4�h^�+!$��޽>X(��p8M�~פoH{➹���Y����w�ޠl"n̼�Y��s���-qˣP��A:�2���yܢ��DZt[��3���� �W�_�4I�".�=�Bh�gb� �0�|����(����},���4a=,hd�ݣ���d<`O�x't_����e�;���2{&׵��j�cqST�t$�/�t�,�HH�F��W:��<��R����^��[=�� �o��5��t[�`�~�b���Z��%������R�Af�|'n?"�o_�0�����d�[���e��J�[um_�S�������\�W9œ{NI)�	}����<����/�G=�!��r<L��YJ���6U?>��G}4��p{"qU�Ų2�a��h�.P�3fV�H�jSYWv����W:n���葳8�*f�<D<�ևמ�*�uͦ��������{C/���t|���u/�L`��L�<�*�,<�t�1/�7�� E�\/tx�a"�$�OW��(N>�����<|]۰nc��.O4VJ^�)��^	ʅ��]z�:�r�b)cR�٧���}�i���O�K�p���Ֆڟ�ff`$[Ja?��'j�&��(=f���D'��WfK���A�"H��h��L#wGD'�%�%��>�+�~�R�#2�MgU�_2�
�쭰��i'��K��݊���ӜJG���[u�P���>���Į;RܦB�.�a&��k�#��Ǐ��3^p����И��t/��"/�}0����n����f	�c�Al%܂@T�9��q"� ���8�XN�a��Y-Qa�
i����&m��h)�����ՎER�s�Q6�2Ĳ��_1'J(&�`p�6L�Q�Z��f#���-<;MM^(0~��kȦ�9��9���c�����I���k���um�IA��X��d�U01�BB`r�e(��q���<�gey.X���Z�s��wA�����$�F`X33���B���(&I�[�Q��v��6��Uq^��z�B4�a���I�ɽ\p����<���Go)�����[$D�a9h�t�Bo^���wx;��0d�;@{��z��.t8�:�K`Ág�����z�|�(\EA�Gj���������{ѝ�SK�,��`��[� �!��Xq��U�p*z��R�y�c��ɓ��M��S5��j���v������u5� d!-+��x�5#v��5?�fղ��)<< ʠ�8#�Ӷe��8M�`�+���yͳ�� ��	��᪗a���
��z�{R\S��?�J^��9e��@	7�/�X^��z]j����K�|�������9��Q�-.P�mV��#d�!�8ф�$Z_�1�92�M��q����P�ׅ��ivP�U[I@8��s3����@Յ�oԾ��UѶQ>��r�e��G]@Ġ��܍T��}�����r�T���-7�	�Z�lv�ϐ�t n����˘pi���_NmL>�p�$�/��I�]<���gucC�#�-,q��>�~��ݎm��=�̾(���+�ر?F��:���c��f�3`�)ivQhT�����ؐ��r�n�^��L��#�������V)Og�\�>4��LF����U���lv����R�h�[��kF�j3�!9���|���JXw�s��o~�я"�)x�G��ReR�귿ѣ�k�b*	-�e@f�d�+$�E����E0{-�.�=�_�5g���&I�=}Ɨ7 Eb�ff�XvLY��	Q�XZj�~[o;!MQ��a4�̽�	01��}*�7�s�)NYlb}�[+jp>�fχ$J_����K�}22��08�ә~��L��`_�8x)�<0iC��E챹��+9�+���k34��ܡ�x_����	���鞃�h�p�R"\�hw��g*�H|VÙ�ک*h�'\��#�����L#�yF�MIB�mQMWnz눂�^o���� ����w���F��
�����g
�H%��o������8\ P�!ap�z~0�^b�<g�~r��f U���$�޴X��N����|s�
��Y���~���IU�1�wLt3u�C�:�JW=�Usn��͗��I����AP4 ��J���Mm�鞮!d��D��*����Ϸ�]�n��ҍ�lx=j"15�DZ)W�(�&W��D�u�f�מ����D�L����rv�]�f�R�Cv�]>�J�`hC�5H ��%��iD��\��X'f{L�c,�Yi@}�@��O%��Ut.F�a\yTd�v���dM`"T�R^i�=%E�� M�a������5/vl�����0ᴨӐ	��9��B��d\q��U4E�>̫.��H�h�B�? 	�މ��m�\=W~e�u1��e���o�`�U��E�oB��M����X������_��gȷt�b`�_�r����vB��!��˂�<��T|�+ס���`�I.ag���Loy!x�?'�����H/�%���mg��0q6�1ADx�z�ڑ�ᖏ� rE�e�j%v��Z��}�mͨ�YJ=`w�LG���M�BtH���mmD��}c��L��ENR�$c���E���0P��z~�7CEx^	C��H��({SIX[G��`�ObL����Ϣ� m�0������mͲ�KF�R�qc��Jt����͏�F%d����UU\엚�>:����|ܞ��@W�$7�K����a��y�	�����$L�;ذ��D=U�4�Cɮ�;�'K�\�`�.}C���������G��FBK%��盕 >��@�:B"���ҕ5��(�LPg���m�?U��Ļ��4�Ư��+�u:�ݛ7Gh��{'V���U�)e�
�\'� ��6B�u!�����tܥUz�qy�D\�������r���jWz�0J��]�)V_�z �c���q�Hp� zYo��o�n��:`�.S P�S%�:y����b���e�;�|�m?<��ϕ��|���L���E�FhfHZ�����`q Z��I���P���;�Q%<��1�W5��4*e����~��Uj�E==S�~F����`���s!��$�v��,w#
mښ��ۧ
+��pQAZ ���VM��F��mő㞚�d����qx���۵�ݲ����L*+�/��9$}�B�k��U��~K*��o������Ъ)�#j#H2<��z�T��0j������sk}p�Loe	��&��ߨ�I��ۿ��"C�L8�B�n���¸-���r�+^��P�@�I���Uw@#
�Ŝ� �:p�d9l.��m��U����Lm���=�?m$x�
�Sl����Z�)�x�w"�8�b�\�+߸��W�C`���^�D�pB��y�|���Qr��기(zK
�_�����@��%^^w��_`��s��	B��2!�4(x�ܙUic�;��	��)�m�r�h��`tu�m�NX9\�ʨ ����dM��`����y��+�f�9��<���R���z�@՗��!��b�Z��B�`����G�;�&����`<�e��D�Ł+��}&�]��]=ȢY8/�_�6@}ݽ�.����p�_�P�=�R*�)u���er�[���U|���|.}{�I���r���AbS��e�(�Ū�iyu���T�Z��	
�RD��\� ��&�6�u�	��,-�(�=Qv�5�!"u�R�Rt�ck���FGo�� ��T:IoVpZ�k�ZBNQ�u� ��Y�ٷ�if��U�B� �?�s�_�揦k9��$s������gc����Ge=�����^b4$��ч�~S�<<BUU��ߐ6�%l<����=*;a=,��q#��z*,�&>�L*x�kzsI#�������W��P;2�$��je�+��E����_M�FՌ��j$4������p0L���,E�ɐ��F��){�Cǧ(��axۤ����Ǫv�Eg���ݙ�ݹ��h:䩶�}#w?�_�)���Ϧ�$���G�����i6��8ޥ2A['+�k��y��X�����:`�;�MI^��M:y�"��拷�����M����܁�lr�2Ko�1��]h�^]���dDQ�����E{�*�g��	4�鰴-��+�L�x$H�����*�(k�3X�� �����
����0����2|n�����-U�ﺧ�t�]=��fü��l�.+^e��m��f�����V�B43����/�o�^�<���,̒�Wُ$��{a��r}�:\�q�e��+g~�ݑ�ץ�G��.�8@�@������
}�����#>�#e�+\�{�=x��D�OFMy,����	�M�}�#��s�p�/d+����b$R:9�7�|t%�g	VS�	�#�p4�?�8�X֪�Zf�b��"}D�
�� G{�T�)(V��	S办�7C���M�g
�Sz��ŷJrY߻�IU�����R{��Z�ڿ����M�k��?�ڈ��$�6x~o�}��	.��"jiޢuvI:�[�'�w��-9�VL��	bP0��攚#��5P�Ohco%���~��}�B�~6��]4�a4.�)}���f=*&�q�=^�؋G˜;��3tӃ���� 3�,>$Q�'~ �G0,"��:l+נ��t����Z[5�)j8~d�6����<!HI�݋�xb޵���c����	���)bt���d�4v~�Zda aq��mװp�(�����XK��_R�TkA7���-����e�1No	́W����L�=��~Ok8Z�7�3p�\��ۛ䛫�K��o�)У�R@� ����3�S 7'��s�k|Q�]��h��,O�,�]��~�c*l�� ��Gѣ��i��t� <@�6���cIja�E2P66Ψ�_�LDRK�t}�@���� �hg�h�����"��S@e�/��Z a�o��À�e�9c�k�< >����4Ӷ���j]R����H���2����#���Qm%Tq�I��{iG�Mt�P���֊��L��RX~���o�9%�o*����&YuQ���vE�@ϩ�A8.
���0r!_�4��R45��p���(聵D����Q�Y�2q!g�:c�h1�ue����<b:�d�J�4���r�_�g
�w�	W����c�D
�{�'6����/��)DX�!�1��KT�v�~s�ԫ�߽qݜ���B���A�i<�f���em�2Qߢ��"�������'����l�O�U�d/溨��2�b	M��iYw�4�9-s*L�n���ѫ�����n�ps��WΓ��<����%��B
�]��)[�YX70�(	+t�=�SF�$����h�l!`�5�y
%�3'u��&��:��t��`ab�����{ԃ�����$�0���!"�$2����*�Fd؆f�g=�Gh�d����5C�
Q��褴������󿳡��`��*�l�[+>�+����J
oS0�2#���[�6�*�wX%&
��k�Mf`p't�G�m���t$��X�FA��..�P��ȝM�O�r^8d.�7A ���}�#.Z|!�-_-�=r،�e���]'�W��������_+�d�Sc*hID	���L�@�}�����b�^3���A�pAz�p��i�j��V)�����\���o�Y��8�"��쮐�تl_yY s� �Ϙ�LA�C>�ʝ��0]���==	���j6't�k#m�����6��#qu^��e��\�z�Gg�"/o�<@�#j*c(�r��Gͫh����T"�sZ��腯�6�-�=��7���y���/�kգ`��V�~�6��qh2X�s�*�#��	�:;fI m!�y}D[t���L@q1�Mag��PN��I���_w7ސ������2��\a!Zo�oO��盠Ev-�J�,�;��YA�(h�4�̫vg��Q�9��WRp�t���pJy<S;��"	��y�����Ď{H�8O$L����~Oǔ��Z��U|
�Og6G�S�Xb�P�9��ɘ-m�{�~�H5�V��I��Ww܅R�z�@�������T�I��S�NCah��M����A�3��0a���s�+����NUP���n��9zx�V�\��,���M�	AclAs�j9ali\����.!�جI;H��%v��U��>��쟑oe~��%�L��>��x�-�.�x�
�������L&�#�)]���z�^��OT���։v1k��Oqq]�vXT�*��"����C��;O���~��d�8�XjA�I���=6��)Ka�a���1G��TߣC�xn�!w�ݮ��/-+�K�u'ȧ�u�+��+b�11vu����{k�6Ӛ�#4\t���}���3���ʉ97'z�Xˠ!�{�~�+�	g���*�T��f����� ���Pxi����{�a�
ڙ$qY�!8���v�[�S�&w�>d[�ۗęI���C�G�����A��h(�ەncx�����ڝ�buv���Aa�u��c��F휛���K�Đ��tN�����'?3l��ׇ��FhG.�˻��m��ְ)��W����+�-OЄ�a�V�9���Еh�`c|�1;h����T���v)xS'�:�h�_F`�I)8��O~�)HL����#�m��c��������[���!H�:@���(���=���ea��\<��Nz0�����~�b,��M.�����G�/oiqe$�%����(1�eǛu0���󆧐�;�f������M'���n��u�PE(���c�Ӧ�%�:}�i����9)0C%˪0%�z}DLz�M�=Q͖h¸��i~�`D�i��pgy&Z����S�:jf��<l��*ִ$�[��u������3*�h'︣��<O�+�{e!m&�~*I�[DA�mHj����d�Ã*<��4�~�I ܩ�M��يO���s��gT�B"�" �,��\�T�Ɠ��*��`���-���:~ 4�*�.G��T�D:�Y�V�;n�Of���m�B�PK���d�&�����/A^�ƈ��"r�Ѣ*�Q5�ݬ�,�=xW�<.�y-�έ3:ñș�uIRޯ�Q�5���B�������b0>��߁��u"O�f�Ã�P�ӿ�%�����m��9���j�^Rщ"�-++�7��O��s2],������2؄_�\g�������(>~�+*�q@pq�2)��^��n�S{�y$�Y�V�­i��;T5�윾Tbz�[a�[�=�f*ǪQ�/�'�|��(��$�{�{b1Qυ���: ���"��"�8��a5@�B� A���]�/��=�/f�������Uk˯�����e��jȸV�&� *��S�����ш���={���EC{V�u?������ֿ�5���3��+��h��^�85_*��p�{��HQ�q����I�t����H#�����p)�j01I��ႍE���$GP���&@q��,��'���c������O]�������L5���hl`���� �P�&��&
Bʵ�����H����:Nf��lç��5e��V�8�R�O+�Un����nu�2x��Qs\�gt5��y��Q`�5$��B�T>�v_�R/P�% ���u[iҧ�M���fQ��ZFXN��(��K[%{�Q�^�<_:��79�����: ���>+]V�y�~IOv��{��g���׼��c�heZXn�)�LM�fCz!�O�ɈϹ���\xp�rå�왘o@_�CD�U�.�<�V~�:Ľn���3&S>����}
� ��V��̵�(JtA�f %�8���Uj�2/�����,������ ��a�=w�����{�?���?��+A��Q�`ߎ�\)�C�89� ��r���S��Z(�ɤ����|i���Pɱ�����>D��V�3�k���m�+/�V�@��+y�T$����cF�x��eqߎ����"�'X/��� y��	�g� w����Bn^�d��}��=��s�2Q鰶�
Y{�ΠHӦ�~��^�pp��g�kTu9�H���TdzK�.�?S�Sd�����L�;�v#�C�Cx��@@�7�R��R�L!D��P��B)�;IE�>��������e�Ҫ�&�P���[;�)[�V�_�����fW���&d"��u�F�`�q��&AV�]���R�h��=&�(� sK�^�F9%d�?5�
dy��&���C�Ɣ1�.x�υ�?K�$\������z���4�h��*
���}D �H��G6�yN�Ѽ6O�
��Dy�fR���!�:�cꎮ&����ձ0��zB�s	�9��%T�p�E�>zLo���`��joV~$��B.v����Wڀt����}9E����*%2�9~�g��g���1�Sj���!�ѫ��!b�E�P�H5s����0�`r�b�	Kha��b����8l��ֱL���n)�ܸ*��Y��B	�ゎ]^KkK���q�P���f�bA��U2���˥�o�l��xZ8m��q�U0 kH�u�lg�2<�Τ���GE-��Q�N��<�w�{�+<y��n���u:&I�*��@�q=�?����"#d��������Bt%�����fOLRF�#�#7&f�2�jGk�zJS鳡pcu��1U�L������;��v_<�A���
ZN�u����/�f�o�
RV�s���$�C�W���`��qX�ſ��pK�w3Mn���qGi���Wϕ2��TO�C�;�����3�Uj�a���u�H�Gz���3��
=y�Ϳ;>"&g�4�dG/�+�����$y��ΙC�f��J��\�{�@�ϡ��Q��s�2W����^,M3u�2��0�$"����i?���Y��c�!���T��@4���KB��vIX,�^����J���N	@2�K��E7�_��?��ƛEK(��A�<u^$Q��3C0��N�KG���?���V��C)�N�+j꽃wp�a:"fж�t\�ER���
�C�̕�	b�w�4"0N|D.4�Jx�k79��~IFA�;8�����𠎚�������3:��Mq�BB�M$���A��1�ߴS��hbĳa�3�]�?�cx�I������ &������N�E	Z���<Ü5���of.��`��l�?o�3��CC3q�ɹw[g{0��\_�D��'�5i4.�➅�f���8�90�̊��
r[?��S;x�>%�9��v�Ҵ�u0���L����" R&!��g�W��]�	s4����X�� ��r-��<SX�1<��e!�H���{�9��`��(u�sb�b�ن3�Ƶ�Zʹ�ܒ�!�4!�F3�y[W��k��<L�]�̊f����+ju�7Y�kwA���
NF��3 FV��H�Ȕ9�M��h��?.�h���e;�h��I��K:����2��q8qx2˦Tpx��{DT�
8�to�}Ч��U��{��܀C~�F��A���aO�,	iq
�e�X,��o��Z�6���T��ȉ�9�K2܀�0Ѓl~��K�zF(�>�lR|-ha��Vv��o�������Bu2�奅��LW>����^�������uh�U�=�0��<����rF�o�W��e_J]�u8~�aY�UDjHk��A��	���^1 �]w�ats����`�(�G.�
��Y�ՊJ��x<���*��7��ww_��x/��ް2w��B�����w�9;�J�@/I*vio&B�6���œ^<�����s޴�3�� �1��7YGo����9�t�Ay!{QȻ?x��#�����̳�r��g"��j,? q�ďo��T��R�~�+�-���PM���TG����F��pSP4o�+�W��ew�hd�;m/�?@ف�����4,�c`�d0���c�/��$e�u�����3,�׏����@�t8n�*�k!Cr��y�ܰanUn!�7>�~���O���2�h5EkV�APRp�oiu�l���p��XV��=8V�KJ�-9AKy���/ml'k�A`B _��W��}!�M�%�[3�ī�����&�Y��qU\�X�¼�$/�GUaZ�&{���ң�Ll�����=��`��6��Ρ�O�`|Y��]}�V�p��Vū尸n��g�A|Z��*�`�8A�m*���� ����F�QM�{{��(��U�&�Wtb�5��{鉻�������$�%R�����ɜ<�˙j��،,Bu�ވ��Qc�WM$�&	���Q�Φ ��4]�rփ�ȥ(~;%�=���l�fr/|���h+0Ȇ����"P�3�G2ێ�����֚��c�<`4��8$�o繼H �� �n�B�?��S��}�W��+(��=<��(5����fA�Qq��H��+���$k�f���X`K��/������U�7���W�Fq�Ǎ�:����̥�#kf�:kE�J��M��e��R��#�+�J�<%���j�\��%�i*����]��P��5:�1܌��Lֹ��e�T:�{�t�0ʐ�˼�nQV�y5x�H�'<�Lg;�(ɨm�����:���EJa�<��R���W��qy!ɢ�C��<�2EgG�b�,b`�pY�o�i�?��ї�,�Oo���b	���a	���`�BZ'�K�c���hyh�.��到��)9��cL��������Oձ>���O�u����M|:Z�л��;T;���u�B��C����Ȏ]�E%<�Ec��	�3MJ��
; ����7�~#v���e��#Mz�"��	;��Y�]�����	 ���$UUB����j��?H8�S�`qEYr�����c��s�u��_"tr��y��`GZ�P
Q�4\�f�Z��sy�}��co�q�#+5[�י�����-~����wifI�G�d�q�
�bD�1�?	�d8̆�֋�����TjXh��@�X^	���f�3W�]�T��4lZ��;W����)�'iǭ��Z-���u�!^�7���t�-��}�'�X��q�N��J1�K~���Y-<��� u�+Dl��I<��/���?�ɾp���R\=�8��15pw5�$/q���Q�C��� \֖J�V.��c|73G¢�aO���^��`h��;-�e�H>*��Y��]Q����Ĺ��z�KR���z$�Oq|�:&Z� �k��#`����Nu�}:�EVE!��c�N�����n�s��C��}Yc ��q�A��̙��C�L��~�AC
�&ޥ�4)Ϙf���e�YP��N0Uu�Y�� Tw8��\���2�Sg��,��>��,z��E���1u�V&�c�g-��'KgR|y{�!x�!MC���Ǳ���f�ĵ7Ȁ��b�]�o��F'��#��b�iUY"���t�]BL��A]?f� �ֳ'�p�����c*r�!�Tc���a�a,����lK�4��(����ѽ��׻��%QB�B�Y�7*R�v�tD�I����C�l��Yl۩�p|�Ǽ�J�4N�#?��X�@qb���5�2�B��uw��o)u��:��ׅN�M�]ثHa�sOwC�<<L
t��
R�3������������e$̴�� �ƏIq�3��
g��^�YG��Ɍ�Q֗L����)7D�1(�ְudb;Y6����k�hԿex����k��$�&97�`��UI�����`�ܛ��5�Fuo���֪��Z�q��x	�GS�J�O��
īP�3��-�YU��b���,S�̈́�y�w+#�����$�L;t�]�4�RB���,��s�ėI*�Z�m2�'��1�l�!2� �"ȣz�|�0Q���F�ϰ 9�a�5��z�Ĕ�,4
������A�a�1�(A��R��r�;A��<� �����A������q� ǈ`��c-pf�
�k�,bqU�����o�y��W�s�*[�L(M^�k�vZ��\��HhQM�XY�d_�d�j�	K�)rG�F�����U��N/���j�"�j��˙,�Ͳv���#��^	NB�����#�G�z�v�ߏ�����rԑ��OrR�U2�xx����z�3WK[o�h�_�k�u]Jv��X���PD\�dO��<�{���翿����í�an�x�u�{�r�&c�R�x�\��:"*s6�����П-E6q���U0;5�u>�"vU��*��E�̛�('`��5��2�z���L�~x�������"�~^��{��ya9��J��uC\���2�� C�◪I")� ű�	n�$L�F�R�d�̎���n�a�@/��U�h�*/�Ȕ����� �\7>�0`Ԣ�Q0�Y�����1~kRb�H��5���s�}� 	[Ч��Wv@�Ѡ�6�;�0���C|,�O�T��CjB�gw���V(������K&CٖE�:�)FW!1��S����y�,��Q�7wS�@�=����h�{tQe�$Ŀ|ZG�:���F4/��"��;�j*�ഓA!�w��@d�Dd��y)W�(#�Á��':��kk�>`ej���
��{1�ل���<��G�k��i�̸`: =p�}��@��$kJ�h��1�y�~z:p������tM��~�h��P�?+w��_+�j��Ϊ�e����h�k~��	���_�V��m'p:j׿�b�rJ�)������\��g�UeI54�ԷE�~k�Qự
Q�,�z�P'�	�w����G>!M]J�%p��Ά(���>������D�H}�x�9D����0dM�ɠ�9i*�Q�	�t���JCp�5�V�54���r��`@��-E���KRc�>h�}�o���sǵ��U�~#\�5��V��Y�,�v��?�];���ȶ$[����&u)���^�6K2�b%�q~/�Q,�oT������>��3q��%!�٧�qo�\�8)� =k��o�^n�t�j�D��/;��|
�v �ִ��/s�|*M��O�̼RƢ��9TA1&C�\�'�M���?��i�?�n����l�$.�=O�Ӧ�ѫ�$����g���E�i\��yz:������&D`�����Ug���FS�Xb�26��rM1��J� �m���4���1N�E��L���L�@r{n	a������Vm1iy���7st�:%�3�B��z�G����n�G;ݬC���"A�5��Jex�Dp��<�]RQ��Yu�@���	�I���ܽd�% 
�Pг9�j��V��I�1�G|t2��K��d\A����8��t�wT�i(�fC��4*�q����
?Z8'�mOI���)P묔p�cf�e�	9s�w�V#��N(�	�0�m�����` �b�����?��LLj�q&�ٻv����Or}�p\U����a�
H|0O��c���ܸp6h�C����h8G��F���� ��~�ߴh(h�q�-m�D���=�i_¾/Pp�F��9d�rW�����v��Fg����t�+
c �[�����?�����a���	�̫���Ʉ�ћ��gΰe�6~����?]������jSx]H3�����@w��C-��>}���a+��bZ�k�轶����n
��4�!���,�_|��DKTn�/�*8�=���:"L���`]|�6O��45���F G*Z��Q��j�&�%�`�S�!Av~\l��v���is��bI��<���UP��i*���,����g�q
o_~�����Bɞ�Κ�RG�n�~��wN���m�u�6��AҞf��͘��H�����J���<X
��=.����5�1�m�Š\ɧ�炲73ߓ)Ǒ	�����|�/.붠�Г�?@��@}��pD>	a>����w���L,�6R�O�S"P��ዒrRFf(<�:\Yoa9�li>B�L�y3t�9r)A�8��v�r�<����N�1���c&4�
�Eb9[/g��Æ1�"���M��C�`��+#��(�7K�^�z��:�)��������1hIUj���˺�Ӹ,��Uo���t��:�iz3䋸T�gJ��!uE��m��/�����Y�֔%
[]=�i�����KC�� qU����� �/����O�ɱ�׍W�!��r�jnF..��UrڗJ R� f�1YSPpU�LG���BgM��Z�F*�X�ֹ�{���px���h���OB]P��b��N�N
$��O�m��x�lք�eǗ��5^�D�E�O��_�(]���"Ϙ��T�L?Ɗ���mOG.��T��ul��Ps�4U�[y1ĝ>��[bZ��L})m!�C���鉁t�b�p*�V�J&��4��֯ ���[�O͑�w6^ ��%m'b�>t��X(���\@w�`}� �m���k员[��?L1���7�n1]����I��%!�q������m��\�5�������S��W�8�P)(Ȳ!�y+�y�k���i�u8����j��)��ך������
���m�����D1�OD���5tj��84~��fcu��1���wNU,�3�_��	�?A��5k�="�� ����=@]�хDQ(e6vf�U�U������A�f p�0sl���J���Y�+��k	�����M���d$�wt�R��Y��K���m�_}>���w��dM��.�ݾ���9\Wb�������_�<��!�?W/�̓�)��Oț�F}~�O�+~��i����k�� �XG�0�B�6���������rl���3�lH�oȓx%�U�(���g�
�s�q݉y$'��7�̍�=a���1�8c0�Qy��uS�����<�ޤ#-�r�ϊ}�{=ba7���?'1Z���4�7�Q�˅�'H3�,f���Mx��'���
7�{���6h��(͌{��ݻf*I�(��e
-��H�����lz0��}B}�:��A走wCS��ɉ�$:�����	���I��;l$؋��
�\�έ��f����v�6�2:_'}f���5�tX���Iޜ2�G�=IH�\��|[��d�xD��m����Q��2,��v����P\.q52��(}�*q�n���n4_i��}1	 ��k-���������{�f1Z�h�Z����D����r��;�J��������K����<�~�d���)���.��q^䤛��̐�ǖ�O@^����������~�qbe䀹�,�8�`��Ə�#����/?6r�G��ت��#� u����;�˙���ZX��������vyuŋXrf��qY��t��� �Y��F#�uZ�؍煂Y��X�`۴ ���Dh���!R�}fxU����oO���14�-E�0�e�}꥽f�m�l��Bצ��~�Y�jo�=F��d�mV�v��͌Ag���r�<��Nr*;K��Qp�����(���}`B���F4�r�1t�/(v��%X7���5J�i]x�a�x	l�o��� ��`����k�q�uF��L;�n�����ZU��oGZ^�t�U�@��^g�Z�����,`U�h�\F�,g9������;�k�!$��l=-<+vT�Q8�������S]<�L1��oE�"��邫�B��u��6}�%T���=�:G}���P��L��rf���Nњ|����hl��C������K߲��_>ʍ��
V�� ^fBґ��j���֘�W~R����#�M��/���lI��Hw��Z�}S~��h��Z�0�,����}ᩯ�r�!��I��C��'M0��hN�{:/�#ݶ/mycF���B'��	=
۩�LcT�ܚ-͊�+u%?-}O��5��\c�(�P�Z����|�Pi���ι;v���\b��	C`�gyR��#� zqUZ.2g�֛a�N����t�e���DƢ���D`��#v��=ބ�8�����x�i?�;M!�8� װ���������|��hfx k��e�:3�L�u|t�� l߯˺^���=��!��y�o��yf���իyLč8ɕ�dK�g��_e)g;�����)=���G��ȭ�c�LfG'�z$�n1t�������J�N9�O?i��;+adyw2��cGԂW��?7�/o�E���V������.(A$1���M�� ai~*z9k��V\Z��Yd}Pv5_�Q���7ɓj��I���d�D�2�Y��ތ���"h�v�x������[_�R �2Q�P$�l꫓$�z��7��́7�j�ϥ��U ���L�=���<�D �}b�+�N'�����[Lk=8���E.�l�*�v*-���}�d]k'T�E%�>�U�6�#�j�1��/q��uE�;�/dG4�͌��ܙg�t]CO�0"��&��+���M:������( �""e\�AG��I��g�䬋w�lpԇ��*	x5md��c�fHfx�]����r'��E�P�g�"߼��N"0�����?���q���*�D%'	�By`�nH���~�Frmp/�.U�m��<1��`�r-s�.oJ�:v�]/V��i��:�K����2e�d����[ڽ�Sy>��a(��(R��D|d���<
s��F�M�].D�&`\���!��-���n�l��;�@�u7�t�z��ƌJ��K{�`ܗ���6�kl��ZvMk�K=��Y��N\	0���A|g�q�:8וv�-�G4���^U��R��4�HI�w���u�)����i�O�
��������C	̐ D;�M��ejQy�b���;����v�Yu���� �|s�|��#%�dN�/q�ݓU[5zU��b�.TO)����{���)�cӛ��t�0p��ZC�@~wDP9e�KQ��#��l����T�0 �+��b���m�IJ��FD��D�d�nm�l�l	��/����+��&�E-�t����5!�(u�X�3,U���c@���cN+��R��-`�=1N�Q�;�_��ITT��=P�Fx ʈ9+ ��%�z�t��U3_q�9C<$�1�[����'Y�����1�ȂjJn9Q��ˉV:�j��F�1��R)c����JjSx�iR�Cb�:xo��!#�sK�>cQT��K����'�4c��O��d���_�&��7L��Y�`D�:Dӭ��c����H*=m��� �J�s+H���%���`���F��	�5c:>v�� _=SM�m�;�S������ �[�e����n�=9�)x����)�؋x�N���;�˩l^�J�Y�:���i�7��%�>(�ѭ���]
�P�K�Xx�M����4t�Øxڜw�,=*ۮW�1�����lf�i�V:�n)�	?����a�+D�;ë��$`xz�/�sR˄�눊�AuZx���r�s�zhN�S>�^wƁ�U��}�Be��N:�i��?�7���]v�C�o���ߟ�`��uYԱ�T�qzx���/��`XK�m�p���UJ�$�>��8�=?��4���%�{����<[Ь.�]�N{:�
3|��!Z�Z�I��]"t��ԓ�ڨ�a����+�~��'��z>��j&w?��`�?�"��?֭�7�ڷfN"W���\s[1�O{��"%
F�v��ʞ�ܤZ�\E���Վ�
h8�̄�磭�J��0�_�	�xM�0;��M0��哩�!�����]�U���	���A�'�x��I-v�#�&���R��CZ{!DK`;5,>��ћ�S�-%�?���j!�">,�f�<`YEHq�(@)��Gbg��5��3j���`d�5o%6�� �J,���]��+�a�H����&ֆ��лɏrij�y����*�q�"�
3���[���F"��J�|ɓ��m��f��AKu8�v�.�k5���#��w{�ʋ;(���F������T�*p��۩w��y��[��� C�с�?�7�����w��}���~��n�f	�әj�.��''t=]�,��'��9l4D�Y�~g[.'��b�Y�����c�~���J\$U;3����],I&��,ۤ7������C\���;���!sW$'���]�KZ��Z��!,��ܳ-G�+p�5B]��]-��ٚ.J�A=�
`�ĕn�n��D=��-��I,d�/���j��b�"c�1Pf�u1 �:A#�.+^񼰓��_�%������!�g������97��VQ���;)��tϦ���-ō=�k_�l�t?(А���"�[V!x�>�� �ɩ?=�3w)�������2�Y36��z-z�[GE^���NLfG�r����`�?�@@�a��=5���J��ޓ�8)W5�TJ�����W)?���y�;`�Ns� ���=���S�L�i8�*d��LB|�PU_�E;[M�t�����?x��E�@T���Y�/��CXQ�7jQ��M5oO�a��=��d� [���`���ta #1��7�[����}��FY��1s�De�~\ZJ�Y��%b2��'�kC�y�"H�W����v���x�j�W7#�Tz�/A	�m�'�z�.tNąϼ2L&�4���eQ�F��Y��5 �>��^3��;�4z�w��˴2��K���]�n�D�x�(F��d���b��f`ē��*Q�� s<�F\���|g���&�3f��EY�"��D�8����;�]RI�8��k���	B+L�V̾��!�jz�Kj|��ޠ<��0��A{�Yo��uNAޚ�i�n��������m�����K}+�Ci'şZ��[��c�I�ؖ/�qx;�O���Rݧ7銮i�����lk��n_�Ө��8N}�"�ג������М�u=`��Fe�*#K'������'���IcP�NϢ�Rg$��L}F-e��!�O��s�����JY���di�I��բ����Du.�.�qe�J�r�="��e`
�t�D�rWJxF�
uo�31]�>���n���8N�Oȍ�����J��.;�E�vfj&�
+?��wW8Lx���wo@s��?%���	�B�ʈGً�����TN��=�_v��/�I�ڈ@�nI����x�v{�4c&����*��VCBt�8�kP;���`1�'��Q �`K�xL�@�¹�]��\�R\�����4�f��L�v"'J]$�S&� �$��
������(�Y꼽�f>e�똽�䳙O�.(�t=�(�U������t9�
��,:����i��_I�ap�fp�O!���mc�fǳ�\\���6Xm�It��o���dEq�cL�o�'�wϕx���u-��pDh#n��צq��|i�)�89�vs�r�y�4����7�`��$�n�ĠL���V���m1��D=�qZ�3<�dH�z�!�M�I�]ǜWο�����$��U�/K��!�[�Nn�(	֭�:G�Ͽ���$�:;�$��W���TL�E�_7�۱�K�'&l�v�p�� U��0�����2����#��s)w4�;OU`��qs�-�٧B�YA���Z��Q�(����:9pL�'�gi߸��t�P�'M��̴H�J�DD=1M0�uBkO�P.NO�S��Bi��AJ=ʤ�}N�H3&��;b�XH.��,��A�h' 1Z?��9J�A"��XV8:8 �X�o��z��ǳ�o�Q��	�!H����76�����y<��`�� cd@�7�X56���E̵ r�����S�����W��D��f��s��c�����Ş|��T���\c�Z�XrP� l͖k�C�n}�����[�p�M�(*^��\O?�d�m����G��Ūa l=��ʽ��f��J!�BGAB�({�~`rv�Eʙ��~���~����fjRf/�95I�9�
q�]7������Դo�a�{elc3�����0���z�*Lb���}�v^����� W�P���L�z"��k�,��|�ye�|  �@y\�Ӽ����4i�}�d**��� �X��I3s��@�F�N1@!f����'�V���9В|�+�R��p��i����@A�5�p�A�����������������o�f�3`=�l��\h
���/W�u�b�6���\qvD	�l� \'RAǬ�P*W��'����g��܀��}����p����3���W����x:_t��{N�8>���Xn�]�ˮ�6�)��)p})sz�~6'�p,
qe�!��3�q�%+�	t�f�g��xC̸%���i@g�J' ������#��"��Jgh缿�tdƥ�n� ň�\S\�M�I02��|�Կ�};r˙��x��w�	�Z�Y��'��*{�ȝX&%����U�;n���u���'��z �f>e�*�=�_[K^}�S�G	���T#�
\�,��X�Y�*�i��*��,Dk\x�33�6a�_������n��r-�R�3�̨ss�ܩ
'EF��O���R>B�t�\�gU�ѡkȻ;�]�F��Q6Rk46h:wo�cTU�fD�j������v�C��z��zL
���>�y��xݰ�L��  ��('����εj��#H�M�j��U��:�[��ܴQ��`�Rמ�(��7�3�zBYa�z>��
:-c��U'�Hȓ�}}��C�+<)����j��K�t�һ|5��=ǭ7)���K�Va�s
P��zГFd��J�ߎ����B�{J�[s����tJ&x�e߷]r����F���x�̃���C-����C��<E��󩅒�=?��<S 'Z��ኖ�E���γ\�E鼏k��������]��	�kY�G.�8�R��FJ�z0���nf���DP97�c�3>�q��SF�F�6�$18|4����}�X�f�0,���>��p����O����I��x�	(ky���4톴W�F�Uj��&SV���f0���b�CN�����Aq���l�qo�l��'Z�ř�8�I�BĎP%��'�k�'����W8���Ӟ��e|�/>L�/������߷��-�H�l��1�5��o(�S4��6h��a:�
��P���'���.]�"��s�C��^�B��{��=�BAI��ݿ�4��0���/��cb3w�G-&CV��k�Œ�q�(��+�%���8
3��W���1�w������G�o�x��w���>Coԉs�U��.���S��Uv  ״h�ta�[�Q7I����RZ�lh�U'���+��n��0,_����Jm��������J�wH����4����Mu��Se���-�=CZ��9r2Bv��Ӓ}Z<����φ\
�WI>�Wf��|y���(�q��m�-o���t�v��f�m�R$a�k��6(�0���:ͬ�2�����f�66��D�j
�i+���H>���3;e�Z�r̃l,�%�4���'�7>�`Ҕ���Q��·��bo>q\*���2i.���J��B�,poT.4��}���H|v��ބ������{��&
7*�>��l0��y�����|�ܶ��1���C�ǀ�KVI��&㎦��v �G�/Il�S;I�))O0��h�XƉ%3�$��^#���\R 5��ֱl��47@��y����R��K��s&�1*�=K���%�,Ι��D쬁F�Ҷ�z�6�k1��D�S���BG��r��S��#���~�K�"�W��b�+Ļի�"���})� �c��)�>k�sGRa|����Y��K�9�:�����>��m��v_�X�7ߕ_�,T(��F۩�f2 4��>�4@��4C�	�������D0 _6�s���+�\�^���0�<O�w���נ�^�>��Ÿ]����ho���'������Mc�:����S�o�c��*�p���5��qC�%�.��RE#	O���!�*���ŭ7c��R�s���k��Y��	.vŞ��OzeX�5<4޽1�C'͐��E{Q >����{��]���ƻ��9��"u������3hD�Q��a�)M��S۰K9W>�ԍ��~��4PPi4zzE�(P0��������a7B�2ܪ6�&V�G�p�y�tp����t�h�}���a��5��4��P�9.���8��TS�L}d��[ �$Ν����Ї��c��j��3Gw��͜
 X�%y�̲�.�rPYuS�����D�A�� �#Ι/�;#�]Iu�2bZG�{��M��@�Α|��9�
�R��B���GD�=^��yOX���zH��B�/��x�9'=)���Y��W���U���b�;�����08!�R2/���(p�[��Q�H��/��PE������K"�Js_j.����<����|��u��Z�[<7'Y��y4��"�T�O��:ZCU��<�Ƽ����4�s�P�� ���E�n"_�xԭ�F��7��r�P���,��ǟ�@��^!'X�����}v�,>V����<��I&����4���C�2Qޟ����G+�0�����nz$�u X��M=޵-=t"VT��(e����*��"k1�.���b}k���C�fi�ډ�MH��asµ�qwԴ�g	�7�@[c������k8�^�@�	j�s�Ar�����fI �6�t5��y�7Im�I����H��I'��-
M9��sNk�1�
�d6�Uo����㉉A��e������t�{��Ι�[8��Tp�֘`Xhz�ՎE�sj96��Fe�fZ��g2�A� ��wã�0���[��W�fl�r��sC�{�D�!���	�L��%<�(�]���oR���a}K���5ʡ�(Cϼ�.b�&z�I�����?m-o��g���X�+w,���K���zxn[��æO�їޥ�,�uNy,&b���$���dy�����9D<,����ZR�+�2���W�f2}���w�D��(O�����~� �|��y��]��ctqf�dTR	'���`��G0R�T.%�S�{a�������K!�!~t�� �C���z��]���O�����j��V��F:�e��"u��T:����g�W�]�5`m;=E:���X4��Q�+�^�Z��Tn���?~���x�I���P����6����'��2�6ӎ�Yz��͸�l�e�=)�����}$���t�5�G�f�Ʀk�ˈ��(��;�H@��9��$��v��}��k���+@uS�df�&��b_v�{C���P��y)ߪ�6>��FFiI�)�־�:V�P.������:9��Ra��7GW�#��j>ϤjV�nh#dI�I�3�4���wrz�$��<�>��� ��t(ۊ_�P��R�b/���ɑ4�����5ӊ/^<�WZ�c��b����W�!��v\jl�d%O#5�91f��ve;=V�#W=�lFG��"vQ�1,���6���<N��Nq��ln����*���9�`��߽��?��G<K�ʝ$����UK������ai��K�)��͊�렰�yb�Pv�^(ꆼ�b���<�2+#x��5]��Ĩj�`��w���m��G� ٶ��_i���
%���n�ß]u���"viz����l�8g3��4��kj*oT/[t,O����0Լ���y��B�+~H	�v�����s��`�3qc׀ ��$%�R�k\��T��G�[�q�|{C[{����L��_�"'�e��Nt4x 4��� �G�7��&_-�ϑSpM'Tr8�wq,�n�J`>���}�v���T�;<z\�,��,az�_�'$Ma�K�b��L,�����X3}����~���ع��~�(�2�4�����?S�-�/E-�� �l�pw5�v���_V�µ%�F��[���=Ҷ���;����Qu����e<��n��ɪ��E��Ж:9� }����S��0:�&P�/{ᔲ�ޟj*r){��#�e;).L�a5mX����\�j�I���J`��6�¯�z�>"�m-܀f-%K�YЊ֞�^�ޱ)��b�����K��eʈ�zT�	��5=��[t��5��l ���_V�R���L�3�M@h�1�ɴS6:ښ�C���{��w؁����<��bm�t�mE��G�a8?66�y�3�~u�Y��qW߭W��xU�E���c��^�|�x?Y���+�L֝ �b���:�oҗ�|M�]^?�7t������_���#���d���� 4q �������4�[�Ooo=�N�(i��� ���[;Y�
p��㔊�G�!虦�*]�
�j5��;m�^����z�r;$��]��"m�1�����\J�U@�����F�7�bɚV\�p���tz�Wf�N���d8���x��}*h�����9��ZA�Q�d�gXu��8Y�� �{��i tX���AI޾�l�֡Bd�`SW�E��Gẅ����»J6R��Rn��L'��\�ok���8U�u� )��"]H,8`�KRea�s��Xa~B�:�JY�J��]�3��I�e���Y���қu%l>�oJ������o�2�U5� ��8����սI��n�����}��h��m�6�ǈabK��
?ER��w�i-�8;�F�6��D5����6��-����rP.�gvY�o	'5 n�Fe	��9��d4������JX�a����!�� �6v0��N��7>����Pi	j/١Ū������;V4���>IZK�d��0Z�0)����^�������hmq;i�`e���G3On�/v�0��xj�-?5���$O"�pϙ��7ZK��+�V���zzǏo�3����}��6|D�����W�ODPF˜	/�>�yfU���m,���1�u>��lR�3�If��Zg���Ks�Xt�kn�Y��e�H�����S����V�1����1d���ȿ~2̖��v9ag�i����I�BS���b��h�g�ǫ/'���+���Ɨ~��/"G�ph��X��<����n��6"Gz.�Z����r�;�הY���Z�`��������aZ��iR���kAD~%RIX�X�{U�N*�s6/���5�K<%<���P�������A�/�����<g��@�ʨ.��R_{���+�R ���%���p���Mw����N��n`>`H�NR�"�ζ����/I+�N�~�䈡���������h�Ğ�(��R�;'1���4O�Fv̹-��T�RۯB[����,^le@c�,#�W�㷻N�Va|�ُ���~��u�ZT5��=��w�	zIP#���.D��_x�����z�̛�ce'�/���c,����)�ٽZ$G��kՙ�o�~���C%���g���<�0�j�D�������љ�_S@�MQ�������	�:�=xc�a�'��L�u��mãHX��[Z�Hf����@N�m�.��?�-X+"ڀ��ݧX�Jy�&?}����䃧�킎�����s��^\��,�4NaYOy}ل�mĐ�H���{�-��M�#��d� ��9��Mr�A�.j�d��x�fP���{-4��Tq��9/�$��F^Oz�}e�a����{�4H��N]B:>���u�b�R4�.�V�4�CU�?'UA_ٽ��f!��Y�_�NS�����KY�l-���ݫ(���,���W+c��n�q���>�!	
��2PAJ�q9S,G���{��%k��m�Yv+47��lz��e;�x�'N ���#��(@x������6*�[7Ő��mA04�mNp��"��m�m��;������I�4�?ȵA���C��5\�V�z��z������m�o��,u�G�4hy�s�/(E�cޠ�S�p�T�;?bvJ�e�[vҴ��)6� {l�L[�V�<�������u��4�����b�Sc�h�?}4�~�W�Y��T����78f���b`��\ĕ���-�<�ʚ)3c����Ҝ�oT�M��!F��y�&d�df�zbZ�S[�A<���.�`�+c*@��Ip>�ﴶlp���-�4S���K�N~��`")@y�jQ�(,2Z���p=wX�R��C����D(U��p����o���@8?����b�����A�2�~�JkZ+���z[Wh�B�����R��P).$�{ȝ��ViP��N5(��n�Q�����*}����R��30��������d��6q��5T,|��O��Ic��wV�o���ک
*E])���Hd�E_��Oq��Q��s6�)g9x�g1�;�������{5�	���L�*�����p$;&��	aq��⮫ŉ��6�Y$R�6澦������C�M}���ƽ`̛w�?C9�Z�A!05�5�]������7V������x`,�8n�Y� mS�w�e0���Gzտl���*˰�{��+�E ���Q�P�BXq��6��<J���}Og�q}3��yz56q�U+~y:��1�3�>αGo���sU�n2]��}R�:FA�Z���B+K�-Z8�d�$Eh2:E^���(���]D#iO�;�g�;Ϣ0�8T���n������Ga��"w6��B/֎�?�L�0Ш`��䑙�a�u��ƎI����T�{�^��\��9M����\Un��s�%O1@Q��;!���"८�S�X���k��(6�*I�pYXJ�%��YI\����p ���fJn�P Ƹ�Χ�G��vrwf�:�ehYY��7*������Y�r��8��%�i���!nB�g R����?���O�)� 4/" �z��ӹl@Ǌ�vC;j�E֗��@D|�4ߓ��q�8VPud�{?��F������'nG�0�x�U�n���S�+�
�൪��{qL�&��7<�?ū��n�����E(v&���'�D &c"!Օ{<��SD��G��9	��B��{�6CL��}�[p�n3���Y,7�I��q36;�b�L�s�9`����Th�^�.�Z�fEp������G�x�i�ǻ|c�����1_�P��B�q��1�Np��J���9z�j�X��0%&��<qL��(��eR�X���1^׋��C��/GPD\�*5 ��X�u�!�=��G��՝�T��Z���n_���<t��<��_�]����;V�웨X*p�@�9�]�ն�#Obֹ��P�2X�4�I����b6t>Rb�'?%B��'魜@�����_Ȩ��|l�-�QD�lՖ_g��Y�N�D7'wÈל�K�f��$q�@�,}��)��ڱ@u���zʜy�d!q����A�0���h_����X�����:}�zK`YD`G)��`hl��}AR��P$�+j =�`U���r��[�+a�b+B�El�ټ��Ճ*�6$Ѽ�ĴȈד�f��P3��>a��km��'(�3T��L�a/�<A�w�IǇ�i6�v�C���@2�(!G���wM��A?.{�κŤ��p�	<��*c��`�P-618+��Gl���,zɄp�[��}{��rV5i�� ߂�ԫ"���\���R��
�rQ@sc�aS��W b5���-���=�|g�/�r_ψP���ˬ��%'`̗����Վ���Y�}S����w�g�s<$�b�����7`
���\�'�pgj٢�����7��EH
m����X��/�� O�庚͑Wz>���M�yXj�k�d�� ���L)	�fa�!���3[�ko~��ߡ���{v�;�B��:��L��<y�f��UX�������<$��"��!cHo�RmpB Q*1�+S�׊�1�o�db7M�A�h�q�JB�[gͱa��W������n&U�тxy�4��=�ޢ�{��G�p!r���H ���bY��Wu�C�.�'��/��.�y�5��<�\B������Fn�Z�U2;��vX�	�occC{!�z�-8�T�q��myS>9����P�lX�)�o����|�K)����&��{��L�дI%��	�M8�Y��Ϥ�5M];A�~�x��wY��t�r� >{ޜ2���^��|4H��P��f?��~�V&�h����� c��s�D���k�8,����/ѫ����8+�T�:��X�E����a.=$e����f���Yc�j�f��R���-C�`����IQe�f[8��j�p���Vd$��غS㤎 @��ټ�XJ��E"vu3����bF���zUN�����\��R0h����~�?4�W�~�n2T�(FgQ��R�G���5���o�E��|s�z=]�-�ǎ��A�Ƒ񍻘���[�����ͿM�G�����e��	��Z�S�;�C��l=2IG�c�Mvd#
���y�٤�]&�⹚�*֡u���"$���Kl
���;��;ΤZ^ci���c߁��{�f�գ='�E(��Z�2Zߺ�o�v��x^�`������zΒ�0��w�ݩY�D铕f{���w��$�6Ŭ贁�\-�~�i��Gl犯������n��Ohzo�a}���K�����s�D1d��*�aw\;L�R`�y	q�o�ƹ_���.b�T��M��sk(�O��e<���,ZԎ�����T&u8=�GO\�nGQϺ{�yH]1)�P<g�M�O��q����k �;y����%&y&/�!R�#M
<��T���8��f�y��`��n<��|.k8SKk�oK�(f_:�h�!�i$��&񏐧�u�&2��$8���CT�E7pg�m�bz������q�p��곥�8���sK�)����0��E9��� :Ÿ�Q�Լn�1]D]�u�^�0+�m�?y�I���@�#S:1����B
��-E�Hf��FH�8�ok���X�Jl����8���暳��(f2]/�c�7�,j���B��O�<�Z	cb�;���b�_�[�O�b������i�Nt��::�`�Mh��m���(���j���-g*�|C ]�j(X��qB����/۲����pˤȡ����~p�`ͪ����"\rW���*w�_��n�ӏtE��i��s�e9&H"�x+��S�ěl��O��Ȱ�s�� 	�6
 J��������t��^9m͹���lD�`���R#�Ca�	������3���s#P�
�/�H\��O���-�����R��1g~�uU>��eL�f�@6�,����jW]�@�������{��Ы��kZ��\y"'��eR\u4=h�y�ٶ ֓򜚕#�8{�E��EMF�\�4�e%9��g�ZU�^ꦭU�"؍y�$���p���_.\.:��z��@�@�E`��%_��d���{'���}�x�D���@^��r����Q������Ni�SρJ@}C����d�S�a����,��4�b��n�߁���c��?�a8\�?֐_��*�Le^��6IUU	��a�<�J�b>R(��[F�o/h��>A N0�Q��:�m�z�o����0:^[|7AAp�Mu��LG�D6J�7Y)! ��^(&=D��0)�v���k��O�g�@��9�k�{�~(٫X8W��2i��^����z�L�kO�/}!^��[ �緣=aU��dLM�,
�2��9�M}�U��!����"��X"�z�K��K��?�x�h��(4�z�J��K_�tijz�9Ds��J`l4�p��x�(X�3M����ȵ]�9�0W���"8���&���NE5�����!��D��Ix��<�$M��)o��Bj��#��d�TL���0���gX�s�8��U���Ӑ�`����Z��j���"�<	�jl�`��l.��E̗s����g1oJ�4�%����b$����N���o�`]�{D��x� ��1��B�TIrxƿ���\��e�u�����p�R�Qe�Q;�f��*�i"���" &a#DXe�W��<]j��_&vKL�6	ƍX������}2z��V�?.5����Q�͎�R���v���S�8{HF�{�9Ӕ�s�Ш����ܦ�1v��#�>uţ���2�x݇r��[��z�1�O���.�_���RR�C�hFc)�^c�_z�^�R��y�3
ι]��d��デ��Ђ#�c��
�v���m)2d�v�w��KH�����y��+������AҶE��e궄����cJm�)����j�i��V���O�H ���|T!=2���<E���c������B"��gd�wz9����j����<�����j,�݇�*ǈ�"��}虏ޝjQUK7�}	��-0)��m��2�s)L8ߋ(Y~�5�}|��8�٢�K�?�E4���8&�v#[�E�g�fZ)OV�skG�b~66W-+fs��&��.�����=gD8H�f�o)}x�&�^H<��9u�*G,w;����w�(ڏ��M�Eu;�^ETiFx��=���h��N(K�I, �%t�)��6%ߦ�[�~����ĂΛ������&�!Gޞ?l-j��Q�W�Q0�H'���ؘ�O�Gjܲ�[�oz���Խ�A����f���gH�J�;� �GA�yv��-�U?6r��S:�L{�}���'z����&����x	}�+E��%Mh�B��.�������6�x@�%��y�=�6�<�f;r�tE���O f���]b;X!��*��5��#�_v�,-�x
��1*�U�%N�����v�r�>Iv'	>���OQ��!\X*�s�3�)o{�A�PX_��;v��&�Ի���̛��z���n+����;>:/�c5L�y�V=E`�1Yp|3��V��S	������X��	.4S�����4qs�[�?�ۢ�����C�	��-%3BC8�|������x]�ks���,�\(JS�"� Q��t��簷�LyQ��#\Q�y�@�k���F2s�L.���.��_a�xjk�5]1�fy��y{�ܖa�W��ׅ1IM: ���ֽkG��(�$#	��}[�1y�*�կr�0�,�'�/ޣ���/!A޸$���6���xiq �&F�+�o�%$J~W�9���p��d���_0��Ε)����Q(��^(
G�P��Cp��ޏ�]ay,����76���נ�a���X+��b\ .��	����X�V?���_���-�%e���%�}��:U�����^�������L���E����t3�=gI���8�}��"���t,��23[s%R��;|�����B�r���(ؾO;�����V����u����at�1ѠI2f�CJs/
5���)�,�|\^|wC�݆��(}�PY���"�M��֝�Ҩ���3g�7�D]8�u�d����\q^����5H��>ٓ�mk}"ΡJ���b��mꄗ;މ�]I�F���k��O@_�^7T��eZ.���R[ަE��,,�P\������_��$��n���b�(��O��0���_� �
�8��Q� KK��򍉖�R3�i�}x��Ļ5� �D��!�ߴ�:�/m�k͍G_;D.�y��]��0����Q�a��h�	7I�`?��	4�j�j�C�����G{T�1,�:����<g��@�M��R�/�,�$F�U�#As�)Lc
X�S��ϋ냋��M�s#fD$������Y����'�ޭ뻈�Y,���N�+`��z�v�o�"������d�t�W���ً��pՐ��ӣ�lk�ue�:��O��ɳ�*`)ej��yq�0M{R�:���uLY�\��IH�Y�{���������¦w���X�Ykd'��n��&��e�u5(ji�j�-������]��}d�g��2��h�1�\}޽G�����)�y��N��_�G����J��,K�E�'�&;u��(J�z��PZ_��:}Nr�ĉ����5 ;�-l�Yo�s;F �
Rձ\*�`��wY�;b3��E6���Fn�� i<��燚�w�f	|����j���(�>�ݵ?�f��!O֔�p/G��VW�LS �[��/j?�l��q]/F����ƢH@�B �Λ3����^�W�6RVE�j;A��P|@ @�]�$Z��-�%�J�N8�jM��b%�C�m�V^ߒ������f"�,��Æz��h�H�_^_j#�Lr>��?{�)rX��YwV��e*�xX�M����S����v�p�#�&uX�a*�l��g���
�1��hc+�6�X�U���6�;��,�q
	uV�b��Ӄ�'��2�a���ftk�[[���v�"��ӛ���6�)���W�&��\fo�̆������u7)�yʸṖv���>u=���L�{�CT�W��N��Bz//��(��"�B":{�&P7O�H���b1?��A�-+�)��eL�ݙق��XVx* ��eV`�3k�N�����&�6W��gh>�����$c�~9�8|nt(��Qn�RH�����ۓ:���X�6�| :����jJL��J8Λ�� b�U"�co���.���>��#iʔ@�P�5 ��2�*�M��磊�ar��œ��62\�{��1qV���}aڛ�ө�'f��u	��	k�q=���	�n���t�g��_~)C�)m'x�L��8��a�36��[�����\
B(���i�I��9��Q��r5t��U�%	����ք!��dH`@��j�`�<�tU��,s�[݋� �B�N�Ui.bASQ��,P.���\�T!Oͦ�-���V��6i��J�o\�8��o������N����x�j�AEh �'s*}p�ɓ3�.�b��*�l�S-C0`�`H(�W����צ���A�u:�� �P������	N�O���|�H�(%��Mv����W#~���������C4���������*���r��xڞQ����`}��%,�ٯLؙZ�m�M��'��'�
���z�Y"%�̤!!d!9��ci����c�;��q���U[�3�<i�eˑF	�VB��{(c�А���bl�W���Q�t͗��>�,�n�(:�ʉ��K>����=��`���`hA��m��>i��|pQ�_�tLͷ�5u���ns�������l�dS�@A1�ڬ��Ox �.c',�d.����i��Zz��ޠ�P}����,NkM�9[�{�ߴ��]:JIw���+T�����Y� ��|$��c�\$���P`Τ��Ǥ��&����t,�8��Kj����z�.�~���7O@M�����5�����p=(��M�C���v�ُ�N��T*u_]�i����F��So�J��a$]\M��<�)�P�c�ͻ��'�F��P�yM�..�m4㱈���[&�V:�c��:<�-!0,��>�
^D�x��ȵ�<#3�1t8]"�N�����L���\��>�P�f��`Q�w��r>�5{9m�ғ�R�ٓ�G��	�GZר�a3yRZӺ�,�&�f2q�U�WWjX�K���r~+Y��.�����k�4���]�
M����+j��8�4l�Ů��p�Z���Z��p�I����k�%]� �H���Cdk
�LD��G�qֆm�h����ֻ��L�� ,:f��ZS3�Z��Y߮�:�ˈ���2����uI'iC:�Ҕ����PL��J;P	ܤY�F�6���{D��@�H/D� o��v'����E��$w���{�X���%����:/9��q�����֓��d�\�a��9P���8ɨ P�_�i��V��X�1�!�Pe0|������^n{�l��z�q.-��SЋW����ˬ��SAUh�?[�g}��a�J�;}�O�5c*�1�"�$��U<�A+[�����SDGFX�c�����xA	YJ���hVAN�D�Zݗ��#}N�6FJ��Q��O�2u-�'](���.�INہ����E�����{��l�-kɵ#	H���c����V���D������?l�,4�2��� �����KZ�~SF�s����4d�9�����"A����JB���ډZP_4V�HeFJi�eΤ�;���}�p ��q�U�DܺU��.X�{��r�7T.?6��tlAU��z�
��P(82��'����4d��\�=>���Wh��%��p��>�xK�y�t%[h�f\v������'���J����4�������$0x�\7wM
�������8Jp��|bj���������UB��KYڴ@�Lݴ���h�������5�t�b�/����9�c�1�ѡ�&��u?�}��Xyy��4���ǘ��J�2〬}D�rrt�3���W��v���3�8���a���;Q,�q"���ҕS����o��f?��ˉ�άyI�t�HY�^�uZsFA_�21�Q���\�>�~Mm��H9D9��@I�|K��Mߣ8�g�O(�x��5�e�y�I�Ez%��H����Gi�؇��{ϴt�>���y,n�M�{�2�/*�*�ާ|�ej�|F�@,5����2~�]I8>Ln��@�4�W�v<l�-�]�!��6Ȃ�͍��ȣ�2zf>m�Ev�@�]f�Q����5斀��s���DLG�p#kb8�i8�.|�3�DC�p��
Im+��Ÿ��-*�y�����1K��RG��eL��1˰k�d}�ꄤ�+�-MN
�%��a�|�{�\1���c���Y>esנs*t�z��V�$��l#e)�n�!)O�[Z�߼��
��rr�E��5�hÂ��]˛*y8H��[@>�����X�C��ɍn�q��q��V b/��.� F���/��^��Us��,y�r�E��KP�\t���Sw_*ʵ�7v2��G�i8������?Ü�a��\p�j�0������D' �\�=���I���]|��? 7K�V��k�"WE����ZM���B���B��6.�)&�brx�yTD�E��q��%�;F\{wreK����ݫ�P-���m���(�%�Sd"��~w��Wv|��M�p�"~���%&z�8���U�)c-!��I����
���(@����8GZCOӖ��U���|�
�4=�?���������Ġޔ���j{o̚���|��#�/�Q�$*�߃7t5l<b'`30�r���B䁹磩g����-k�lݮhxk��$*�[�N<��`$�u�F�Q����v��8R��Ƿy�O���;r���9�n4�e۞ې�o�Ş�Գ�b���j�QW�Ph���oKM<ύ�.m-�!F���h�6\a?Z�����1D��3�1�zr9޻
	;��[�tݞ����>�	3i���Qf˯��\��S#�
( Y��W�R㪤fuUr�o��c��\�5vI�5�,�u���Ĵ�ߖ�JO��������қf>�1TkԹ�����Brg�{���ؔ��=N��sD��%~٤t5�]C��\�QG+&47�n���$G�\n��d+�I�`�ӡL6+/0��!L �\NِR�K	��x�ɜ|�7h����z.��:$��$2����@|�,3���V�3�M�Ve��u�@� yG�-�wtQ
��D�v��\X>��I>Y�_P����J��%�-d�B����Wi(j���$����z�HAX�Ï�A��,��"�6�]�&�F��N�ʅN� ��łEC-6�~��c��q`/K�+�~��������9e�ЧH�+�>�*�'��r�̢)j��X�~�k&�Ĵ�7�j�`�V�&"���N����9���� ����3�;;��ʎ�;����[��T~�b,@�lKv\)��'9�8:��bt�6~����$���Ҋ�<�PZ�T��%�H��(iv�[B@�."�MS�������oz}�s����1���DÓ��cK8\�����i!����X��V�U_�~�x�������*g�Yn�*�*���������)�� =�'�(@����d�m����t�˭�A#�Ev$�<`����暍���HN��Ǔѯs��#�鐘�L�2���؛�l��:�	34%o�r�&3�8�!T{({`�D�;����� x��z�W6\*-W8�:�a�R��P�1�r�dZ��0�?8	�@聸��m��g)��O�i��W~�c������2�76�y���y�󟺨e2���o��K�7�bbi��@�LL�E�SN���@���|Lﯬ�+L*v�:�b%��D�6��թ��Nô�[W�X���+�S�$�x�a\t�q���:*�Xݯ�:��r\<���m�X�_F�<^��[��x�{A��vN���u=5���*5O�� 3=�ۏ_�Ņx ?�q�K���B�-ӝ6���:aQL�ߒP�2F���d򺬫J�PbW+��6X)����I;��%�g�	�H���Hݚ�Y$�7��MÆ����?c_��˜�;����K%\r~�2����#�j
_8�Jl�i%��"�H�Oa�]tZ��I7�t�-�.p��J�6�#�e�NB)-2�6)���s�m�؁�yң�M�9ZSṼWfR�t�z�du�t�c}��1�kEf�f.[ �^�""�B���sj��Z�����|�,F�awj6WL����!*��4f�_�F7<�SE;qL^0��qݎ�y o(yn:�+>�������E�3Q~s~Ǫr�'���q���;�CCR
R�N�����m�g���T:ķ�a�u����e���N��2	����{����2�58����\F�Z��A�*7����[b��YN�9BM����e9���I��s���U�5�j_>��l�?��A��}���/����l쒝�����=����HY"�w������%D����i3,��Vϔ����*<�MD�?x,�4�̹&�䡔��L�W��Oǖ<\͸EV,B��NQJK��iY9��$=��X���շ��v2��ʸ�x#����K��{�{��5G`� �9D�;���E;ΰ[�f�O, ���a
���e�F�@/�d_�;�*�;X�81�X����;#���b�4A�jx)PpKG�,�O�	E=Uj����nһ�N�(s_��	����gi�o4�1�>X�5��[~zx�/�J	z 
�����\�(M�"���9�}�e���-��Ɨ"owi�ה��4�_�r����e��;��K!�L�_��O�ׂ�i �b�2�l���@4�;�7i�X�<�~�H�O���~ʐQ��1���~9�y�_�գc���ږE���t����<J���â�+��Rm:�P3-�����K%R�f�B�k��Mz��ו���A�{�9���l�i7��BǄ�s��g*���6h�fQ�9�՞��$t��QP_r �����)��R$��A�q֮;��X9�-�'�V�DТ0� �r8d{�j��ou���'w��@X ��R�s=��V꼰�� �f�B�>o?=��e��/����j�	ɹ�a�DBw�5�X��x����[��//i\.n��,0خS��#.M��R��ȉ��c`��ׂ�Hh:�hIf�I��Yr� ��$�#bN0��`����m�	?u����;���!�j���,�Wj�C�+x�?�2C��eU�	T֫y)�^Wa�;x1.��ԧ���ha�$��,�0��5��2���3\�GuF���A�\�I ���� 9�*������+�+�3�4�`�nz�`�q�ZE�%,Dw��J�=��1�[�J��8�x�a�����(���C���#I�Y&�s ����iwf�ZԀj?���Eݐk�#�Ec�(s��¥�;�z��? G��gh_߮S�u�1��;��%�1�����f�W�;|q�\q��z�����!���_���/�Wt����`SfPr�Fᘗ�����E�e1��z�󍟛�4�;L�e{:#�F.���~�w���XhS�^�^��R+Q��T�H^
���j^�{Z0B_S[�]@�'�JJ0���30R͖~e���K"|��J�x�����P���=v��P�\�]E�1A3�olşQ�O�����0#X���d�t�E�̇� 7ߊm�rfD0��V�z�WG0����I�׺	I0��3^����ٜ6�}w�'�%�7e�����IU�'�X&�d)˜��5�{" ���F��x0y�+���\�=z�\��_���v��Д�Ѷt_?��wo7֛��|�w�]F'�Y�^_$e�]�YE��pe��;g���|yS��>h�6NO+��MS�3d�d�O�2N�z*���t<�R>�Q�ᢕ�U�w�c�=�����n����M����8��R�b�Z�޳IZ��]5'�3�|�0Ds����1��k>���\�XR\�-��48
���W�瓄����Os� ��g�b�K�=��;�g�������{?�}�qԶ�QSz:cLUN�r�m"{˞U�c"w�O��1 f}�M���y�D2W]UM%����K�J^�@Uo�	L��fJ�����lt���EjC��.3�E��T�d�~g�i�� ���\X"����:UԻ�i��6eW{Y���E� ��Pw��Hi���y5���[8�����P���5)=�q8/�|��n��\�sd,��bL@�۳���Xܠ	��3�Me.���1L@Ps��H2�¨��
��Ha'�B�!����K�UU�v��7�:�7εٛ!�@�)*�	_U�7 b�-:cxTJ��[\�`��\��>�G�d�ܡu��4�������EەG����-� {=���8�;��e����m������.��ژ�hM:�Z�3X=yb!����SR�mi��C<Ê��p�E�sa�;�s!�����4x�ݲ��a�F�.1ŕTVK�u�vo��:�����E_g�:�A��� ��2�&CS��T�a��5.�a:��V�Js��}�FHkͰ��k�' C�D4@w�ڛ�۬I�[��`��B���^N<O����)�gt̏�XF��_�6f/#��#��d�5�*b�S��81$�T�,dZ����m�^L�g~��Ŏ��Į�8,��Ǣ���̄ ��E��G��rm�́� �!���挼N@��Y 9�������E+������|����L*�׏�",9҈�]��"���o?�&(�:��+������?Ĳ˯`ss�(�1M�^r��e=D������A����"���XZX�c�g&D�_�����u��bO��8&:��*�)[����<v�"c�P�㸑�$������w9wO�lVrz�����:`��+��]������iPq��e�.��ڑ���G���9L���~�d��4�z{��V���1y��nG-C�5Jw��I�+���M�hw�:)��=t����rhXA>@وp�����۶��b�<��1K
f9����� ��Z)��K�x��z|�#�L�a��o���-N�_}�%�&O�Ct�M�dkz�ø�i�FỷP�s��妏/��p%�O��)�K�IZ�Ny[K�b��8�6�}�^P@g��s*$��2��n��b��k4�q�_Х������sX �U�(�vS3j�B�����-p�h�|C��X�P '��'+���X6����2Oג/���?q�^�?$DN�������35�R}tf퐜iihl�0���&q�T�d�"Da;�eV#�������%�&�4Mu�e͍�Y9�����TMι�0�����9��h@����u�����FT��o0�ʮ�H�R����=����g��%���ʊQ ������
��Dۊ�)xd��u][cK���Y���E�R��8���=�Lj]ʏ+���vB��\ڤi[P�߼NV7�� -1�3���YC?��k�a�����"�y�ϴ�;(b��^`V�xMhLȹ��,��ʎ��[�9������+�ʧT�
�?Oe����#��1��M���H�P��ft�W����k�QE?7��?��,��d���b�9�h�?�m>�vL�*��?rXa��L�-e<�ݹ��W��TO~�0�A��WA�F.�^���f���J��U�E�(Sf��O�@�#'�?7��X�6^�@��By�F�7�|��{���+���~�!vs�o�	���h����_���w,0�M�QKM����fŕ�7�Lס\g���oŏ�Yˑt��1n~��ύa�[�a������0V� 	��T"So��I��ȇ�g�\�:��t���V��r�c ����\��_��	�,��tI�����1d�KU4ܫư��L�+���:�d0�W�Y�נS8H�i���{[�;�9n.�Xc���;��Lq�ל\�;�dKw�#����8/�du�T���E�\ߚ" �T��u�^L����:�;R�/�:0�h:WK�H���a��a����o�x�0��ƋL%��fn��}��&i=(9�[���a[S���;�G���	ĺ�������n�+�Ns�M�&$�M��m�+�Oi�)2RPdK�%������ƶ��`�����a���d+0���g=�ݠi��A�=�r��/������7�s0O �`U��'���%�Ke���4�O�U6���'�mdCaV�a��K�7����5|d�� F��j�؍q��|�8V�
U�n�_D:���o܂G�S��V�C�A{�Ս���N�i����RZ�j�f��b�}��Kng��=��ϝ@�+�{Df�؜���!��.s����ᒊ�HGCi���#N F$F?�U�^�N7D��aX��Ekx�
�z�x�R��8M�v/�U��W=��<���eV�b����	�´�[�Ѿ6�{�Ύ?é�S�ai�%񩳛#8��2i�	�]!&���~�:cP�����]���Z8?�����D���9�=�����;��a�(�ɔ�V��?���]w,г�U�I�"j2�=����#*��K&¥���\�F�	�}�"���a���1����r�e�_�~�M��;�^���ňk�F��Y�$}2Cw���@����:�*�?�V@�^8�9�-p�����*u����0� ӎ��v'�/�̰y5��,@Kx��k�P�j�"�Z�����|���,��h��)$��"SX��
*W��R�+�V����I��Mg��x�?��riq����𲳚��^���h'}a��UH{�ј�ΦBrpy��&�r!�^�TdA�o�9�UgzT��9m̖j�h�a�]C$C��v'����m؂~�uouA�ADi;^�"����Gf3�.q���r
H��� ��ߜ���Fv���h��@��^ښnM_��b���3��P'��(~AZ�H����8�d����������!& �r��>��Żb��a��vY��Z?Nwb�n!�ְ�s;3w�Dc!
���9�������f���":zw�1��,���|�$^��0�����k|pf��3�*�QvP����l�������U�K��T�[�H�[�UŞF��^h��K�3����wߩp�F�̧���Y`T{^l�t��K¿�}��$J(��wkk��]����Xp�}ڠ�ą�V�	4���i2���+ێa�j�+��i	�& ��x�Y�m�ŶJ��M����M�G���wl���g��ѕ�=>�Ю��H�;���ؚ���i>&����;lC����Z�s�l�]�f��?�DG�$���ʟ�21��"i�K��q���7�GkׂUEց��l��\ŔX�$�@��q��;,@A�g��e�/RQfE�k�J3J}2��S��I?|�׫�p���ȡ�u�oU�[���R��3yR#:�$Ѭ�z�x!�̀c5�����߉ �:gE�t�\��0�{�]�*�B���f��ckG2�?~-��w��;�Q����i�,߉� E3�ǃBx���Qm��㤜�=��F"��>Z��BF�,����#��98=�iS��e����p��(�h���n}�!�xǔ1c=��"Of��3���s�o��UΎ�7\)�I5 ����,����qB����¤]V@�]�W�qYWG�"�]�g���� N�k�t����m/��D�j���%����� 6�C1;�'|w����|Tp��o����GME���������C;�+��v���z��ޠA���i?	ј7����\(��w)u��$��3u9��K>p'��b62��,׾#�Z�~=_��Q�������࠹�}���^n1�L�v ]��L��X�������k��,r��§}�d;��Z2���8��TI*������b��� /⇥�$�X�N]_k�˕!�=�a��~ЂR��-�O��1&��1�Ry�x����1�1-Qx���j_��d��J����u4���B�v��(J��M&
� ��3.�㫒L4%7it�"/���Iy�_�}M��f&�Z� ����@9Z21H�W�<���?H��/;P�P?!m��ӢV�����5� �\��ȆlI ��#�H35�Q�����������J;���g��ᑯ�e��eC�����]��W�����W��xB-b+�j�9�z��U�L���D��Q��a!����f��eC��:J1m�*f9�g��x�pR���D�i�p.�z���_n����t���#� �^rf�a%sޙ�kai+܊>h;�����P?\����k�l�~9G��V���@����{�lжrj�hV��5Em9�.����b��WeQ	_��H�A��0�f���+lW$��uz���!��D1��p̯�"9���� ���sЁ�y�z���m�LL����.l2�"G��{�r?�R`�lS� �ؓ1��9r&I���bE�I��G��>�l�ü ��C1ɯe2O')���r�r$�F��'x1?�]-�3�;��0�g��|�M����5���B���7q�i!ADo�[�Ӱ=:��G�;�Ҩ;l�_n�B�9Ԩ�q<�Zܼz�5�.�.K�����-d_���q�R�1�g����0��Ⱥ�P{�E.�MOQ�_�Ġ�'V��V5��g���r��=�(*�6�L����B�<����կ$ /��Xx@�:C��E���#��!�=?���Օ6"s^��~�� ��D�g<??��7������ �A��������k�c"�ܴ���B6Qz����O�I��`VF�����{|�C5�	�'�Q��wo�~��z\ΈP<��3�K����~�R�ǯ�އ��[�Ix9Ƒ��"t�[t7��h� �thJr�4�I���*�~�7���!����*�WӉ �*�����,���2�M5����)��vg��-c9�	�=��wz�
MX%#�[%��`�a�7�^��ӻ�s|���������Al2������.!�ޱ�XJ����g�W�27T��SEk�@�����ː9�
���u��֜sM�>�����	� ��+4!?8r��]�j���E���T�1o�a��&P+0��%�"��b����:�O@���Z��F���
�ś���-��{�:��m�b�n#E�����Ӭ���*#:sH�T��~���m[%�fd='���W�+9�CG@�̧}ٌd��Ki;'laZ�~������m��������P��Û�4�â�)���L����Uy�v���tw�_em(�r�.�p��B�ZS�6`��8�k(/{���w�rx''����hr�"ч�救�ڬ��|kb2>
�:��&��jzcOAJ�C/u��crXǚ���J��K�:,�ƣ�e�k���s~�Ɠd��H�pn��(&\?|%�$�8���8�UWݑ�,�Q#�\I�(B��k��	�s�h���"��QP�V�s:�6?�Ɗ���D/¼�]���y"�5nZW���u�B�,�>~q��6Z���9��v>����5����.@�������U�I�}D(��T�M��3ba?T�Mq��؆���~#<�5��~�㦨�,-6�U�_��xx/�oyY^q�W>�vQ���`����{��;��Y���>���T��@m>}�s�r?Z,}9����;l��Pf��g0���xC��]�y���%���E�JB�|tz�=�?EcJ���x{]��#u�Y�AE���Q:3�<�Sp('���s:��*�@Ѓ��8�:?��8NS	�>���0_XJlĤ�DZ��rH���kx�@f��{��2,=E�x�_��m?F��8q! ���>�2�F&X��:��<�?_�Чp@�O5��_���		�{����|��g��[`���>�ی�vT�����jzCR�~'�2D�r@����V�wM�r�2����U(lTU�vտ��w��r�����+p���5�I�DN�;E�E$.0��	���"����[	�&�����FL/����v��,����F������[���W1I�?�p`'*����z>!}7A''��BV&�{����F
V��x@AB�#SL�n�%H�:�ؖ���z�׽+6}�g]-t��?�����gy�fZ䍜����.X@"(������[]t��|rɛ��w̒E����闭��i��i�)l�v�b�'��HHۇ����.�r�o��V蚟/=Zx���w㫹��m�!ߋ�g���E�O�⭣�ks�1C*�P�+���/Ɔ� 8���6dX�V�6��S�!�e���jV���٧��D�nu����y��h��i�7V4�͈���u29�O1���uԴꑋ�G���%Y��4$x���U�7�{�S��e��{37XK��z��=b̾��б�5�X<�$����� ��[U�p�9ũ������Zq�/K��P���TYB��I.|���-������Ӥ�N-t���6)��Υ����W�"2�]�t�j�������QS�(�?uc�|$��D�g"Ҵ�����`��x�h�A�=��!#�8Zt��;��E8֓�!a5�̮]���m�����$f\l}�"ǌ.g�����?p+�qLZ�S�%�!���j�h&�{"�E��c��W���[��
JJ���O�_d"�����x�>^�k�T�6�Js��&���j��kB�n��K-��C�*�i�ƻ�Wy~���t��`z��%Ӟ�fZ���7=�oo��%^'w'\�0/����)�݆���Y�O�icZD��s�T_b~��k���uQ���+��Ĺq�g��!$�'��!d3����̑o�}�+��l��� �c���Yc�f6��B�����C+�oƇ�q��~�ZӠ��x`H�K��!�;�W+ı�"�U�qv�{M�U���Kd% r�P��?z�7��c����c����-4̙Z��ݗ����hkʤ��%�Ւ��H�����w��v�ԍ>�ԉ��'d`p��q)vs��G��=�n�;>nG� �"����nr=h�2,��d��,��$5���; 6��>'�hB�������F��Ó[d���8.�*��x�MdI1�Ă����r5KLԟ��&%�a���䍈�
���j)f�[�u��W�7��qS:��}����A�s��h�T����N�J�P�Nvv����
R�w��V�GG��	���Y܊��
,-�)��i�-��K(v�����J�ۜ����*���<F�a=����qP%��Z 	X�ӻ͂��9+3i�]��N,7&__�z�K�r�G^E���fS
r�xM�
	����&ŗ1=Hh�=E~� 
@cvD�T�EH�*WVh >��V׍�W��%gv��U��t%K�쉥]�Hs�ߑғe�eR6�ڡGp�,>���ꔦ*A\��m��֖�����ֿuՆ���߅�]T����,�q@RU'�ª�b�Y�8��m�)ȓ�����5��(+ϙ�t6*��9]b�5 ���36�ܡ�P���v�j#���j6d��8��,Aۓ{��h����ٶG���mIB��2x���x�A���N RGp3��/�S�ۜj�3��=%���:���K��L6�?��ڳc}p_�����$�c*¶`��7+��%,?f���Aֽ�ANV�z�ؐs'�d���	i�d���G�g�e��"CRM���VÇ��7�.K���|���ʪ�M�Y�BBkmW8ޠ��3�X�Qʓ�����8gK��3������L +7����)�D���#��x�Iֽ�#��/��6-��5�����u 2�o��E1}�����HZ�?p�Mkm�/���Q��N֞��oS�Qz>)覺�X0e�^#R&kQc
��[�K~zkQ4]l�O����|/��9�Ra%2�p�|����j�<0��n1Wvk�l�+ �&�ѳb���a���EC~l�7[�;t�iF�FE�l��kU�3�ϻ�Hd�u�\ҙ�.�Ȯ��.��S�+F�Ύ8/,�i��`1+����ZY�����a�?���_�����7� ���S�H1kFYd�W=�Fz)�Bm ��OemP�u����Շ>����.w����UD�b���M� ��8G�4���.�W���`�m�c؎��=�?�6]=3�t8��=1ɥd��(�!�߲jfkK�
�+°�����ǐ�AE�ٱ�L���Q�^2���}p�)���w�3���nU:`]�/������� ]��ӻ� Χ�E��\%�BJ[꩹L?W@Э�8#b���� ˃�4��;u���c�Y�k4��ix��v��C�ކ���8h�� $��\�T���"�v&#A�\6:����z����e�q�S)���$&k�+dÝ"/kf�(�w�1�8�����V�9�_�r��W�w��֮�k���M�}�U�?_up��������r8*���ڙ�]%�u�y��B�D��qӆ�U�l�P'�_o�d���&8��-�r�Q�j/f3��zR �L�!�� ���tM�5�cB��e�ۜv* b�^b\n�`|���xI�ԍkn���S�Q�q���A�kD3c5��O�!��"���y�`���!�G*W�����{�(�y܂ݓ���ė��Y��
A��m~#�'2ŷ���j��y�2wG^!��T%w�~�%� ˘w���u��GX��^������4q �	Ոl�s3�w�@��%�*\��>,)/ح�ᦡ�X������R�	o��u��(��I�i����on��Y��m�6�
c�D������NqPHXH�H���#3%1uDk5�+�^?bs�߰���_�APY`F՝�S����I?��˻:�\����9��G��qX�GȕHh�OfW��說A�>��!Sm}�-����PN{gN_x�Xs���KF���7��'�)"
�7�������[<�®80Jx`t�6�w�=��
�̀�����4f���79���Q��l�bln�7�7Fz�7_�d���ڑ7�"���F-d��{�w�lyCVpt�ouz�U`��V�lE�_l�d��<=�j�N#����tҔj���h�Q"�V������^&L£��	�E�k}�F�^Ƌ-�������̮��I�p�'l͇N�����T��˶��d�-�CJ��)��)�nus���$�%_����b�t]�t�/:�D���)��O`��*9ݔ6h�)$�]j��
���|���i!'J�z!�`tiJ�ȷ��k�B���"�'�q?�`ݞ��>�O��g�'��m�QY�8��͛����	�,!�}w�)�r���6��c։y�y5�ª3��g:�w@9��E�dZWN��y[�Z�^*O��m{�o�b{jb�]�A��al�ߡ�y���X��� �*���>�kv@��E�z�7�HPO�2�;߿�9�HN2�415^K�4'z���g�/����R���v�DM2��[���M�R�0�Y�U;:1�����e�LX�؆+g�[��j̛%��"�m1�r����x��$���癍&?��*g�u�Z�I	���x^�yܙ�������<��f�]X�{u�9;�ɰ(�{S�p��P��]fDV�I�%����8��?��Si��ǔn���?7�j��!��8�ʰ����pVA���P�0�Tj��<5�e;1e]�h\
j��!7a���XK�Z��	�\7��k� 3뭴��|:�Ū�aFd�m����ԷD,��(�`���`����\9�)�唭wׇ4q)2��4K�Gu�PJH|A�[���ܐp��
��@2�APE��m9ԍ�'��me%Qܥ�h���������:��7D	�>eM�
x�9a�t�ZhnV�|���`H4 [L��|�e1��4���չ�=Y�z4Ha��V�=&�A1��Y�(F�y��m�o��f�����Vc��}���>Z���P������YG��,�V���Zo����Ĝ��'�ܠw�G�f9J�PoH��ߖQ�H�[�p����AO�$޲��5	6שA1O��p섟$�-��U�;�$z�Ay~Bۮ�o�;�}`��-��zx����'�6a�4�F���Qg�IA�i�n��=^��>��4���:+':߃Hn�Ǹ?�T
�y���z$r(jA�]j�7���
��:���yd��3{zQ!9��H3�0��}�y�٦�쀐eI�P���Dޢ�c�f2p�06A@(�7�1��>�8��'5W�����Z����D���m>~�-�iٟ5��[e��[>P-�����U���f��>wy��j��B�J�<3�I��I�bo`+�:6��ڜ|>P��u���kMP�x���XS� %�/(�����J�U�$*�ma���mQ|�ųR��V�^A����^��+���D���]���(^$ɢ�;I��0�ej�]��b�Ȫg�BkG���ָU+�a�@�t�I/�X�/3�f8|[�,�^�4JO�9�b��k����{�:po�ձ�5��F٥��1��q)dյ)���;pp����vJ���f�C$H�40�9)d.�C��!�w�f.��v�=�£���m��g1ej�J3dk���d��X�R����K�D��κ�,ӘL~���R6V�Z�PQh�������h�����֋[�L���:Un��j&z��Z9"�W�"��=�s̈́�s��?�igv�g���^�4�Y�s��z��v����Q�R9XW��!���;d�[uӶ-��.O`Z�������J�C�>K��1��2)D��2�L�5^�w%�E�c�� ���W,1�fZJ��ކϽC��l�w��^L�@��e��� ��Ѭ�]G�ҽd��� g���
IgӅ�HZ����!f��⢟���]⹕D�WM��ر�$�J�2�3����Y� t������-�/�n(��CGx���9�j��*���R���kЪ�&y.n'�	Ӎ��fI�5lN�%��U�x�����We�K�w�����fb�����\7��=h$#C�3t.���u��)�ټ)G y�g�%�z����
��DԶН���xߊ8*�z�c��Ks����xBI�:<hj
�%�ϸ�����M�HJ��Y����JV�cx�F�ߧ��Rt�w���}�G���MT�w���P�"��gR��K	�ը{0���hqZ
\��TE{�;�ո�*�4�15{�ni�&O�	Wy(O��!�w˴Q�!�cq|;ـ'���nB�0,3�S��j��bpk7xQ�Ao��膿:9oyÆ���ɷ}xDS��̐���o�K�mߥ`����=��'���~}��3֠���C-��h��Yty~����+�6ov� 2I��ߞp�����?8��'cC�����&"�~��\��f��䇹�7e��E6 휩y5]d�E�+0k�
�0P��A9kv;�[YG�j�&|$�1�^sȦ:u���u���m����� ��3�{x�ߌ��b{�M\|�y�)Ļڹ��|���۱�rU������91�ܪ�;����4(�P��@Zb���_��H&�ɬ٤��
�`�#֭G�ep���7��a~�I�U����ڪv��X5"��w��O�,oŒ��U͊�B;�.����y�3;�f�
65���	Yf�&���s�f*117ެ؂�4�ϾE�%2��7�LD/��	d���"�#S�7��a�wѶ�a�1b�(�Kx+yD6P�y� ��7�}1���Sp�]8����1*a~Q�T��س�f?�/A�X(�:����L��9�i��"3\�}�ݮeIa��]i8E��;�3�p�v2)��ɯga�\��e�.f�2o!�$h�G�1*I�W�G�煛o�l��|�r�W�d��eثZ�n�Iq_~���&C��ޢo~�A�F��/��p�d��f-F�Q��<���SR�[��^��ވ;���Ƒ+�"�s y� �#}�4� ��qݤk*�����k=M}�(�)[ͷ�Xh��q�5�qq���nӗ��1Z�5�%��7DDI�o���P�����&��л��|=RO��>'?�ȗ��BZ���Dr<�w���a�[t)1��o��Y1Veԭ]�d7�P',���讄�$��8܇�V�#�+b��a��3��/�[e�?�L���?�1���m��%P����H�Kʥ��έ<y��EJU��+eU.L�'���Iwo�r3��%=?�(��С{������et�/�C���Q�:�,�SF�|�H�wG11�i��J3�D�iF���)��Ǻr�� �-�@�
�]+SeC�)����A�T�-=����O��'���Ɓ�R�sm>;��y���Hf�k�FQ��0��𿼑���p���5�W�H>, r��&l�/���}���0bҵ^��6��!�����).�����@v�]8[��D+�w�m��O��A��N&�LO������*�.��t�`�-�m�v����#c�8����s��:�u�{8���8�LG/��tM���������=�B�'�uN��.xNf����sFvebjJ4�.2I�Լ��bd��Fnq��o��!h�t���VȦ�0� ?y ��Z9=�٦$�wɻRwH;2hm�Ɯ\m?���.d����V w[�cS�6���N�q5�� }Ԕ���&���@�`\�7��-�9b���V%S���̕!� ��G�Ӊ���@�#^Y�G�.��5�i�5X��%�+����*Q���b�V��('܉�#u�A+�o���ĸ�x���ο�&v��Z�z� Y�JL
���^��W��z�}וâ�,ދ�S���C}'�+U�s܅"H�2�C#�x,� �g����	�f��C��?����9���@�M���2n�s>o�T�т���ѥJ��.��_=�{��Vp[��jZć�?�S;��e�;�
���աk��yC诿�/���	����G_J+W�M�zUF�mU4��j�"Ƞ*พmTGD�梅��5n����a��x"��L�{tfʐ���Ç7{�"�A̬�P��ҋ��� �ΐ��`�({t9����$+ �U���2�2�(��H�aB[���R)��}m+M���oU����O��(��t�����+R�n#���Y���5�&�KB�zY�C0��f���_�F	XPB�,ҍ=�,kT���)w2�����8�V��o4���t�~z<�/˼^���}B�sm��VUv��g;��֎����$Y�Z/�c���fZFK�,�|�� �y
ݧ�e\ٱ��	dl�o�z4�g4�j`E�6i�Ӝ;���ͯlĭ46�Y����C�"����E�o�S~�tսnk/�,!*������â,G�VٮO�v?��~��+�.��ku8}µ���Kd�Ö���@tz{CX�93#u��xw4q(3k�+'�qf?��[�S�ze�/��!;��� L��+0b�6�K�l���n`]��h���2@%Y�i"wr=�(�����?���CK碷�l)L�z��>�@�IY����B�i�5�����/�y�߯�����j�/*�#3��V1���=�IwӶSk�rf7=E!;�����hy���Qǘ���^!���f�f
�ݔc���Fp]c�FDl�z� �tx�c��E���oEqeh���H^�ӼX��E���uq+C�*�J��'�$C�A��.�e�	����<q�KfC9C|�DRaD�4W;�{�E�wT�R�a�Ǖ��p�1P����Ku��O�岫����:��4���?Ԁ%N{ԸG�:�)�Z�3/��2.�3G�Z�&�J�&�2��8c�oq�m�3���I%�V���n]%?�}����6}���R��꧌�½��7��G��hM����	����E��o" ��6��
��2����q����HSE�Fr�U>�mm�)k��\�h,Mْ&���V0�5��c^�7�=r[�6"P��x6�x>-;�a�S�O<����z��7�\�WD�?7{8 �������2��
'�+���ӷ�����
��g���ov�[F�
��f�4�MV�`�d���޳�;�2�f�R��ي
-��ҳOi�M�Ë��#����i����@
��$*�?*�z4%[�h$ƀ�Vש uޖɅ�/Y�6VڧA
�z)!99g�M��q�D�J,<�p�pp20y/o�[�uY�s�5�H��Snh0���ٕ�%+��j K��@��1�0�!s"h�f�M)X��k�|Lߢ@���DRCa9�Ch�U^!6
7��N�-H_�27U���\�G��;}ҠC����!�aû�)�VnO��99���n[i�h*��4��bk����D5Ů ����\���������Qu1G��0<`#���Hm���Rչ�i�-����n���yzss��Qqݟ�W#UR��`�y���bV��] �h!]5ӵ1Nx\P�I��<�l�M>JFeN��Z��擈��;D�E3/O������yh|^���gۇ��b\M��q����'�����ᗜ��> �*�}m�~�Un���S)m꫞�P��&���>|Zǚ'�#ֶ��L��ձ;�52�{|�d�Fb} @= /]�����c���^yG�n��9x�Ù\��R������Ť����ސ�[��c��hf{S�<��@\Wz=ikro�U�B4�I������!#�ֹ-���v ���J���}K�Ƒ"�i
�p$f��ی�O�H���Y��Ƶ�V�ڴh;��b�V���%��{�Q��*ϐi��������u��C�}�	���r*V9�$o
1�����8��k�lc�Wlڡ��C������{����;*�b|�Gpn�w���
����i}g�����So��F[9JV�[s�U�'�]uk2cj.�����&���S�ؙ)�uwG6!�on�[��M�\�i����_`A'�I��z�(�tĥ�r�%,�G�������|Ի��e]��������Ͷn���O��)>^��w��D�=�q����%Y��m1;�W�����L1�)��v��PXX�1�2�ｳ�99�0����S��	W�@�nn§��.����$�Q#Eq��8i=�Bu]�P��[%��' �*@#ʯ2�T�����g4��J"�-�I�j��m��|�ZD�rv,��Xj*?�����`���;���Ҹ[B�~�A
�Ғ��B�U��dr�9��	.^��;�C	Mb��}�!�a�0�l������;��;7$�����z䍚vh�����^��mjm�Y6�:s������<	�;O&�I�)���)�#���U��C~uդ�濡�)5� e]���-�A=*�u�k3��4 #;�P�%�Z���|�.�FM�����a�V�萷h�#�:�B�/���Z>A ����,"JR߫k�n}xO�\��Ĵ6\L��͍:��C�����rA���8���F��Y�$ťe1���A�5'������C�I�����l����$�7���(���m��s���������}�a+���-i�Z�_P�n���":2i;�����	�)B�fV�M���k�����f��/=�tAh�FB�
��!'ʒ����(J�~$�~o�x~�����"&5s�L<ټl�Pv�կb��u�75��4ɖo17���+�ȫ.p:�9�K�bg�V���r�o���y�2m�_���1��kɈ��P9�J�
>�_b�/��l��elv)�P/|�7�;�a����9��1�7� �?KkBI��J��5Df8�e�2rv����U.:��b��G�*YZc��t�7�:zC�Uql�{�d?�/o�x�@�V<�Nwr�c���Ȍֻ���;)n�v�O㻟羨�J��'�*�֢�圏�,l��lJ
�sN>���S�d1K�@z��'��cn"�`�)���?�,��
�̠;#a+]9%�2^���q6�)�d���A���(��=9)c̾~<73��-��)Cjcub��~AT̼�A[LՒ�-\-�U5�)��)vV�W�^!H�nz�0ikO��Z�g�&�ܣ��*lVY�l����^B��@o kg���7a1�j�B8*�����V͙Qc5�l�ǏQn�BǍՐp��!�$�Rp��a�iٙ�^�b��3�H�0ϗ�t?�_+U��7�`ݿg�=u�Vż�2���g'���/�E,�[�
����ؙ	z�����j��j��߳��>�䱰4,�D�3,S�ޒ�Tf$��#8��B�M��^�2�BZ�(���l��	������4��6�YzӦu�H0��R��h�*��U�lo�����V�Cj{�p�0gr] �Ц�~)PL��5:����+kI�De�o�Ph�ύ�Ӈ��\[���`�I�r����(�'PZ������C���o�>'Zx$&���CX뾑@��������d�{�,#�����N�6�Q�� ���^�	��	�k�P��BH����%z��|eb��.,����U~K������+��pf�K��ѝ��N�}�����H&Od��Ddc �ۤg��zPVХ��+���0`�^b=P�~���`Y�6vS�a�y�e�,���0P�T�&�Xd�uF5.#�|dx��z�������+�n�_~!
||4:�2?�ލ�5wա��$���L�i"�iۀ�x�ͯ�����I�3+�u��v痉e��o#�i%�:i�s���8�Vt`����g�9��c`���ꨮ�@j��_�#\ݒ�� ���'G܌�'ߚ��T���؅ar� W�.��b6!��}% 4�P�P��Iu����\� m`w*gג�]ދ-\k�x��y' @���S�e1���n��J�����h	�	aR?1��I�|-Ä�H'0�����ITf��m��-)d7=��3��qx�&���<�q�������K��Z*=���!��&��5xej�"�K,���\%���Z��GN�m�-�V��5��Cg��̾��"�
�g�;��Z�d�/��Q!?Z/��?�t���<�d�z�~|/��[3��Gn��u���xl����?��\�υ@�ؼ�� `B��E�ǀb[ܜ]�rR[f���S�S�e�������P���r��(J���Sv�q}��߈�wd{�Z��������hF���o^�X,�]���3�'0���n���}��_Ǿ���v���Y�eҥ�a��=:�x��'6Ԗ)������y���i��ʳ���!�:�#�KP�.��*͸�'�F">�T����\�����ϧo�5%�
��u1}�Ҿ�$�Yy��G��6U��&mk!����� �Z��Ou�C�A�ؕ��=�&�&�D���P��C*LXt��>��W%�5d�&	����vb����M!`S|��s����0�3-qԬ�zޕ딀o�1�|,jf�΂w�E˖@O�F�N�D�`D��S�/�Ӿj�__}p�V�%x�_]�4����fp��`���r�B��P�A5�k�a7Z�X���y��:z)���z��㽲���?�2�2���J�$��	#�Lrr�9�w#g�A�j�C�W�h�X��-�_V�01��6�U�^"�HA���F�9E��us+U}�Ў_�5o'T���4 ��	���?E�R���\��9ml��G�iOaƷ��7s�Db�����[ȃ�������f��d_�k�|'��Ӻ >�g��lZ�rŁ�Js��
�U����xn	�s�rV��K郛�\�>�	#��,�d�	&��9�^��H�Bl�������b�*��Yoۦ��cN=~��`D���~�����U�}�T��w�y�^�l�u�T�X��;+Q�ó�sv����q}����,�`�qE>�@�Ld�jb��o�*��$sɇ�b������o�&���f��OC
ٙ)����j��L���:  ��$z�o�Y��dG�k;M�ya�x�[��`ʧ�`1X�$�X�>\7�\4,@ �@�Ϙ��s\s��������M��Io�Qvw1���=V��}�9��i��\�%T����?h>� ��m*f�/�4&�Ӏ�@d8�-��)<����syU �����Z�e��kx]�:�A\��>��V,!� �*\�f��yR2�|���#r��7�Ә�}_��~;�j��e��|]��ykc�lo���℡�А˵Ҿ�X��$��Z�q�K��mr�Їh(�L6/�=6���5T�楙|R֗[���Z2�W,���ECP���af��p�g2%����@+�g��:`��U� ����f�Z�V��5Thq���Q7�zH�����'�=���L�:�+����*��:�+��R�i��I���	��<Cx�C3�;�k85�z-L��s��r��u�3|�7�۾� f���p�I��9o�sN2�͞�+h����SQ��Uޓ���ʟᚘ/?(d4c�n�9�d��Z*԰��̲R�
�g4�����2�TO<D�]K��8����h\h�G��v~@���&4*�<e�Y�\�as�a�o�_6l���N	��]�>����'5����J��Z�<�Ms�S����n�r��zr���W�	k�XD����{�ǵ�p�*M�([@�~�"��Wk�.�2�t�$պ���>��>X!!��X�ٛ%�Ji�N6Ǡ��w+�~�hb `0>�:�{�L�0k�O�4�|5=t�C�<
.O��ѹ|�E�����Ն�{��m������V�k+�y8�p)g�ia�,�2�8Ä!��y�Æce��p��:"�(aՌ��I_�4�2"�΍,w��|nf͈������c*��1_�Y.�ݷDA���>6UK"�Q�܂B|��݄�/��Gk�!��ҧ�\=R�aDi&��������mL9�wA�x���w s�|R�ȳL��g�3rup�'�po�����Ļ.7��*����R$��x=p\�_sb�C����'�GF�z�V՟�v_�DM/z�
���؛�׎����N���������bAn���[�_�
�qx�r��|䣎�V?�k¬�T�[��`V���ث
��90���7lVK��n�Ow�]�!-����]n��q�ooToL"�~d�u�J��>4�.0϶���z[�5����������I�
7 l��������kީu(����!늅��0.�H�	��[�_�{�!�"G!��b�6�G%xl�ħ�(��7��/���>,��fs��Nm�۸�'��P����+������{��g5�+/S�,�I�c�S�q��d���>֕��o��{�6�Y?
�1{�f�I����S���w�����e*�{Ĕ��z!)*ʸ�W� �$`�)c���p���A*�0E� 2M�Y�y�������l����D,*�Z���3�W�R�~��S�C��2n|�X�^�LF�϶�m��X�;�"}8�-�.,4e�	#7�VS�˔�&�e��?�p���-Z�6�,f����Su�j�7Hs ��lC�{�Ϊ<�u��S�u7��Z�񙀉�@�Ѭ
�2e�M�rT b ������uRFga�;�6�$�^u�5����m�R��jD�1Ja�e%�#�梒�%�����)M^��t�:	�0��gu��-�����֛��;�k�����c�;������"��"t]��&L�Hz<yD7E���(�^h�k�?�*��	�ܢ��w�(���T�����!Mِ��NH-�����3E�J�BC�l��b�M���V��;"Y���5�7�Ϭ/%~r�T��柼�*�;�VxXˤ�ͩ�~��X�Y����,N`��9]S���#*Vl��e�|:��Zvf�"��]���Ɋ��u���T�G���&�#� PE�	�H`5l���--smއq�z?��*�P�Z9��:���#r��0*���y��LufN��hnKx��~?����b�t|���ΐ\�k�)?$��e0i��3{;�޾R0����������$Yk�]�Q�s�A��g�S��L�0\�~�BQ�F��~i�a������E&��8�1H�@�:����m��8������O
�R���Y4Y\�|u�cTڢ�v�
mf�3k53]�(~`}[��G_w 6��S�^[�U|�h�W�h��g^+T�1�<"+9ʽ�1Y �o�0�_�Tv���3 F��\8�X�^ӊ�Nf�@s�o*2�Ԉ�!}�9�Әd-�����u���
ܲ�b%#A�B���K뽪����j]���a�"���1��fu�[��:37�7*�Q����!cG�*�IgF����W|���<��G�u���Q�b��e�a~��e*Q]�ܸ��"�O�̫U�B&A�;�������\�	���z�=�G.�{f�N~B�'�%��1��ys1�{$9-��"�gӚ\�
 ��׻Ͻ�X����
:�k��et�e��#d��JE���Y�4�6� b�������x��SG}����4�G>��T%�G�H���<�5G�}�1o�����*��ڏ�JoT
��Z-y0>8��}�5o��r�6yթѪ����5�Ʋ$��D
�m�Xgj$�����dOd��b�����Mz��fg�3�.� ���f[���b��UjZ;����2��E�ţG큿���[� #Mo9��)cc5$���:(���[���M�X����4�y����:1���J��
?�^dww�V�fۭ�I�˨�PbuQT&���ROl]���"#���`�0T�$VH�O��;�t�T�,��+"������dX�w��Up�q��Y���Z�3��Ia��I�r��j��Z����+N^*_M�L�������.T�wȫ��a�&DQڲpe���AI1_�a1�l�%�VN��we��y6�����f�!}��DQ�X��*�[��Dŧ�Z:��`��띤�X�F8}H��)K�$b��:.��67J	�H��0�Ti�����EuG�a�~i/|�]�~̘_5>���ҝӶ�-c*��Q�������F�5>�%�/D|��`�_N,��j�]Fi��}1��L��ӈj�供THY�Ѯ�]v��R|Tk0>N�PhLV���g,�lI��8K*���-������ �����]�S[��08�;�a�~�I��L-0��P��	����*;/�N3�&6�P;3ߎޠ�&��,�s��Y4W?$��@϶A�2�Ë &��?:r��͠�4��%�5V�O@:�w������2.�mi)N�@UjQ��2��)�՘�N�R�����k�q�4�g״�)��ŕ
�]�h�MIFY(��|D���j���&A�y��=�Ʃ�%�~�W��I���W�h�%�Y�>��l�Р�qYcP_������'z0;��U����d%�P(�)���B�]i 1а���Q#��G)�%�Ֆ9��qI�e�Po�5�^���$�0��cs���] ���G�#	�Si�8��i�7� �ReS�����9���J 5��/g� }>�E�k���"b�jr[�SC$���V��V�>� dNyR��=���N���cr%}��13;�&����T�,�S���!����w�w	�������ޭT��ִ)�M���$��Hme'�38/���=��*nIwF���>V��[��C.��D���8�fGY/���ܠM�nF����c8PMg��l�m��Ŀ	k��Iդ�'ͪ\��8��)��|-�p��=��^d����}�	t��BF��*qp�����8iA5w����I���R���@Z�m�#/�O������9)oy9�$[h�����D�6�&y{`m�`"6=y��=�N#��]��F����9�aēW�?���=���zh�\��K�H�z����8a _��] Yy9�M�෵�Z\��ZA��X�h��F��s����x<k&��3���y�k�K���>����D��t�ᨹ��KK�8�^Tt�r�����_ A��EeON&h#Hˁ�&�K��C�	Wc.='
����1��h�Mm�	1?M���~���m�����R��z�zL���YE'� k4�6���X�����:a�:~�JV3⚴��/h��<P���~�/p�"�0�1kh�q*P%�MC���n����	�$`&�}�.b��qN��-�����V�5������PI����L0b�ccŽ.ӭV1�&�b���qH���W,bゞdeS.��%HB�j�w��M�B�h���7�P'�r�s�~)�w����`���`94��o�N�Hm�4n��m��+޴��f���n4�W;R�����"����W���)���|��YLW���g�Є�����fQ���<k�k$#�If>�jZ@��ta�B���Q��qv�L(�����*w��L�Kl�w?�Zq�����p�9}����U���U�"�,n;�T���ѝ�E�-3C�"��F�a���"�t�Px��>������?i���G��g�x���S�-я6���h���M��RYP��T|����Q�#�P���jg��˛�������}�h��?�[��;��H1ޖ!F~���Qz,��h�~�˥�YA��V��:;�֟�n�g���·���J�7�W	�'Ǻ��&F���sx��� �"�ى��m��p����l���Rd�rI5Q�0aPh�I���z7�?t-���豤N �R?h)�To�d�K�N�^��k�²��W�{��G�B�M#3�q;�V�MD
I��O)�\l�F����;.��X�da��.n�A:��G�ַ2^d+�/m�e+����ᢍ2s}/g���;.�
��ffi�~�8[�C�)�q!�R�8qЍ'p�}�}K;eJ,Cx0�z�J��S2F���^�ި��������&��1�[�[��dw�a7r�KN�$,)���E�+I���J�x���ϩ:*��8w�99�4+�R������V4U�-{,�.a%�����AE������鰜��	��1��p,D��>׿��˺����k��R|���,j��f6K�1�amڛ>��NZ���>gf7W��9�Z`΋���I̔�:N��5R\�oz�X�j�ޱxrbԥq��儻��f9�fFF�2瞮G�����gI[# 6@n�6��!�jԦ�uA���{ >P��C���4���O�D/z�B��#'jq�|��}F)���0�蝪P�_OfĮe���1�QP���!+������R?�f^E���HC�4�����\mmż��Ӟ�����m�f�ӂT�a!�SF�i,���^���uK~Rv����̓��V|~~��>r�j��S�9�PSQx[�P����)��>{|�Q˘�0u�KG"�p��K�4��S�m��a�
R��B�$�dB�wf@�h�Z�/c�H~���,"�`kB8�Y:0�/8-�%�i ���	�z��ҞZj��)�ӛ)f�O5��I+�r����&���'�+k/��z[���G��99�� v�0��#BWqBE�x[�^�/,�0�����flv6I������}��i��Y�{JMA�ZK�l�vqؚ!~�(v�(�|
�%һ����K,�Δ��~,Z�h&�6��7}@�L1հں����5��`%h�$)2�&��/�w���V��;(g�}�L��q�QɃJ/N����Ҕ��<q�����C?*3�Y©�f�DA{�������fi�+�^�ksf��9=��+��j��G ޞ�@ZƧ<��D�"���\�^z^�: %�A#��Ä��'Fl���0UMOe��{�T�!�K��p�!��	���Փ�~���ÖѶr���kN�s��z0ړ�D�,b�����9�B��ڒ���)�WS=�0&���L�� ��M!����'��U�{���WsU�uǛ�%����F,D$�m��>��|7�4�hJ��,�w��� ����Ֆ���fڜ��nz`x쒗�r˦&�V��d�,�P��kY� �/�B���C"1��;a�a�H��(� H�Zt��]�PD-�bEL�1�u�	��ֈ���k�9�X3�>�W�� _K�w&�)]�߰A�@[�Q�L�NѢu�ƭ=O���(���F�M"{�����z*c+�V�&�����?��\�C������+{��n���K%��Nbr�]X���@RVvmE�\A��̜}�E�Vs1���M$*\�]�%N'ɉլ&6aI��KR��A�VĒ��H�S�G�.��Z*���tm���[9|��	>T��-���gt%������]�|7�[e9�	r�n3���"�b�����GDv�}�(.�Pۍ�4^�4���?F�R����bq�+����G�&Q7Y��Y���{!�1�R�{��VA���՘U�ij���cɹ�x�c�n�}9]'�܆�m�����/�"�i�Gl����l;e,Md��W��zz�Z(�|���j7$]kQCTC~N�;7��=���60�H�(i�_�B$L�.��vL���f.Ą�[����q:�)������9�y�!�YR�3֥��1��I@����O��M��z±X �@N^|E�������a���!-K��a:��T�|��j�a-��I\��QM���]F�g��dyK��rc������eAoq�|�\��[�;&e,M.c��4���F��@?#��������3]�&h����(�%�"Y~9�-���`]������������ef�z"�s���e�Ḷ<}W�,�2,�$��c��)��|V�1�Fmg�����-,OI~)z�p��������������?��޶(sI�v��pj��U�Ħ���C];8H��wdN]|_&�u��Mr�5t;��E�&�wVX�!�;1��1_�:��8؋5�d����My��NK��GpBpa��r�ߞ�#l�O?b:���l���4pH��4F��ǚ��3�m�+��C��)ͬ��@����Q�#/� �9?,�,�i	�����r+8DP���{�	���F��;-
Iq�d�#�z6-b@��#g��Z��="f\��=�wNE.�_����]�~��%'�[�a���(��C�Z�*�����z=o�1"	V3�y"mˤKm-�s�~V�4F�M�����7�}�'E L��؀t�} ���[�1��`o���/�� g��&��\�"8!JQ"�)��Q�� ����,f�$w�kY��]۴ѻꙆx��[Jj�'hZ�n8�II�Qb����K�k��r�/���^Dk������wٴ��}l��I�uJ�Z�����䣩��a��1]�g
�����I8jk9����ӄ3K'����fSr�ƈ��ς���ZJ��8�ap���)t���]!d�8�,���>�_e�\�AeG�XJ���C&��I���̽��}u��>�S�pi�Qf�F틠QNR�2Q��<�
�i��+t9d�|>���w��:�|K!�����*��g8W!g;��@�z��V��#5{���"[��k7�Ԗ�����~�{�$�k`ז8f �*�Hμ�rgY�)�[dMn$N�{�x���#��F�k�E��_H�Y�H�Q��S��b�{�OD��W��nt.��73�����D�7�ob_�xb<��=EM��j?&҉%�1%���v��o6����cz[9�Y�L����]C*�MG���a�y�k�a���`�U���8ꄻ�h�zn���RX��m��7�'��D������!\v&'N`A��@�Jۋ�b�:YV@�����w��v.�HQ���Ŀ�.��RJ���� �N�o��՟���Z������[���CzV��R:ͨ'bԃ�"4�+����]�R�^�WBg��%��8y��$x���8VBd��X�����t�Y��[!Ny�d����>���a��4�dx1�F=~"Wn�N��U'0� �e�\Yx�����r6Ý�I�{���?��\���U?��]!�3=�Us��X��%��I�-��px���|H���}�?炇�
']��E��$r��|�'d��b�sʥQ��'�uq""(W�H�!���C���c/���kY<�,����:���=ǯ��	��,�u���(��Q����>������d%vl�}������L���?G^���?yT>o	�xK��%�,)�W��?=��W0�{��4;��`M$��X�@�v�⊶>䩕�c�F������-c����VU���Є,dkJq� B�W�*�ݮ�R�v�kя�K�	4�M���I!p��&ɥ���ư;�US�E���������h�5F�H/Ă�q�"���2C�BK"XWw����L/+���Ͳ��rg���L22=úCx�=�2�U`��[�O,�K��f��R��NR���]r����B��/��c��ue�;b�&���	��-�b���䩤J}c,��z`��yy��*=��ۅ��(�ާ�L�:n�$� G��X7����	�U�+�����N`��D;��J偖j�
�#X��La2��M��3�t�y�
�>��2�>_�E��i��K��44�S{��ʍ�ǎvb����kn�i4��X�j���oϢC�'�r�jz;�#���ê�7k�)NӼ2�%�Ĵ7y|�����3"51����z?Y��ic�?�����C���~�
��/`�,R�\�G(T������1G�W6�!����"eh���s<���A��;�j0 ��g�̈́�F��rcz��X�)p����ĳg�RZJ)��%}%Z�>h-!O,ӯ/��,�_Lj�qJ���h�Sr�S&���G[��14�3p�F��ˤ3	;�݄d3/�j)���i����$r�I�� -j���O��5!�F�ZAq�Α�mp�U���8�Af���P:۹z�i�h]@aR)i���-�����x�����3d>���z4g�u�QR��\p�N8��L4<�"�x�@�~z�U� 5cX��2��jZ��\���(���δP�Xk-NbE��%��nR2>���V���yV�H���(o�+^E���s�Nٳ���hGN8<�-���;L
���2 �T���9�)�%�V�]VYV��I������`m�h�6�[�G@Jx�C�V�ENwT
l���0�)\
� ^-Al���J���.��I [ب�B�,oO%t^��:D����e~�ܰ�a^��K��������hag�/kWK�x���ǝ%��xxO��n�8H,g�2�pM^1Ӵ.3���v���7��P����K!t�\��ײ�wj_�/�q[3�D�7�Jlr�W�E�����[@Q:�ۮHP;�c��g���X�S��Je�8��mL���,����:A��l��W;+�#"a�F����<1�`�3^�ic�0����s��u`3��K_��S�_�\b��ɮ٨.��u�bX��Sā��$���1y�s����)���j;�1ݱF����Fp�8?OI�\CUWl�)jA�����7G�L8��r��0��}�9��Y���	���a@�ǀ!�R&��\��F��B�����r�p��ϐ���N�8'�*��p���� ��}� K���h�AE�L#W��4��Sg�������������\^�����ٗ@�߀�7`�j��4l��A�3�YJܴ��d\�YNI��W�`�؍Y�E_n_D�����Ã��f�����+ָO�7��o/��S��I����C��ą�|L��s�i�R4�%Y�|��J�N�E|J3�j�}�څo���t��A�G#�4�|l�CԌ٠�^>�{A�_��Hs^[`�gF�Y�F6��--�$ida �X��ާ����_Lb���XϘ5Ҏ�^�@�Of�슄!q6�M��f���o0�p�쵒V˛r$p&��.6�	�%���{Dq��"��[w1��k8�x�p K5���սP�R�{��\�?U���uтD���dib	 �o���+�CYcv����-(�e�̰ќ�)0�3U#2*�3��W���-um�N������GE>��s�zO��`��$ܣ��'���`n��d�N�[6%�3��/"k��VfU=`j����[1N��#@:�����h�f���ҳ���'lfu��?h��0�`DG�ʥ���cA�v< �Ԅ���n���f�k\����w�f���K���~��ц��C��8�Vz�&H,[�����G��QV�k����G�wH9�.`��|�\V؅�u+��2�+�c~�	��/Cm��L-�̐q�U���z�j���[�ۗ�p��%���f��C9�Z�of���ֽu��痊��|�ɋ
�8>Ќ+�����TcQ6��g�)F�FH9���g�G�k�ĥ��tT=�X��\lH��'O��j��jL��B��$�+	���'���i�ej�9�L� N�N�F�y��� G�TE�&$�ϋt��=�W��r(��BmkspB��X�A�p�
��������ٵ�|�9/k�	�G���+�Q����.Q,$o��3����G+��i]$BE�4��<�~8����� ��� ��^7dA.�i�@*I<B��L�RYN��/h�r��h�SCd ˻8y~�k������s���"	�ܛH����=4�/V�T8GޥRt��	�QM�(>W��X-����\��`j_��wif��i$5��J1��g����n���A�Bt��Z���KV���q�-b���RK���Q]G��k���`��X
���k�<�g��$��K���2G"��)X�a��H���+��`�Le�v����9�߰�u���Lcl�v(1G�;���v,�G�~V��j'r9���\�*R� 8{_D�L(^j!O�#+���%��wȸ�W��qC�
���[e��"���ʉ
�Z���(����\�o���sݵ�v�cS/2�1��I����GC]e�-wj��Yc6Ś��a��=	��\?$�[L��:��:�q���OK/+uk�KN	�;]T�g-�*�[�������`�b);r��R	G����G/�y+T�%j1��m��Q#B�+�5j���N��i�`G0�����P �� I��/W=�i���N~nMH����b�):�7�Q��%e7E�y��ϖ޳46���Vػ#1Yo�!(�M� �GC��b�L~]sPق�N/���Hl�����ଈ#�3��e��o-|����r�j�� ��( Ч�� �llj�P �z��2����W�q~��Mu�X=���v�l�l�q/a��
I�xPP�:�/{��;��X��E������2}!=�'��_�pΜ�5D/�Q*��y5o����IY�I��ع��މ[넵�x�?�Ő����}�h2���P%M�|\⍩�ގ/
\�F��@Q�� �ԴxҖ��8�p:(������h�J@�tP�����uY��f	iV�� "u��o���?�fogH���"�7@�ۜ�UG�AH�-�|r�K�G2��컭oȊ��j�ohߩ�H����<5����mO@-�@JV�o� !��qk�+�����5#�s5���1�6˟XH��o|E쭛�3PYfi�/��.���~��K؆V�4Q��L�\up��y=y�;�د��R����UM����;?!�b���m��%5����9])�3�u���2���{2�A���㷈5���Z��J�*�g���8s�b��Rϸ�09�B����������Z�=h3����z���{A�[�����W^%*��V7�_T��I v��o���~_�}wE7[UЗ��!��gRTwI�
�4X�|'P}��,Pu���W�Q�'܀���V�[�n��p.E�kT)�� �r(�C���7M!���N�5�\y}"7���Jy�Ok�K�ã�������X�J�b��|ʢ���m_��h�-1���*wjٞ��4w�(���!Ra�`�1���5�p��tq���Mj.~����-'�!�=�u��kZ�=`Y�Z~���z<�qr�9\S]�|�85��x.�nV^\�k�°�����o�/�e��l��752_�<��=Fw;��}�/��)���E��Q��٪$r=��n.N����β�Q��~��d�� ƦwhT����*�8^�c�����C��H�#t �`���+��Z�U���d�<���-˦Μ�Ye��8�TO^��Fd�1�x��w/3��C��@F�RWA2��h�{��b"���s=����&��<%T����k�j�a�4T�|�������@�y�����&�Y�:LiF��a��9���� .U,�@�Hs��
�%��1�����b�l�D��w�(��'j� ��� X���|��k|�����M��!D2Q��Z|J�r��C�ث���z�Z6�:E;>>$�w��e�x�� ��D�	Hr=�O�˒M��(�w� �ii���!�q�g؟�e�o'|��.��B�4�|"N�Ct�D���ZT�ǥU
F2�#A�$�e�R3I�� �M]%k�Ȉ�A��,�Y܇�ߪ�5:5�w�o,{Y���GM5N��{�X�J�_A"E�E�7W��<���En�^¤_`��N4�A��Y�Q�'8��~�u8X�v��޾��x�C ��|Mb�*��.� @�.2��b�״G��A�\�~=�ro� &r`����4��X��gl�T#�ȕ������+֢�ʉ�,�i���H�������{���q]�� �k��j+D���\�@�]��������0��V8�ڏ�
�� �D��l�E̻&ȗ�SZ��V
ʇ��q0���`�9�1 v���/�u���aQ}{c�	&o����V�����%��~����K�$4:S�y�c�>S���H>�ڶ��f��$��[�� �@1�-�Y�΂�O;vF�|	TU�l����yE=c��Z񲅘�
�\zU���Q3������%� A��|���qW�����;�~����,Rvt^En���ۭ��gnN���I���=T+V��y���C�A�Ɣ	H�����,�!_�J��נo����ǸQS��ý)_�6��)!������I������R�"��P�#˻%�{��s��`�?S�I1g�=��KYM^�e�,�Q�K|�c`-��S�(��|@�Y{N&,�?�#4���N��} �S�~ܾ�	�J�j��f�R�o�N���_�_t�q,��6p�Q71K�.I���Ԑv��m�ۆ	�CNw�'"���ډQ��/7�Ĺ�=5��2�FId���ˊ��rSd�eu>v�Q��x2���4Oޠ�]����(���Y%�-�$���]�%��TfZK���o��������ܸ]W����Pk���p�7-X��5Ԍ�,'ܐ�n
��P&xP�����/~�7�MI����(�IN�o	��T��Hł��M�P��H�0�Қ����($+�v:�K��~�(;��D���8��[a-�����p)W��'׹��}��8A4[`R<�Zw�z`"�|��6#�� ;�cV��_bãt�ڟs�G�g!3�_�w�D+�<K��pȸ�$a��]Ѳ�#�6�N,��eo��b3՚� u��7ؼ����,U٦���@���:Cّ&��Sn��:�0~	F��f�"�ǹ+��n��1�` k�y}2j�I
<�h�h��K����du�a4���C�٬���DX����oTeꂪ�X�E��6K�]�,�J\6��� E��#�O�:>H��-���9�j�}�*�78��K(��e��{\6#��ES]O6.�ߺi+�B�"�Q��)�3'�$�0�F�j`���s��E�N�������!�P�{ w{65hM�-�U���j�+W��f�����fA��B[*�R<͕zO��fS�N��J\3��L����reag�JG#5/�3�m��}��R�B1s�q&]?��w�����]����^/��T6���D5�n
�n"�oV��7��?ܢ���$,��Z8�97��@�E���T0��maeٟg��1�ȅ���ArV����,��g��"����y���8��%�+�!K�%A�JXX[��^ߺ*�����o��M�K�E@e� *6a��n�Q/0��T��n�c�	?h�R)�W|���k��mkt�a�ge����ܪίw���|�1G`�|<�i
疮�G��Nj���j&���:YEp6�}�
��tں�=��'�]��+��V�	� @x�
�^l,�v��7�[Z �΀�Ԯ��`�f�@n�K�$w�!��r���c��V��d�+K�������h��
��<Jp�-Z0_�9_�WH�V%{��o�����Ԝ�ߝ.,�%�;�&3P���9�~��6Iҁ���SG����j����@Ibl�)�߹]�a�����dd�ՄX�Lo���	r.N3u�S��>bo�*"��v@y���{�E?=̈́���,d���Y9�-���-~U��,�O�.� R!q��D���?^�G4�df�:�����Q,>������^��H�[P� dD*�}��~���'#�k�ޱ��UԂ*��܊ ����#���
�1���%H����1�����%�����LN�|'�?��ͅ�a	ܢ/���8�'ݚ�nfcm��O=�y?	�ʹ�q��g�ۗ7�w�r;���%O��`tc�Q�B� �
Q�گ|(���H��,�������!s.`��0k�8-J��*������d�u�ߐ3�����	^�el�Ii�IG�b6"�|-P���?�R����h4�
�#&�sX �	����V�@,:�ݓ��-KbVk�E��w�;��0���@I�_�í`��f�G�ߗ��	u$��3p@*��iǙ4cqU��;k�Mis���T���:9,>`�ۊW恷���� �̬3�6�}��-چZ��ط���� ˽*m�_#�cS�ZG�j a
�1�-yG2����s�gZ'Z�e����Jj��[�i8�**��|�o�!��u;�����G��ձ���_�>���ڜ��[�ycO�ycx�'Y-y���ф����aCXN��V�Yk�'v�x��D<�{9�6E�owti��f|(F4�"�%���-P0� ����v
�2p�FDe�\�·������-��c,�6w]{!PD���Yh�\�YϕpA�3ݾh$�"�f��T�)P��n+�ߤ/�I ��$���xtvd���8 ��Ԛ�j��I��4iݙ{�L:������|}���W���c.-W'<��6��"#S�$�$7gSk;�B�>�i%�"��Z���3�OEa��ܲY�bI[WǓ��g]N8I+JIb�Iv���'r�e��$S7G����fY/)vM� c�g2����q(�/C�ӋF�P�г4X���Q��Ձ>�΀Vˮ�!'�j�̰2kY����)L������������m��zI�q��G��;j�j@�x�_L�Y�t��Қ�G�ׯ��'���)�ϧv�?i"�p�� zW��ؾ�$c)����u�3j!Ħ+s݄�$��7Ny�7�{CJr4Q��PC&ϧt3}��v"ɕ�'p�.������
Q�۷m�p���,.�i�(��(�-5`0y@me_�kMʲ�m�c�G7{�)����F�v���[�9,Ǟ�k�9���9�X�u�.��S�k�@{3�#�}�--"�l6��
8gΜS�	�2L}h}q����.�GgeQ�ۿ?���$�F5(�)���N ���&j50�!P5Ɨ�k��Z�1�>ܟ9�s\�vK���JЛo��f{P+'N1�髲��q��J�6ɤ2N��F ·2b�j9�
�Q�W�9t,�#MU�G�#t7sW8�@��OV�H�|W0�Lb�/��B(p�8����Y����ЫVK�Q@��څF��Ro[��;��=�V&��+T�/�q�8�i;F��rVâ*m?l8�h�8J؍of�'\8�5��e�u��z����ֻu���\qz��fc;��7�a�䡗�l���㛎x�v��[����}*p�� '����������+�jM�(�dh;��<O#U��\2����{�,/;��`(� ��n����k�Y2�0]y��Le��!c�e쁲I�l��ӳf��v���r4v����l����61��we�[��G�n��򛉕�:�s�S�����;��a���Z��5��u����_�$�H��yȽ��2[�`�9U�������Jq d���.u��J�$)��Jr\֬�q/r��	;��`�6LA�?�x����3H��V�u'������jK���m���n/���U+3��c/b�vF$=�a}UW��t�ZS����=h�d�gV�	�~��[߿v�,��"x�EMge&M�Β�np���+|B��5�._���m ���gf,� �Mc�w�ʨ�XM���{���Ñ�jn���Wo� �o�!:iJo�N�2x�J�ꝧQR)n���^��FUA�rfL�
��ni�[�CM��`�|J�kC�uE��1�1�U��L�L��"|��r1��yA��e��;�/�G�1���.����֔���]*��r��;y �j��������R�xi*1v:���n���tP{`���q%!���-q������n�|����M|2�M�گ#�*�<v!E��l��J� ��uM�{f�iB�ߎ�0����c4'��|�2|�j�`��q#^�M�*�Ј��M*'�Djz탸J&���':��m�ߍ̭�%��?5�%�"k������Ss�3�b{k@\�2�y+H0Je?E��N#w~��!b D)��[/_ȽÕ>��Š�`�I�-v&�S��{+�l�_�j��Z��0hp����µ��q��e"I����cU-viP|�a���@�7�c�+������$�wn� ����V��%5R�X�ɠ��&rD���%�p�O��ᛡn�� D���ޓ��K͕n1L��"iEE��Ȉ�#s�����TH�p}�ѸEBln��W/���b�]Rﱥ�I��[Z������B�b��9	me�%�W���4PHc��7�=��V�c�>ǻ��5Ӓ�s��JO䉄m�\ܴ��Z�43��|�\T{nNW����@^&`�=��9)V,a3�u��=��v$O�~H�#$p��x�;HOK�� :�hc��?ak�������^���QK��p��A./|}�]ֶe6�n����1�#����D�C�� ��9���KK��Z2���J�t���T���-������k���V��V���]�k��4�O���^�zci��?���(m���(�%Y �KAb��;����'��YF	U晍�8��[����dn~˰����I��|Z8I/obd�����FeW���6DWl�7�uk�LY}�3'J�ws�K�v�AE[�ؠ��="�c�w�U�"��ڃK�R���C���8�Ӂ!����Iv��-�M���tw��*J�UyJ��d��Oc����;���]�p{ ì��zs���?�}{ &mG�lv'��e������aI5JN̣�e�R\�D�#�e���.0{�RJ�"�o:�V��*vTVxS�U�M����˓�g��I8c��"b��*�G1���s���L.6k*ނ��k������_)�~�i�f����(v�`0�n��0�z�6�k�c��іe��5mʤR�h����UGP��A���o�e�i���w1�N����(2?�U��b�hȬ�:m8q��&���x.C�B2�}�B�THv�����*�r�#6y���}�FL9���AӀ�%aa�ٚ��ZY�}�Z����ת�l3~I�gX��O�����߆d%�iÜa���@C_�cI�h�2��u���n�qtc�i��:�g͹һ+B��W�. �<�#}Iy�UԃX��L���>�T��K�ۯm�i}1�{�O}e����Jw��2qR&�@:�p�>*?���D2��Dv-(��#"�Ҫy:��􆬹n�-�ٮrE��pv���_��T;C����g�\1e�d��O<Y�2iR�;ae�5#�Cw��:�ţ���!9��3����e]�:�w����TST��?5�'$<�!���K$�[ς�xY5���uT�CE�� 2
o�HJYʈ�V�)�~l�*A'�Įkp�UH�s�G]:ￖ`������6y,]X=�q��Xh���y���j9`�Yh���5��xO�ֵ��jq���K��V^=�l���0���`���5Ч[b������уٯ��|��/.C��Dz��1X��e�>R�'�7w_��s΂%��e*�J^p���?l״d��z�<�����拽�z���lئ�4l��Y�)b�Fd��)�#!��"Pau�|���ٰ%�8�.�=&_�{��Q>�s�VM
�FvC f3VI1�xG�I� v��[N��"^n���.��(_�᪭N���
�]۟�ޝzt���h��]b�d�f�.:�7|�����ڷ/1�XS�TU���\��7B�aPP����4�6�3�"�[�����Ɖ[(�e&���Xj��=��� ���Ǻ���;:���L�SGB�4h�������j/����joD�j �}>����DK�\g�	X�L��j�tӭ�,M��9ըF�����OJ���5�	���_���'3����z�/b��&dE�v��S��~L�\�M!��7��j����^m�u��5|�a,Go.�	9�i� �g��q�j�1��ů��i��blӧ/���ckLʤ��!ok2����ٿ�h�\�H�l��.:�~m-�S]3�)	�����gD�P���~H�x?�8Ҝ6���y�у�cF
�/2Z4	K�Se%�;TU-�!���8s�F'�c@~|�$�x2�JVYK+�����5��iۦx<\���������\�����0�s�IL�;��ޗ�P����Kd�����.�Vo6���R�f"O�J8�>]�'�t�]�DMcW�i���!�&���1�|tR}h�����i����n�4V���5z�EB�2���ak)�ȧ���q��^�ȞsSӃE6h��0VC�㥤[��	�p��ɉ3�¬�h��G��~���LV��h�Uტ����so��*��JE�]���yEl�MNH`E�B7t|��&Q�0[z�nȳM?��X�s�(�ϗR��S�ґ�k�>��b��@^����q�Y�F�еj*�R�7\��#:\�T���R�]�����#h�efK��͢�v�.�Q&o|�`�\����J]ڢr�@�9���v�tOޠ9���c�5���v�į����w��_�}Ý�W�K�g���i-n[�ڄڮiw��D>Ƥ�/�dK^؇�DD���d`��\�o7�ថ�����'T�M*�"��ſʼ�0��M�C�XAU�.$�^�ۣ3o3-��D *H��4�Wm��a v�B^,�;�z��>u�I'��m[]��,?J����0�B���ҹ�,b=�At�+�������ž�p�͇=�)��g��g�_;k߂�0N��E�Ȫ.D�����E2,�hx�:�`m��R��r�b �5&�9� �J�Ɣ���H�č:r��85�F������x�Vi�/����U��|Q-Ob��ޜr��÷v{�wu	+�xq5D�/�s]�U�r!
CL���5�1;ey��y`�S}1q|�#(�'T��}�e�?���'�&��c��rǯ�E~�8�q�]g��Qr�*�v� ;�k�,Yw{��_��ὦ�z�p���L��%��/Ұ�.�aN��K�s�⺒�\���8'
��z�&h�8:�IŞ$J?h�p��Y�Et60�:P%������8��FB������)Ԁ�E�]��r��p�6K'T="͡mp�xlr/���u�<���}�bxf�1t
��d'��}��x-+_�P�d{	��m�t�莢�&��O7|熅�ֺԘ���i�!Y�}~�1��zH�`��{���u;l�Y�S��IZ�c�=�����(UY��,cHKm�P�{��F��� s몐��6b{�[����h�boG���^z1�3l�t�n��qQ�T�]
�TzU]`���L�q�)u�;�y��D
-��ޅ�:_���A���AkmR��SuO��þ�I�_<�݉�Z: �N���!�0�.��(����0�tW�jd��^I���c@�hH���.:jV���`����z�07�y�´�04��D�O�ݽEM��y3a$,J�?`����B�;u8ٸ�4K��6�dR�o��g��[	���pv�P�e{E=ڃ{ ��vg��h��v8�)��4�����::D"bװ/m�k���+|qxe��+����V�i���ctg�?�|)��^wU���D����G�e�!:��E; �(�Js��Tr'��em�8#��������jww����j���FU���k�"�_�z;`��bd�a���9�7�Rʇ��p5���jY�����;�;3$:�$�͗\�M�Q���t�,@�G:���ql�H�a��a>�2G*�e��z�[s��i��h�?�:M�6�Ӱ��t�_��%�o�����s�?f�/j]neҙ(t˾�~�R���<W����v��?O��b�U���ɻD�
���h�4�w��'
suX��2j�4��9&��
<^�f�h`'rԕj�1���׷�%������������� 8\�����m�r�jMtW��)�bj���ཌྷ�7Ir��:��"���v=��'@�r%^��0�>��iy~ZL��q��t����"���/֠�������J����)��؎ǲ �B�#?����I6�T��J��RAUi޳�D|{���Q	`�X����m����I�Ʈ���������y��{Ҍ?N�..�@�'8�S���I��+�6u��DE�t��֬��):a�lYx��z���(ء�vtT���PE�(�+q���ҍ�B��-�I��`�[��r:|�x+p�q/	Q2nt1D[1>�2�6�q�/��F)��-됬p)�_�uV����X�k�#����L�W~����Єm�(�6��Ox�uS~D����t�ܖ5�z��1f�o��w�h}Z���$m��N�_fj�B�;�(i{�	6.�"m�9ħܣ�ֲ&����(Yzˬ�H&��(E�d�t�Hf����s��&��l��4��g4�Uw&� p�9�EC�|(Q#8+���&D�����p5t,?��Iq���:4xVQ���HI{�(�[ѩ�e2���U��N��؆�'Q�XZ�޷?uF�c���SZ2(&V�h���F��5��JRHїI러o?�~�е�00
��� ���s<#�˴�S���囓=��)9,U�����"������r%D��X�垴gk(� �{�;��,�}�|Z'�*S�~�$�vg��L�<OU@Gf�Eg�H�4t�+�j5�G/�Φ)	������<ou�u�.���!C���[�\X��&��d�v'�qf�{�Kd.����N���np?ȏp���9�r�����B�:����'�^��H�^5��� O�������eZE�-�a-���O��Z�e���a�"sQǧ���rO����p�b��*��E�	J�Ζ�fL"t��r�#W�&��
��z�JpS�ϋI�Σ6��tq�3�x��d1çR���$�C������(��F�f�T��}$���ʹPlG z��3T<�B�F|�r{ub�O�-��vÄ�Y-^�ӄ1�jR`*�����:�����ޣ�z�톕��=�},�D?qߥ�V��_�D���ߠ�?u�g��RR�Fv��ċ_%����o��)H`]*iŪ�E(m
�H���+C��s�z��hk3��Na� 嘋�l�{%�:oC�U��cz��u"D�c���^�ϗ�"�s�\��cQ5�hRH�� 4�QLѲ�rh0�=RQ芦'$m�MS�gr	 �躆�90�iE�E��H�u�	���},�kP5+A�z^�a�	�K-���xx��S�H�)H���n��&��5|� XQ����xǘC�z8��SX�9A�I�� �>��p�O�|�᧩��cmS���HS_��bR��r�r��,tlǌ<M��}��6�hr�5:�Ge���D�����"�
q-�z���E��N���@��/��Ls�N֤�#ϒ�P�T�7��Y����iv�%�1	�m�`Za�m�Cp�/ߝ�� �Z&~	b�!`ޘ���؀��ђ���(g�E��>����ژ��!`�5�
����j
�=�zh�߈�S�'�A��|N9'%7�D�W��}���5J�����Z���h>{��"�|#�B�[���`Q&�^���������?�	j�B�!�v �I���΂�uC\�,/����fY8N�w�a��Y�¢׺���a��6/����l�6	����~�L�^���e�U ��z;�Bp�4��N�Tof��*��(6�p�Q�,T��΂�Uh	�&)O�?��w ���<���\a7	 2�L��"R@��w����xފ�k���<^#�)��\�4@K'�HP��᭘�~ӂ�~vL;�� ��\���N�}*��9�(�H�V���We_���"��{X�7G�����)$���w:� %��P�~�����g^�ƹy�&n8��-+}3k�h�|����	oz&�S��s�����˰`��?c/+y�F1m��<U�lc��G&������PI?ېX���h���ߛ�G}�ђYf���"6�
�ջ����It�UOg�>�J=ll���>Y��[�^������J�t�O�����@��__*���KU�H�u��?���S�K#Z܄����W��} ����8q��v��¯+�p�Y��|o�%瘥�t���v�q����z��ٍ����%y�5P�ؤ�|��T+�Ԯ�QV�Xe���F�Pyɸ�w����梨J�u߯�����g�/?��Ϧ��������{���n�~�@��H��AvH]�q(W��Y���\A�}�[��T��
�ݯ⭓ے�	Uc�N�[���H=����p�!�ŎXN��ȩ9��'u�t	�a5a+���?�
(�E�b��������aF�][�4þ�S�
�Ҝ�������&�\��g����m�+D��y���Y�A�e�Ͱ~Z�~�;f¨���|��l�<9{W�����8ND���+�>4ދ�I����sf��l�Yף�� _\�v��A��(�ް����x³���(���ѭ�č�[G$o�w����V!��/u��:1�v4�
ב#vZW��[vv��D�W�hm�V"��v�A)�$yQ�|�DV~���>�y������*���)*�W�pX?j����|h��.��_3A�+��� B
"��
��V��T�lUH�anTW�l_� 1�}��d�2�'�-Y6)@&�M�့��i���%����{��S5��Ig(5��9\z� ��z�ޣj6y0����O��3ȑL+�U�y]�䅷�Ґ"�@Vuz��%q�P����I
����4�f�o�;ǩ��2s�Ł�c�Jgn�g00K0	���J�&�J�h}�`+ƣ��Խ�[�I�z$}��w�E>x�~�d�jQN)�z>YB�2�����^��xy�`�s$/py��w�#���J��qn��@#���=��%���w:�(zO�����z
�Р�J/G��8-{�"���F��le�1�a�~���U��Q�Y�������hC D�,�E������3�/�C�7� F8���T�/��\�:����;�0��u_��+�%�)e`ڴ�l�l����{���e�VM{�s���h�̂v�CuSB73Em���*U|��߻��QA��.k��=�]�m�B��7c&K*�e����'Z1���w�a�+���wAU�f��Aˀ �Тf��7;<E�H�(�qF�E�=K�6Ş?waM�AC�7�&�zp:�Cɲd�q8P�M˽}9�vxmy�e�
�`Xc��^��۹�T�>2�Q���,g�o7�r�,i5�泑�Ӗva�9q�%K+�$�s���R"���m.�&u��?�K�b��#��}�5P#D^�Py�����$�NK���uu�6�)�BL����Q�&39���SO������f�8�ki��{�tK������O��W*�ip:#F�9s��/7��w$��_����uٸ��G4ZH�&T��?qt[HO���.\�������Ŋ��Mn/�
8p$��̖�9�m p��F���J����\A����:���l����{M���b��rh�N_x
��*���'���f|����]ꋝ�±��PЅ����� ��#*]����C?�R��lɁ�c)�Qv^Q����{Y?���n�g�K��ϟ1��U]\ro�وT�7;������`ےo�gLYn[����d�4�L��B�}��J�4���op�A*,��<9l�@)�Y��w���@�I��Rv���4}�Y#��*}�`0�Ϭ��i��ƒ	����Fpц#H��Q"�� E���̓��*�@����w��K^=�3b��/����y�>� �o����N5��P�LM+iU>��	*��=�����Uo�۴��J���*B���xr:����?�F��J�՗�I������d���E" =����i7x�%�c{4����Q:e��=����R�����LG��Q�~�rH/���u��ͅ���3U���:7�#��x%έ!�[I�7|��D�� �p��@T�b�0��l�"�?鹮,�T(��j�����M���[<���5�B ;��aE�����7ܨMÁ5zͨ�-8+Y�ʍlҊ������5#�ӆ�D5�?��yv�ѵm#���2�sv��Fp�h<U�[�	�J;m�����0 ��}
&���ɚx�sv-��z�&&��b!��+�!O^�:��-t'?���kx�rh��F!%sT�M�9�f>���!��K��� %Zlnv]i4�}E����Vj�֛�c�,'�
��s<?�nF(�Ia)J�'v�ø���#�|�ZR��sj�g�9g�ˤV�.Ϭ%�UT(�rj��M+��l�[��}U~W��Z۷0W4Ӑc�´��	�O��{rł���?'�[�)&F��%�s}�h�A�};\���e���O�V/�佅�"AO�\��;i��J.�O�3���G �k�皗@�mv�ֵ0�,�jݽ�ik5��!��gS��"i���,�~*�QYBU�P�;�qY3^�\P�F���`V�	y&ū���]tt-��=��f^�2����>]��qT�m�K"�	�rr������Ay�LTq��j����1u-e�?x�4ip��_X~�h��(QT	ȵ�~�'��s���.0w֠����(�����/j�~h'r(�7�|� y��~��򈍈�ZD]�u%r$y�������6pNI�[�E�y⶘jt�},�Vy�j梄6���{�T	N̽��Ĝ���s}q��˖{	s�p�LxU�R0�v�e�*H�m魛�}�@W,�a����� x�4ŧ9�YPW��Ma���!|-s��e�I��[=+�j�	�_��&�����LL���Q�� ����L��e����x�K�)Jq�1^�g36�$ك���43�Ȧ� +�v�l2����P�ߦ�:6��yh\Ty��q��*`�SUDRl�]/�G�dCV��t_�l��kUm*M9H��&�P���˳_�����_�O��5��M��������o+��T�I����3�����&��8�2�j�����0�Z-�E�W+m�{�s�"~�����{�[����Gx�5d0�;ٜN���HG�Ӽ$[��A4eZ�#�'�	P��-3)�`���1B�1z��Hi�t����F��X��uQ�s��v=^ H+'�.�)ńuM��J�nڪV�[~�w�\�+"��G�0�z��&#�;|fW@���n=�{+2��br6}�i�no�֚���3�GV`��tǲu�O��L%3����%�lfL3���Y�o�nk� A��/x�ݦ��6����[7�<4�1�N�F�on�l��i1�_�w��Y��!�C��r3�8��3�I�c�������*d@	ݣ�X�#�D�E����e��K4�����>�g�rU���0g$
�Kt��H��g��ɺR�ߍM���P�ֵ�Z�j��1��Cg�=�K�OU�%��_tYN䟣�ΆՔj�:�ݟ�^�@�-��ށ�E��F\�p6�˹1�MT�e|�RՃ�V+���V��#�Y�؄ݴA7��~Xo�+`��y�5❅ť��ޅ�j��]�
�������o�~��Տg�n�ը��Jf@{MÉ�}>�^���-o�˳��遁��#�]��Z�ɱ��u�jn`:O\�SPM�0x��~S�T����r�K��'�%Ad
�����f~ɉ�xoF�;Y?(������S�h���2%��v&:���ש_#�v���k�fP��g~�5��2�tc�(+���\VR�[�n��������M�Ǯ��4C�����7���\Oؿ���'GT��ɋ��:wB*�==���?;l8N���y��/�3n�E�����Q�r��Z���k�����B[�<��
w
~�`D�����4(ݎ������)X�Ԭ���
��2�gJ���ը�'���TD��b"�԰/�x�/uМiX�0��U���x�*���Q~E9���2��~ ~]v����^��C�J��ϱ���Il�����I01�.�=�:����"��G`+kbp���mNhd��L�ߘ�Ib��bp9Mgx�#�R<�A�J_(uz�8�̂�;,\�B��ԗ�I7���Ҍ�����N���oΏS��MԱ3n;u��1m�!-oTm.��0/��C�?@��ʧ6���L��m���L�@IȐ���&�;K۠߉����]+��|k��n�N�5��T�fU;�8��~�8�x�[J��G��&n��Z.��a��{��� ���#.a�y�W������ ]���9T�2��$V��3�&H�;��N� h�M&p��k����V5�!c�lKGPN3�4,��¬X����àɷ�1!1�A���s�B�0L��ri���$-�
�vf�#n77�Ϯ�K%6�"�H`�\�~�N�����@mvcR��W�m�ą�a��KG�8M�>.sb^��1J�7e���pgQ�e�ә�p�������y����^�Х� x64�f�����I�o�N"$N�nw�1�L�RSf"}Ә|Z��u&����<ݽ+5J��/ޗnz@k����<��#�-�^c;5s�{o���)k5��٨����P�>`:��O Jꐞ��2�,o%��n6��T��7�H6��Zo�AgA{������:C�B�#���p|$nWB(�����$�M�=�iVI����~N�J����
��Co��Q��)����9�Q�n*;(`WS�v��?�[��?~�O �(��X �&����XoJ�u<�#XTU����A�W���.����ƮFܞ�0x�)��5��Ս�T�hƵ-N�\�5��·�T�GK� �o�]J1�r�P8ϗ�����_�%����	�
���{���Ai��"����d��WB�4g���`�"������nJ�ȕ�D�)�!�S�y�n��$E�״�A���!вc�@���ae-�Y�;� ��UL�	�O!�����OB��1z=!����^�l�P�Q~j����u���B�rS��J�����8�]�>��U�����f���ߒ���U�����g�A���T��|���a<�d�<��|^�ٚ����5�"�qWi	��+5�='�dHJ�=���D%.%���'�4����de�h�w���;֓�ؙ�l"���q�y]���]��S��̇v�1��)�>?��
!�3��`��4�����M��d���)� #�ӵ�:������D��ۙw+@F4C�D�N�E�%���U��v���ͻ�/�	�;�T��-OEw���;V`��FM+ѳRϺ��\7�ϗ����SbłU�`3�1}V������1��LJY��Wwg�Ěa���p�H�uOt��%[��OPtR.I�\�Qy����3�k�9�J�v-, �IC�������~iNɎo��ɴQc`,gb˙��g��N*JD�B\>�l�cC�\�#MT}�:������>Λl۵��c��8�1�g��φ�W�˽���u��9x��ϟ��|�YP%�>�J�噤��(D����@N���uk
_�W ����bA+�����Wsƞ�m�K��X��hOB��ǘ�/���}�+�1ַ���3�!�V��i��(�f>��h��_�N8'$���~����y�l<ͩdk��@/��j�È�}<@���ȭ� �w�J��v�N.@��1[t��+$z ����&j�J��\�Zs���"���@��6����O`���=�j�M�syh4����q�d��\�r��'���*��W����#��!Y��߆���Dp֌&��� Q��u$�S��E7o�A�GJv�3|���>� zeَ��sr�%=n���x�(7�\ʅ-�fӦ�\R��cZ�=�6G����� <�W�,�S>{X����݆�80��_�tRy�lU�r �XIX�^�ʅʒ�<�����{YM��u6컅��3���M<Ο��*a��:��}�DC�:t݅-�1��U�e(�d�B�6��3�^�N�e�_��([�R֪�2�|�������7X�^߽<��F/;�=�#b��xa}6Vv�s/�`�-�G�}�@d�f�سｄ���2bC
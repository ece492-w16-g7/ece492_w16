��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d้�^��r-�>��s �8������h�Tw#���#/�x%������N+*z�ăZ�4;L�
�K��R��=!�[���l����yqip5hd�qF��"�(�$��SQs��93ڤ������f����.�:�^o��}�I�ഁU��ۢ:I�V9���|���:�ܲ����n?�6�W�ꠙ�e	m�G6���{Dɨ����0��<��U�K����:%L	ix#c��y�=�8+~Y�Q������mG
z*�̌{�3�Y�~ 4�o����[H�#�r�p�!���.�eLٵ�w���5���߇�(��0������OF�#�C�
�Q��[k/=ʡF O������~p8�л;mq޽�'��\�<a�K��72��4��p�l&A�{�T%���;�@B[��<"`?D5'�q9W*�N�ͷ��M���RO�M�4�����r8�]�y��|�M�ش=知k�<����I�z�k}�X�����������.�;�^�����b�H��L{��j;�Q��֮� t����*����I_'UN��R�����w��:K1=���E��5�yEW��-(�0A��F\�b*��X��mN�M_��*:���3��%0�?�P�Q�(Gv��+�K�Q���A
�|�	�)�{���^_�>�li5E��ˆ�P�M��N��q�!y����"*������o����'	�Q	���x�F��뫛IO#ոs���h�T�,���u: ��v&"M(��F���lKE�=$WQ���6�T�2�:ٯ����%APexRL�J���V
%�������\��p%i{�3��n�!��R����Ϛ���e~q.~�p���]n?^�A@B�p��pg0{�/�ۢ"ɢ���j�y�w�>a���L���f{�k�b�\��L���G�Q���K��p V�-��[����3畨�j��������J�[�o�}�ڕ�����{bjʰ| �%��eE����ř�UA�%ª�;0Ah���Ȁ#�<)�:6|Ӌ���\��Q/�O{��c\#�Y�#MAf�ZՐ���O�`�* �i�g�Q&��O���3L� v�.[FنT�C�k��-��bs��5,b�"B����������Z8,��%��	`�f��B��v���n���F������S-�$N����7 9�h�Z����>~H������O�z�fx�P����J�r� ��H�w>�c��j�*���\�[㞧���5js=U3~�ЛX���;X��.��O)_�D��!au���-��˞}G�:�*��sQœz;����`f�V�}��O\�����Z�-#�M!!@�^֤��l��9C�6�S��N`�A#�JJ[o����ff�G<B������r��Q�@��2��^V�ԍ�-�ޜ��K4�|�k.c���A��(��j&j�O�GHg$��~�GG�Ԁ]����"g��Fc���r�v (r�k�yT3CKgv�M{�j��/�x�OK��J�K��[��I�KS�����HN��/|i7�-ni�D/z�4A��4�n�eO�G�
�7������$�^u~R��Ξ.��fg�$��gOII*��.x��.N�!��M`��=�li5-�<7��y��f��{Fw���y	Bu>t��9�O?���?�
"�n$��.M���,�P�蛎u�^��-��(�A�%��Ϯ^� 	s�*�.��E�an�|����&P�o������V��,��ˏ��}�s��E4bm�=�QK=A4y�`�I�0 N�)hl]�z�@U���Yp��</s��U&�	ת���{uôa�ڰ�L�J�9jT������bјfA�r�D���|�""�^��_���3��ڮ=�.D�=�r`�֏.#I$i��R��Q���+�	�%_A���ft\�%|�H=Z�I��9;�W���Qn�~�q��_Z�+Q"+�^ס-��ȹw���<$����
O�QT?�-z7� �3z�l��]:u�f��N�m�\x���%������+\���)�J�cp�B��sF�g���M�+�D�$�oH��o���CN�0l������y7�'���]Z�| �t� dD�N�]����U5%\��
�lէ V�wŁ�̲��>���:^����D���]��8T�/�3���XvBM��i�a��)� �J=ǑS_�M���G��s���;���O�u�V��L��<E�p��=s�,u���U�����?��S�d��<8��]�q�j@�V�:&��F���ߛ�A�y-��z��ͻ�YvI��e֓�Ы�c���N]����dVl���i�r�����ph�
 }�U�,R4�N8�&��%=,��:�T�[���@�A�s`ê�[���ǃ�;o	0����/)W{x����SϪ�}��.�jb�{�o�*v��lM&��� ܟ���7q�,�-����r��զS�S
�6�H�ؠ��Ƀ�	�^�U(*��i��ԘT�i&7���FN+j���o-{� CdD)�d�v�	%����{������B\�`���1u�rš�ߔ\%&�L�(@y�2�W�ŗ7���ɺZG�1��J�8�_,E^N��������p��y%T8`ʈ$u�D�  ��i���/�rҥǞػ�Y�j5��η,�j�A8�%J�گ -6�xӓ!��?���34�i盳�Y�=���*�Hb�������7]��3�t$L�a�PK����M�Y�K		��A8S���'��b���=������6J��Qd�����*��D8η�oW�0�r�w�0���]���\�j�χXT�)�D�~�Ψ�L�@��x�My;��TiG;*�x����9.�A�Q!3}H�b��c�U�p���n�(�r]�y��!��/+ۨ�}���mP�:�9q��%*�Ŀ�f����	����i������w�$�����0糣�5\
b� ��@�+�-:��	1�\���6��w��تZ9�5ҧ>��+��N��E�[�_��[�����&0��rV��yE����[��E�Z���;�
�l.so��%��;F�����\��e8#c�9����;�A^������3��$������	Y>��Dz|2ؠ���v��2�)i���`i�*`أ%eɗЫY��j�,m�::��rW0dgMGC�6Bl��Ew%?۴��{����]�O��14�*��x)t߶�����(���u�,�n�(��\����ȹ��6-E�8F���x�+�.��$�_��9���W֨2S89���h~��hAǃ��9�\1�������=�\�pی��i�h�*�Y��	��ڔ�%��S�=EZlqOl����L�}�g��)���D6SY�M\����`��"������ �xr�YV$^�]K~�8:�yi~H����Ds�'k�"��PJ����IL�Z�z �ԭ�aX�m+���{�`���.ݎ�5�xD.�c{�O����x����XZ��v�Mf1�Q�N%�*��6ɪ~����Ӽg�lҤ��J>6<����WbM:~�T�r��,inڛ� oD��h|n �n���j�%��Pg3���V�)��on����Vg-�88c��pL� BTY��������<��M���i��	�H�sIpԐ9�BR+˚��8-@sC�͈����l5��Mn�PH:�;c\g�r{d����΢�_��5ĖY�)0���c��Z5,�h�ʔGSU-�&��Xx�e���zS&�o�oS�7�q����x�p�>��@��P����l�/�:h�Z��V>lQ\�Jt��qg��i���L�i)[��߷�>�xӿ-���@MzRYZ=:�򉈩|9�/���P�[]�2�N%�7]�h�k�#����p��>�NV��������ƶfaڟ��Dlnj48��9�������\@��8X�bHLM��YT!�=��T�]<�8 ��ĵ��<��g)w �׭�%���I�2��run�8��Rk,����dv�{���V�^�)J�_��1��&��ԈZ�t�?[F�'^�#BH�2���@��w��
7���"�ӽɬ�1#�4���t͔3 }�l�F���Q�[�nƗ�2?0V�3����Ù���}ɿ�[Eb�ڽ�'NM1��KS�m\��\�柕 E貎��X"�Ȓ+��j�̏��u����!j<�����:wʞQO���?�M���m���&�^�a:�V?3��c� ����1��M>)A0�{��"��Z �� �ta8f��Q�fɦ&���Q1%���"����!׵QQnh����-�C���oYJK�#�a07ѯK�g?�qʒ<�@*0���eU�!��8��B5vKX�G����L���������~0�[-:N
,~0��2���'�׻�V��(���lNϭ����L��z�����Ş�s��fg&D��z�w�n%B�D�*�T/�Z:��o4�R�Ծ�ǖ�
�A������}�Hd w�� _k�Pl��
М�WO��N>�d6�\(��M���rW���"����^�5"�K�?�-*2��O���;���ja�z!dσڳ��c����O����������ՙ�:����ZTDȖ���(�i-��&�qN�RZ����]����`�V�1�E~%qT-fSL>��.����J��C���!�qo?��з)W}忭v� ��	V"��H
�=�}��i/	0P��>�(&0\˹nح��W�Y�V3s!�]s�-s�t��eG�|rW��L+"�/����n
ƅ�upJ5��Я���+�01� 6V�|fG�����_�����\�"�w��|O�3�#����U���YeZP�$K��M9k"�N(���:Ҭ�JMА����Y��Țf��2��FJ�˿�� h{{&�$���R����ݮ\8+_�W0�L.*�/�����Q�����kL���3�D@��43��5c�(R��X��:v�f0!A��/�Pt�g��}�p���6��e�M�f0����y�������
��&�(��Q%�?(�����hu���?0D��jС퉲YR��a��hu$ny�b�L�d+��4�jD�\z���P8[y��cm�S�h��Խ�Yϫ0Md��b%{$)��$}A�����4e�#ە��;�KqsX4��s`�"v�j;n��|�����qZ����
�l���jd�#FQ��`��Y��7��Y�x4��T#h�}.G���N�����	�K>�e�ۨ|��UD���*��&���6�0&�$Ŭ6t}��W�h�P���?#���C2"�!��j�"����GՀ���I�Q����!�R�Iʫ}HY����=k���XO��W�+p�A5��Q�V�����a9���,Hk��t�������Yb�qQ�zF#��R�0A��ŇG��Z�{�E��z%�g��m������ֆ��s��׾��UkR��I$�#��I��a��{�3$}�UP�=�j�ɵ��v,�� ���5�sd��0�>�k�:e���^+�\������ �k�.�aR:�t�2g�׉���qpD�M�DþK��K��(���".��|Xn����?-�P�D=[2C�1�~���!4=߃#ϫ�{F:�G)�A�s�^Ŝ+.�-����y9�J�)��&��}V�`h���7:�i#k�x�{�	���t�t���-݇LO�׫��'F������G���DX�pU��C��G�$%�5~����p���f���2J�U�H��{oZ���>���kg�cOt!���ɡ���ZZ:��aLf�zaP��]!%����)�ԝ'��ԟ�bP~���7[r����1�V�Ϸ�V��M3�M�[ha� .�̣������_��q����d���)�F��ś+zh��u�	��'v\��ƌٽ&
�H���b������ƿɈ'}��W&Ӵh`4V3[�	�p��[�JT���� �������wSp3��L�"RX'o2լ k*�Ԭ����"_m�ZϐHU�+ơ&�4S@<-EǦ�К��E|~|O�� 9,��6_.`ѩ�a�`�t��p��$JM��xE���>����n������~ClJk �L��/.��M7����L�)2�^ZK��#�(�L._��K�:[���e��2���p�!��H�$�#s���0U�+�4����ǧ����?AP&��6�to�e�Y?�
5���fC�1z�S�s9�X��gB�1c:H���?!��<{�%Q�]8���M�
�Py�Dk��ȻJb��u��ޚ��d��;���lr�����-c0�# ������c��VE�!���onő��m�,G����7�ނm?��B)��9���h�e�a���_�_6A�[�>XL2�g�5m�b
�Vd8D;����g7���������Q�&A/����@cz�[ a�k-~�������{.fL>���`�EV�*��߭?�Shh��oO�E�hsP��Sp�7^u�h�������>UwN��a���oPȯ
e;�m�Q����.�SG�z����	⟤ub����RW0/99�����Uegu�_7�����q��Ћ���V^g����K�m��;%S�������蛣�j���x7gΨ��.ἄ/���"oh���~ۍ4Y���@ϟH��Z��g��1yh�Ha�I�Jh�m�ە��P��L?�|�ɭ��٢ld�s�+tY ��k.T��\#�&��5v��I�h�!���VW&�l��S8'kT�j~��+����x�VV��a��c{����c�{}:�%d](²��46��w�4d�E!j�J�4���\�N�tHT>�#�����^d_g��:�[l%��3�$�O�7v�D1�����/з{�nP�>����
Ùk"^�w�w��9>=	�}��4�����v(��&^�fd��@5�,��
5��X�;3��� t����Yj�N��	�����HS߰�(�
:��Ri�!��JN��n�F���b%X*�]�ں�A[���D��pl�č���&?�Zȏ�-�)ƤAx����%�_��9��������`�\���o���E�i�ǰn��쪓�".�����T�ˋN8xKK]��X$�{u����O�#���7���|���8���C�1@������z�s��#q;��b�B ��Φv�s3	�V��~����ê�	�n5zE"u��]+��(��v���Ք<w"���\�ѱ�j5%�/��b�BdK޼n�_�Pb��Xf��ȸ� �Wo�s�w)�cu<e-/�0͝Ao�
�*4�j���cw@�}�<k�b:˄e��y5�`}��Q��7X�v���>6Υ$�W�=�������|p��j��چʎpR�w��D9�3&�8@�>��������V<�D�Rɮt���MV��4>�΋� QM���4�����1�|a2���Q��i\V����1��:��5]J2��<�b�!��Z�����A�(8a0vm�����k������_��%��}^�ʍ[P�f)��-t ��l;Y
����Rm��Qʃ�[A�<4�?}sZ�?�5�*��úc��%�\�1��B�#�(�* ýߋ���<�w�iV�%\�qO��,�AlӮ\Q790q�(1�F��J�j�
e�^�A ��a���t�3Ƣ���1ƣasi
g"���yH����T�P���X?i���D�Q�J.2�Γ��<xI�D��ނ��
��Г�(Ɖ)����ܾ�"|��J�����dA��G$*O5*��Z�A\�m��]I��!��}��i�JӞ����B�S��mC�=��k��N�e����F�c��?Hyg�H�q)�L���#��;��6ţwJd��x�Q���٭��%�׾1AW+��Cz��xrf`Iz�P(ϭT�ys�^�M�B�ߵ�3��k�f9j��<v�{�_Q�c��9�wf�dM�K=�N��ˏ�P�T��%����Hƺ��6��!��Z*�o��6o~E���������i��b�\8���S�B�\(MD7
�eZ�p�Đ_ '�_%iK	��?�t�����p~���h%^bK���k߷6pд����0�#�}���T-n=e=g;ek���	|���B>;H�r:��M�~S��X����ܳJ�W
:��rsp�|rB⾈>�����ׄ�ΗY
^�7�4�4)�H�0���L@1���U��yiW#���Z$&W�<�(��M?ܻ����n>p�&̮���ﴎL�J�A㣉�{c��3a�馱�č��~��' ��&i
�[.KN�86��kV�x�(��}�i*����	��7]�D�
�wŷA��ZT������	bC�h7�VabA��5��M�c��C���u�1��®wN����ȬZ����/i�{�,�c8�	(r�o#n�-ι�|Ca�M�.,(���f;o��6B6E�Iq6��ϠS�_ͼ2��WsZ���s�ŀ[uu�Bs{m���k���O��=�=r,�
o"��R�`D��a���:���|�-�ya�:`j�zډ�����*�]�$���X�`gꅭ	����𦍎���5�����"M��D�g[��}��=]w�!�0���Z����E�Y�����f��1�#g|9া(.�;˄=�0�)�
�Ȑ�_�Y��}�T����/l�[�2����z)/�����3;�G�W$B�����u��6���{�i�1�D	���_	�ԗ5�#�S�	�lf/*�%k���f�J��0.$�z�o���YS����_\UeIWX�C�"��e�շ頳�z�>����֭��!I��<f�/�������H&#V��H=ς�?x�|WzXT�A<L���V�e�#�X�����F�+��bdHyz4&��j����ɩa���(	ѷ��ǥ�q��|���?A���F�P0�^{�_z���J*�J1�#A�(t����.��1tQǞA� ~����|g����h'��K	w�741���[ɶ��˯�E�}Q��Y�\�O��K`�D&a�Ջ4�u>�@�W߄�+/1:3K���.V�%$�/�T7�a�{2q#���������
�P�t��?�?�
K�~C %�Ӈ*Ae"��FR+��!�
-\
a9���qU�ܐp:+,���kF�%�b�ժX^�dY�7��7B�-��;�0��M��:/*�%���1�
=ؓ��i���֥�=c=�����@��?&hS~��3GR^\��a�M�`�f��YS1�'Jqw6�5���ƕ>�������ʐC�Ŧ><D�/�݊�ʇ�����<��՚
�q��u\��Le����$g�d�)����%���}�ƒ.��wr �i���rYj����-��J��}������-�1��u�K̡�F0ֶfa��(�H��:s��#]�G ��Q-����M���_0�||�<��{��E��+��S+X���ũ]ۀ�5r������/�XnN������M
�ںi�Q��k�u�3��-L�re�u���s�2���</�������Q/�� �R���`��K��7G��/p�4h�ң�fg�3*�e�?��:�';Ǭ���W]��{������L���s��4�����nh3���R	�XU�i��t�U-ٕ�F���j������C-�����O�%`\g��,��:[c�{_Iٿɉ'�c�"x������ݒ����(I{�X��f]Ρ�(��y������PM=�O�-�ar����k�C�k>,�CFHP��!��t#��+��	;��Y�yB���X�)rl�J��Ԩ�"��X'���7�C����P�ퟸ+Y"��*_���6�j$4c���K8Ŕ��%rWG�����O�Of7�UF� ��ִ�
v�
�x�*2�?]m����#5j�HxW�=3ލۑ��?����R��j��K.���6�����eԖO|;~u8�H$���/v)�&c���{3܄I}=^ᔜ)/3�е�:GV�p=��ڣ��r��-{�����\�*Z���"��a��Xd�@��R���%cjX��+�����mb^�H~Ȇ��,����5v��4O�ߘ��D�}<l �P�*��&�":�ۃE�{���%�BL6��_�V=�l���8��pV�ň�k�Dv2���D�)t�VC�{VE 4��~�F�b�%ҥ������V���3^N�Y���2����/'���uLF.V*�q�
*bW ���T8�t��/\�\$���,ιH&u@��W:>䂗TK���J��a?�$7=+J�7u?��xl K�GJ�A�����x�^?�k�7��N���i��\���=[Ѣ�B��J��|�ͤ-�8��L"J��^��
=]8 GDtٛ����)�J5�V&J{�i,���r�&�w�ld��6:�/Y��29j��[�{�I�h�H�^�:�0�ce�`��<�rx�;e(ܭ�2zW�t�<a�(�Z�_uxD�Xi:p�\ԇ�ߚ����<+b���t�`
	�K��C�:+E��j*���tJ-)�bԣ���qt,.�f<�H3��&V�}�>���� ����v>���I�-&��(5>�;CfV�tg2���X�3��t̹V�0x�E
pG*w��9�:�]�1F/v�#r�&��M��w��Z�<�pH�&�ש��N��1rv�4[��M�h�#��W��-�/�����|{��"��g�a,-1�Z������MhsN���\}G)X�zY9�v2P�=N�y���CDA/~�vzg��uC"7�A�i,��
8UVW-?��~���2���&��7�̵���YrZ��xeB��Ë&�Eh\��.l�	}��[9#��,��vG�w·d��]�4��SI�P��J�f��3�rH���+_��Pg�(B�ro��H�7a�`Z��O���??��I�����?-�Vkpw�������oDd1XW2V2;����*���Wc>�y�_��Na��&$�ɡ%�Z�c���g-��j���sл��{lb}����%�ֱ@�`�j�PwF����ih����d�=��cFI�s/(�����r4Y�cs� ��q�*���й5��߰�\���bVv��I)l��W%�Is�����ܢk��y� ��^̽3��y]>6a#W�Ͳ�����(ɲ����!��Y#�$?&��?�9�8�;
���h�Q>F�~C�
�IW�Q�f3�D�nT�ĥ��j`bH�:�J�Jek3Ӹ���-pc��ee�w1�$2�Gs ,A�nb�;*��'�+nK���C�\"��h�[��o+u��c���ݞ=K�v@�8Rq�������@dQ��-b�(O�	g`����uǙ8k'{�R��i��-����~�_ŧ�j9y�!��Gˍ���2%�x���̌�Ҝ�F�|m�}�ή�L���!��ru�m)2�}��Ť�׳g���.~˂1�_EW�4�цV+I�S��+��-��~�5DҴ���m��w=��.�_�g��hx]}CuD�������f�u�|�A�r�1-�ן�芑iD�q[��]�5ZuFW�
9i��$v���+��B�LLD���T�N@����-*�@Fiw�<�/$5P-?jYfQtL6��Ge�`,};=t#{�[Ol��ޮ��>A`f�q���].7]���f9��#ݝ��޲��ȳ+�/� Y�I����O�Q
��}يM߂$>�'n�І�Z�7�j������D�a�y�S��+�\�Ҝrj�q�#��X���M�S�\h�@bvy��b�C	1�Bw췤���
%#}ɓ��t���y�]׿[��};����{�7�(1���롍Z�_����n��8;3��O
cti�~��a��l�_���f������|��䐌���6���}$�en��Md;�֘�fɂ�Ix�s��df���;dp�>,��$k#*:�Į�b�{v��1�^�G6�3�q�Z�~��X�F��7-�u�4%
c���a7�t���dl��Y�dWG� a�d��г�ESV�9M"���{0
���u��67F���L �Rxz���C�c�9J�&����Ų4Xl�~G��5����4��y���,k������cm� w[rk�5����S�E�K�@W���/F�nvU@68K��	��N�]B��p7�f6����h�����\ �R�'�6�����tfz�P�t���<ō&E}@�d�)��uw�˺��:^+�.pG�a?#�����qѮ����k1��T����,�J,��$�w���Ą�	�{_'A0r��d,@�М
O]h�H]L�[;1h7�6Cc�ތ�O�pڨwpF���n_�\�s�%�=��i;��[2� x�=�e����k:%DeWd\��;,�B	��̣�8�H�E����΀|�o�8�"�5��+_�wے��z�/9>�5	%�6�y�!|�������q���xM��Q���Z�p�G�+�Z��a��Vx�-�^2�l�*F��[gn:�����P�G��k[��{��Uf�
`OŇůe�W��ܘH��l�~{��t;�+&�-����������2rv�5��-�@�g�%���Vk��q5{ֱ-:�����G��.T���i�D�Pi��@��?ێ���,*�]�9̓�� m�
P���� �r��G�����]5M�Q�����Fv������������9˽��FlE)��-���q�Qf�����K)V�Z��_~@k�O�����7�"_"�U��k�����זw�E�(G6�fC���N�|[�w����?lf<�$_V"E`P�7���	C��!����#c7l�x(��@j4�B������q�W( @�q�k���p��n`j�Ǵ�dcoЦ�_|_
$֊�,��
 ����cF�� n�9�����d)����(_q�gpȩ����Q��
��ק��k5���O��yz�$IPfGD���Pvt(��� 5��GQ[MO����8�ӻ�
�3d*�\��nU�-Ѩ_j�xܼ�4w�6�
4�
���+��u�:z[5���l�H�u��6�DX`����n���`9ݻ pD��-l�K�Zhx�>�_�4�a�U.�SqH"�
�g�T(�e���,&��A�V7r�Ks���\St��H껽v�k�6�*��j�����e��U��_k���K.�Y}����Y��EB�a^X4����}}	��Zަ:p�4g���z���l�=}U�`�
�{�n5H4��zC������@�����O����[��4>�伖���rP�I�?d�\g#y�Η��VP��̖�V�r.��5�@]�6ۣ%��:6�r�'������R��?��l��t_�û���Is����C�9�f0m��.:b����)j����j�nIS�qc?1�i	�97P����F_x��Fd���mSP�QK0x K������|ڃ(1ajdSױe��l�AV�S#,X��**��$k�1�d��]*�}�-�wJ�e�Y��k�kɠ"r�6�@
*|Y�O�����gc��y9:���d C��/ �b����Y��N͊�l��
mJ�0�٨�˧�4:��y�F����nn��3��t�F��$�o�	c�I{xj�9"G5e�SF��9�_3:M ׶�Eh�m]�GG���F��p�LUh�'�ꎱ� &�^CJ�)9��:W��؀��$c3cx�f���Pp�c�:�b�1���G�ӳ$���zxT�&%�*��}��۞�6cmN��si��l��rdH������ϲp�����I>�$��d�Ӊ��
V}�8��h��Ѣ��l`�`��?���
�:+,Z*2v�{VbG���CM����Gշ��8�i���N_赑�d��D��h��i ]ME��N4�M6E��4���$�����O�7���"��M����L��^�l�^�����A�u���q�HEfM���1�o_@}v�J�@n]��RD���[�;y�����1[��DO�Ǵ��$�#�D@��#J��[���h�����4l=�?o�λ�lK����x�����!q[誛�����=S>�6���/E#)5�ݝ�LG�9�4W9�'�k��ؑ�Z��y(����Bq���yL�>��5�El�"#l��!�F�(�<����q�Ү��b�Џ��n,��^�&!x���:cE4
Hj��(6K\>I�O�x�.��2dMy+�]3z��2���5��ɯ����ˎ�J�`�� Е�k!����7M���js՚o?	/6�~HY�X{��b&5�tXl�^\)���o'e�iÎg��������B��m�:;�W�Gv�c9��Ѿw��aO��h;S�[�}TL��!k�6�_���)��bD�yZ��Z�UL�#�D��D�ؐ�G�lmp�M���;+�#ߤ΁��=s>����Ė'{�$;����FVo}�	�92�d��E��ݽ�z�ލ�s�x,�8�����*JL2 ̚hF��b���_7�i�I���dw1y��7fE���څٗ@��]���T�!�W���	~_�}����LuD�I����`(�E���:�$��,I�3?-�����[��ykk�d�l�k�V!�E=fW�K��y<��/��2n�����󖗹[S!�)JO+��v6��R��
�[.���
ҶG��Zcu�D������OX�5m�L͜���$��
���@x�MHOhq2˸}�r�X ��[Iтٜ�fwMFFr�w��A�¤뤖d5�G� 1�#m�\d��9v�?�O���=�#Wi~i���W<Li[�Wfϵ�--|Y8�Nи�#�@�/O�����B�<��!71�z
)�?�t��]Z��DQ#a'�rpԬ���+�2~.f@�tgr]!mh�Ȫ?���-��%t#�oD�'qG|�v	�ٟ�|/\G��{���hK ����tr�q�����ݺE��UN �zL#�:8�z5�dN%�8j��������u���L���\TN��n�E�)��Q�;���zVl�ꦻ"�-�/@�Td���6�
m�	���J�,�9���~t�z����l�mf�|Q�)F-m^�}��	'diXg$���]�xo�5�?Gs�T4U�e�]Ȇ��`�cߊ��k���׋@�Fa�W�c��:�R�F�&��>d�=h	�UU�@-)l�uu]@=g�p7Ҙ�P�
�G��LY��2���Y�#!��:S�3T�IpٹL����b,�b�H�7�Ut�?�w�j�edFݭ�M�x^:��\w����*�����%�5�[�'˗��`h�1�5�\}����F���X0Umz��O���J�x���&�Xz�Z�ͯ$o�8������da�|8�g�Ǡ#���(�&�ǜQ^PX�#��1O��������h1��0󨸡iS��_�s-��f5�MIZ�Ó.� lC�5׋�$�V������S?w⟿���J���Q�gs�ϝ��E�w f�^p�X������m��V�$���%����SC~n�x������Z�P�l�r��X,U��0�Ab,&����F,/,z>UF����-W^�����Z���a6����1G�'�y�����K�U��۫m�=`��d��
zdK�b(7�޸n��q	�.ҡS#b�º��Y�0��k�j�0�+\K�A"8�"�)�`���o�����l���8�M�F�S��7������e�eKʵ�����P����**:�]jbsN^U���֔��Od������p���t�VPl����/"�(@��b�=,�`����Of�1�0l���p��B�d��m4�����g�E�婔��4�׫X��+0O�S�05
��.����ߢYzm�Ա+��N����@Hg��#jߋ�`���v��M$|�����B��o:�+����J		d�Au{䭊��qZ�b�?Pa�ȋ��z>�o�M$�Y@�DP���C&k9W��=E�P4�}}� �хI@1�'���v+�$�-o��@z��{�x�[$ޙ RJ�X��o˙L�J���f!m�Zf�b�R���3�r��|İ��T߉���r�7�x��KT��l��܆(�u7y�m��O�xΤv=�ʄ��Gi	��Q�j�F�xW�k%��Y����w�ך�=N9�@����]��w�������C�<�
g�����5��t��k���䗈|G� %�������q� %/�)�4o5obZ�LK!q�66��	�.�9�*y}!�X���U��.�7O@1PS� �����
��"'���]+DO=�aG0B"�ǽ�y����CxU.�����@����A�!)��l��ࠇ#а���*�0C�� !��߀w`��XT{�YD�t�ӥ�bMx6�/M@�O�4�C� 2�I��hL���'M5�16�k��iv(��&c��`��>s�rt�^�uX ���n�����ޟ�w6�cK���d�]<�v+"�E�ˡ��[�]5� ������\[��	��I	�B��e��p�׌�v1#\Z�����; �]d�T��9
��l4ݾ�7�fp dƪ�O�����=K����DI[zV��C$e�"�IRT�[�k�z(�.�L����e|�./3�c�"!d�$'��^�[���{�-W��]�A��T���Dzn�v�����+3y�$��J��t2��ЈhC�Z����g����O��b��t_��KH"��,����d��J���,j�JS����a\,��娶Ǝ�^9���������@oz
(k�-`�|')i�9��P
�LND��
���'x�էIkV8b�b`�R%1]��߀��˱(�`��ٝ�d�X��n�+FuWLģ<��X���:R(���K&v4nvlɞe��w�$m����f�r�t/��<��U|�QO#�Cf��.�<��0�N��,�r���F�����#�ӪEq�ˏb���ō��M�u		K�Y�� �0����QM�/Q�Ff	���&�1?`�07�ԙ�
�����յzםdOG�0pۮB�/��CA�A�^���ԍ�IE0��H��䢒�D��-*]{V�����c����+����*Ĵ�! ��{�)�_1�9N���t���ݘ*��
��2�
=B�UA����'�c7Y@���?^��nw��ʡ�`�f��0x��.�_i�{0��"��Q�	l�Bff��b��.��3��1��V3ބ�S��b;NA'A������	�"-��2����n�B��TzօG��Y�O)Q�wG*�MC��a�����.����N��(�WC*O�S-�vj:}��/�e������6R���7�Jt�st�-7 ��t��uV��'񻑦'�_�pf�b��`�YK��N+�ӌY�V)���0׊r�� lZ��#F�E��/�gΑ��R4[�G�L�=��'$F"bZ���I�?Ȳ�O�E��j�=�_�e�n�q�J������3K�ǪS0�0T3I#�D@5���Vb?T�Ld�=��+S:,Q%4X��/���ѣ�t�X^�n�ӯn�
��m�d�8�䲹�%��J'WZ��=BҾ���F$�X���eIwf���4+�m���qy�&��ά��Ĝ�e]�`��O����N ��V@��3�{ RZ�.ʢ��.�P���V��z����a��
X��s'�d*H_%�|�hl��{>�ه*��z1�d �$��ف��f�٦m���wݏ�����c>�'I����|j�S�C�0��h����t�9@)��?d��~�R��:��4�;bi�1������&þ�$�6v1���KZ��|j�	ц�B��a�z��+3P�	��s����7�@�We�(��Q҅�K�����{¤��#����rT.�%@���͈�q�}���	9b�#U��	P�RB+���vB������69��]"��`G{��Ȋ!����8(7f/�?���c7�
�mSUl8_�J��_��v^��>2sx�����C��>^:�<:�,	�0��HC�5��H�Y
jX�>9�<�"���>��\mϩ� {�;	2MW�
�)��F��9����4�2l�u�$�a8nF�Q �+�7u�\������7�[�/����'�����fjϧ����\�p�fVVU������LY	Y)���ɑ��P ��p��ڹ���tM�8s��8�>��� �Cnr��j��	��P~�H�� 9��l�H U���+qCخX�dobǦ�%�����LW�)Qj�0����  �h;WyUDl�
��U�LW�|Fn�j�Ld.��	g�|��)��f��As�f��X��M�gK��� ]��U�f`�:v֑�ė�8�����t��p�l@NR�t$}���:.vM��t��N�^9W�na�oXnѥ��������N����m��1\��\���Y��D��t������2��GMл6�����_-�x;��
a`����uA�wG��yyE�U��+�ieT�W�?������Kޢ�6`1��$��Ki����z�9~�����&���,��z[8��:�_FD��Z����n�,<Pw�Q�|9���j��u�1�[n��a�ZJ.�wf:1�'���a�S*`,�-�,r�B+S����ۢ�1$���ML�����	��#l��}�0��ù�C��Y��������p���L�9J���U��(C��o[{*��r>EpPZ���jM&Q�ǇK���_���h�w��j�ԅ�}�R>�f���z�v���B�H�t���̈��	�n��O� ��'��ur�@T�U$��h̄?�P^ي@�-�^�P�ǽ�Ӌ��M�� E��D:uX�����*%-��z
��	���']CM�#}td9�JV �Ј���֘���b��#�����K�������@Y/���̸El��n�]�8�'��Hf���\,�x�k�kb%����?�$���ˆ�Q؊u#��r,�-��Ɯ�ӎ���>��ԡ�ۣ,�I���A�g�1{'i��@k�k���2�\���}F�� ~�G��8��ج�H$�{�)���A���k5T�N�*M�FU���W�LM���6|'���Au�2�Y��gg;�!�E���v`Pj���;ْ)��V�/�mN$��M�X畛e�$V5�Ɣ�έ�H��]����2BXZqVh��RO���S�GO����� �NE!+�pW��'���=b���a��|��*Η��ٝ�]kS��I�c�e丌��蛍���L{��qZ��5O�P��)�y�gV���ذ/!Z��A��,�����rkJy�g��/�?7�u���� "��ˤ0�]��¦z|sȇ���I� ����;|�ƣX�8�v}A'�:`��l���Ft �py?�d���&%H�b�xnHD����5�  ��'-)_G{�X����:�Y�o�|V�ά�?6���#�N��{ �v{&~�yl��F����i�ù��!��ӑ�-����,�����_ ��؆?7[����4[y4D!�5J}���IM�r�W��<K	z�%,F.V�1F�E~����(2-���j�i��Q���\a��RC�0��i1u�T��Sl�,g�I�*��7O6��=Y�V�v�LBx �lxﴬ����m�����)��P���ň�����*�8"���#��f@���E&A��v*�yB����x�ǁY�f�Q�Y�6/�Y�<�m�&K���y�����E�c�B�����O���bJ|�eMV�6����e��7�È�A<;P�m�;iY+hP�+^	e�I�&Q6���xԫ)ϴ4���Et�'��cEdK�9v�nRu�m2��,�Q `��f�sZ��P�2��2�T�B�p���]!' ���'7:r<�b��1�!�W�[=�.`˨��$�I����Y:D��(�{H�āb�ub��q�4��d�:;'����4��
>�N��4�Aׁ�;M��*��^x΀��^uB�zZ�|���w�F�����6f7;���bA��D���F�z9�^��;��ޒ��ȷ�y["���+������@8�Y�P%�B�e�� E�F��6f�}!`(-����Ct����|!���-a;��.���,p�\>Z2.�{�K!�G�M➫�;)�kr=�<o����*Vy bF�9���cx�?�ɱsk�˞���򼙻�]��wI��A�p ��ʯ#�^V�G�vU� ?�-V�g>�ãd�.�N��X_q�kR�W�ӐR|��G��B*�E��9{��Kle���[@�O�H\�̅�0��Ml����?�s�ƀ^�3���A��$�)6ŝ�q��>w��ݑ����� �o�>0/��(�k/�#��ue��G5=���5'U��K�����tC��)�������>s��hp���(�>��� `sF�����M�l.��Er$$��b����UX�
ǷU����~H�]Ll8�B�E�i�7b���v�c�$#QЎy�9>]�ϊX̵�@�\ ���x�ټr����^�ÏC;��(��!��hÎ(<G���@��Kk����t���`�A �5�۟�Ȍ2��;����8o�#��P���r�݂d�^C��en�X�H/�V�R�����u�V4F	Q��W4+�͎%
#�WS������i"۞A)��Q��;�'��-gat�z�s���P�)k\�T���Q�ꕬ;הMJ�����hK�����C;�PF�Gn�W�q��26+�F=9I�x��k}W�OM��7'$��l���:l��*���TyN�eo�v%��J|�;��W;�0~�9e�`y��k|��}�,,g�,�~7�j�0ED�G���n�i��6���8��w>�TG�+�1A3΋󇃪��ǂ��;��	��u���4;{<337����[K���Aw!1x��}Od{Ц#\��'���Qky��f�w�-���Κ£��3[�eZ�,VD���|;����}��Rv��}�@�ΖE�ȟYi�|<�{�˺�)�����}�M�Rʫ��M��#|�>>�=}���-���7z�']=���5��T�J0"aD@y��Uw�eס�54�OI�a=o0�H��p��7�J_6��O�������0��w����.r�
��"̔?���~:)�j�L�+�����N��:��ޢ���'t%8��R����>�Rx�*���eu�� �Z��%���#��<���It�w+�� �v z�+	w��al�^i9�����P�)�x�u촤�;�|�q�a�Fs��K�`�9&j�W��4�����׏VNV4҉)�m�A0;�B�IU|ś�f�J��1�V%nĲ��&l�a����Yiڞ�$Dfۺ�~z$1����V�� �_�H�A5l��
(K��G/��!�
K� �1XG�~`a��)�>b{L�]���WJwY�K�z	���A��֑�)�h���������~ĕ�� �$��/�Ѓ�݂�V�6ǂw�fw �m�d�^�B�芠�zHA#��p� ���a����9wG�n�!���	l`Ky��7�5�I��2܊_,�)w�pȌM ����/H�L��5�v�8���BaNZ?����#�GZ`B̪�L�z*�iӹi}�?3ӄ�����0��t�z����Á�e��3e�g���*�֞茝f�mV�������25	�aڿ1[����0�(ٌ�^W�j�Mkm�V�X:�كS�֞Ex���W"g*Ѻ'�ˎ���
q�<S<��o�nw`��������fHA�وUl�}Z�����Ga������J��?"v�%��A��b�%��]>�N���BI�ŕ
r��a-��~y��t��`�U��~���,��2i�X��u�7ҹ�0+�����f���2�y�eY�~h���(-�b���!�@���M����B4,A���5�R�ǎ�\���[?b,��nF�)���N;��#�nº��sVe�I-	7r�*�
�eNu��w|m�$�Y@KJ�Z$z�E0�Q�I<��H(\ڎ��~�{r�?�b	�;~Y����	�=U�nޒ8��%�0J(�a�&)ʈH�����yva�L7b��2�0\��
��VN�R8,�
�����ÉP���d<�YPX{O�K�2!S߂� ��,;>;��%�[��g$,�B��͢|?);-����4Q�$q���5Vf��L3����̹�6QOB�x����1���sw����������8��f�t������d$Ya��;��=�騀�+J�U5���2��s�iߓf�����t�kuJ�]����
���1����}�t�)���N���_���Z[*V{'�*w���'=��gTR�q��XV���=$!s��zMϽ��c�u�Ud<)1�SM�C�)k٫�&盤
D��� 軸��|�iF��ыN���_����ؕ\��ƻ������E��eF�m*�*7Ԕ��b !�F^a/�gը��EA ���#L��Rݜ�	�����j���O��i�'���r�lĝqUc��Ê���x�t!�W�!����Z���[��߹-6�nZ����f�m�NN��y��|I`fmw����Z�>�zDk�̫}WeK}�L85�e�H@�Oeh+������O^��u�1㘯�6yc��Soe.�*Tg�6b"w���#��y���T���dz��*|,���η�@�$:IES�t%�l���_�Ʈ�~8�I�$�4�������}��xA����a�Odp��W��{��/�?X�IF%��[{Y�}�4��xE�u�Q�:"�ەN"��7B>8�,�|�d���/�%�r�K�������g}M_���δ��!��&�Kv��Fv�E$�����A�<�j
ԃPG�}MŒ�d�� F��K�X�M�Q <�Ԁ��wA7ܞ��g���JS4�!�փ��i�D�K�
ޜ2�,U�'G<͑�3��4�W�)X(݉Y��Ob��],�F��#5�`A��Q�0�p����zH��yE+�Zr���֮�2>ߵ�qe/|����9�G_ ?RfYd�%�� ߟ>�
�׽���}�r���(��h��RsS;�U�Z�)�M��	U��,�g����a���w}�;���c`���O�O����b�+��̏��9G���kJ����5�1ӧ��]�6�!���s��Ǘ}�蛫7��%�}�pu�j�^���Y�ܛ��eA�@(��|@���Kq�dI85�ѲNĐ�4#q3Ci7"M�f��&�8TN<�%wC�1s_Ū��}?��RS*���.�k�Zk�LL�lip8��e������F��^��J?��#۸d����Z��㡰�2�i��'��R֕|;��m���٤��[��-��d��r��#�5e���,�m�ع�Zr��Z�%�Y���[�}9��0��@n_����.�z��<4B����u_�5:`���.�@�>�3h�Ay�j�W�;"�O[�ٶAښ���Sp�����X�Z�Q��S���,H���0��?%s�n�9���>���3��4a�|
&���N`�ߊ���R��`T�L�o}�X�s��=��^�����e�C�Y�d�nH�O�<>�2�?�s�Қ�Q�^v�s��zhL�'�S���V*���������xM��(Y:3���!8��7ko�k��҈�\��d/��QҎ,K�R{� �+��7H��֞d���Ov�{�(A�ִW��sQ�P"�9��������7����&�[���_~)�����@a;ą��b7��cij��7���;imG+>�;�~��eU"d��v����r��	�#�?ŠM�$\��g���w��?FZ�s��({B��	=��0�Iz7��
e� 쇸�ӌ��XD
 )���;��Ե ��H 9��Ʃ��WkG�k��o+YX����KG�!��������J�
�����zJ�����PVolؔ�゜�-� Z18�!RG��5�m(��B}Zx�wʲ���f6�Nz	*�:	�ӎ!1��d
�ڕ�� �q�nګH(:���AQ��)'�ꞯ��fj�{&xҧq��Z��/��(�<9r���n�K9��l�TXD憨mC��ӤU~Hd�)��Vd �0@-�+�����2�9Ɖ�:U��@
]��S�l�j��� �JA��E�R7��F�x�k���@�-ށ�:�r���媿��1A^/�&��L�@] �~�N�>��!|`l����˅���x8Lxl�j�t�ׅ��ݹ�	�w��A�E	�0E�n ��k$�,�g���]�)�r��4���<�UTDm�B,$1/�ᇎ�h���z�t�yM���[b��@@����Ͷ�UX[=�e5v�Dk�-]�
{I8IU��R���C��g6�'��1x��↔����9s#��-�e�J��7X�7���^Qd'�'@��ޙ�`����OSuh���9\�ʵ��$�v=H�n��q/���+Fhܤ�at�ym�+m�1'���@4�ʄ�� �x��⍞�{�.r�D��MV��NVe���ZÇ��M��M$����Ѹ���|�/��9�a���L�lY��r��ޫ��%6��
���xxI#�?���JV�'exsq��Z�.���b�+5݆їS86)��Դ_J��[_�ɍ��Z��9~�*�T'���F�(� -A�:/�#�:W��z��H��2�L�º�yic3>#m�vn#�,*5rd�2g�̔nP[�>�n�����̥���;��u!���72P�>k����5L{�6j�(i0���1��ػ�r=�v����A-�фO`LW��1S'B4-W~��obg��HR;M��1�o'N����ë���@e�����AK`��\��ǡ���z��(��z�Ĝ� }[y�����U�,|,�A"T�!&�1)|~|V����I}�|l��^�z#3bc9^a�)"ѕ�6�E��7�q@`��MB��V-���(F����	IU �����O�ؘ��p�%�rQ�'�)c��4���y���ن7��`H��&����a��0�?���@XIENS��=@q���Ѣx#/�b��iL�9,��􎬉Tr�dbyٷ2��b��hv ��y��5е.?&|����\X��bp�3�ڜ?��M�A_6�E�I����e��^^Вl��q��O�U�eV��2��jf�ocֵ�h9HL�x�A��&dmu�nxέ6��@��-�(�3�E�Y��?ڗ��0j֜�La�V'=�uMrYvwʚ�|y�H>��N�i�9ˍk�'��yw$���Ɋ|�Y��a�}����R7��/�<D�~L
�k���xʢ�#y/��9�ٰ%�4n���a��`*�2�&�P�,j7m3}�\,�𧙵W����=��$n�%Z��pN�2�%�!�{2ql1;��1X����u�%ӗ_�%�."���۾��jQ#�����3Қ;)P��4�xؽ��ű����W��=�K*�0��I����F�8�)=X���h���ڼ��X �d�}N�.!/IP�<O����}�ݪ��WF��M	����	u�T\êE�SFJy���o��+ئ�9-�H�k)Fato��v�u��氢1�
�":l�GOh�"��r�6K����������b� |�{U�_+W_u^�h�M�4r��
�܄1SS�T�S���CJX���@�"�����g�"�pk��;�'HزQV{T�YI{s~�*���G�wJ�;b�֭NL�b�,�^O��ć��c(m�y���rS�'u����51'�A�:j�b|ۄ8R_�VM�ˡY��#^[)��b�%�[��M8yW^=}�ߠU���{ �6���Q*�.)q�G'Gz�̘?p�V;��N�ՙ���&\9��R<)ΐ󊊯��鶁Vo���zI7��[��,Ud�mս5L5����4��j�b�S#R�π�|��?|��wj�H�-��\�%j���@Zܮ�V�^F��f�� �p'�Cr����,�1}?Ѷ��A�>�Γ�����X�[�������Q� E�����`����o��d�Jl�[ hk��4I�)�l������(����@� ~�&[[����cfL!|~�ie�a#w���?�y��[�X���y���+�Ü��d�C��ؗ�&q.�)mo|�TET��ء�-�G�r��b/鹢~�'d���@_u>�:�H耩�;�o<>�O���5[S��n�[	ٟ����TG	Q6���i:��kY�ɒ�}4OX����F���j��\�/�|�Z�o�%�����Hb� ��͗;�J��s���컂s�_ʳ0͏I�/(;�˖Tt��Gc/|F��80�!�-�kظ� �L�(ȁ��/!Ѕt1#LCp�n��c��"t,k%%M\5�Rk�DU;��UU�֐N�0 qM0�f�l�tT�K<�d�lkO��fJ'�bZ�}^�%�r&�T�P����E
+>�!��f,��SH6���E�m:�9�QoQ+�Gf���%e������j7I�nӞ��b�5����ι;��$**E�hj
d�/p��7�ҿ�f4�'��~rW|g��Gז��6�5��ʵ<����j11,c�[sY�j�l���$h���d[����D���K1��͝G~�Z��@���zN���m�j��ǽ�vB��'��g�t΅�$s��;fgHb��EK�0?r�0��vMCK��0���7�Z`ȯ�i�$?�l+�jvD��yw��K���E<���,��{ qEA��v&>[�'��=����	���?��h10���r�'��K��i	br�,�@>��j8\���F��Ƥ>� NP9��![|~y�X��H�G(�o��5I,����'3i`��X�/�:�p��Uy�b.H�ܹ����BԶ�Ac�˔/LF�����z[K��+�8���.y<�&	���Oۜ�eB�4�N���"c�p�?��gl��QjE�L&���~��k�?��?8[S��n��hJ�bx�C�,iFU��S��76g90Ȩ�T�K�l:�D'�.2�Mb�s]�i�u�Ӛ��#��:!����i�u�q����m^��%������|Y�4C�D�g��m��F��`p���N�q¢�F��G4��8gv��R��8-��p��X�[Q�Ge������ 4:���+�TS��{�Eݿ�����q�a3�H$��;��c}v6K���(����SS�٬ �{�pzs�/~�[[�%-l��Z8�C#��&)6�5i��Y|�U���
X��@'tN���R�@䝫a���?J�����=�䉵��T7�0Dz��x�ߗO��L��f���Z�=2o�I��L��p>�yq���3�&s�I��.�:�|�H# wa�;|mG�XX
!39z�E	�g�SDG�$�ûg������9#a=�ii�t�:pw�k)3��kzp�}A��«���Xpq�1�kP�<�5A_=�9�$��8Ӓ���ý`UQ��>��I����%��C;w�KS�BDs�%�0H+��gj̤v^���P^Cv=7(�����+�ga��􂾠�w.�!�Y,x-�;5�l��l���Foڢ<}K��U�>��'*�YAm�̻�����C O��LqAv�I�#F�̯+�*��6-9��d!	�@���oB Ó���5�o� �[��bՇ�v%���݃�_0"-z�.���^�z�� ���bC�E`sP��;�mQЕU��o�<<p���$�*�l�FȿZ�e�o��q? R�ZI-*��� �L
�RR������	y��d����(�>�F������q5�.��8/d<o�>���o��ys��(�����olK��S�q�{����P|�F�B��[29E<�m���.��:�6�׹���Q�����B�^1��b�U{Q�;� ��0,������[I<�=ւ{N��e��V��[��/�k@:�ת;���X��RG�9�n�+y=V��'��@X�T�	��!���'����͕���{�D*6�O��pY���]B,�����U�5u���s��t:�"H�&(��t��ٮ��,�u��[��<��� ��/M�!�Q�p����w��sl��%�T�eɐ�!I񬘵{a�nY��~눸�K�t���:��l���U�A{�Fg��)R�nm87G�q�+��~ft��1�J2�0N__J҅8?m��_ٗ�	vU:��Y%�%(E�\��oA��j,�����<Dq��H������GSM��1 �}��E�S�	)��k����)���RX��Z	Z5���eC��Kl�M	uW��ސ1��mD% �E|�;�f�9�C��Š�xi���?���J��c�����N���͂x)������Zb��E�ﶣ^���w1 2�I���Y8^ʆ��]�(|�A�S��=IaO�LY�Z�B|��S�e��$B#У���۾ ���sw[��/�}��''vN�����5�x�׈ӆ3�U��j߭�;�J9>G&̻�����JQ$k��P��,�&f~W�#0O�ް²�L��e�
�4�aVG
�v5��*�ȗ���,�]��3 K��/Q���E.a�e '��:\�����n^f� w��f|vJؔ�!	o�	���b�ט�{���7n��FVN��'�Kf�տR�haנ6w�ϗ�om�,:>���ک���:JK����"�6����Ď#:���a5�*v�����^"����Zî^��G`��U�	˃�kh�'�L
�����dL��p��FkB���T^2�X&�t���sȓj�	!2q��7�F�E!r�Rrv~�S�Y��m����>�<�ԵY�ʭư�q�q�F��)8XY��f��J
��!ng�)��Mri�q3�D6��:��q��c���K�y-y|U�eL4/>q��0F�����@w�
�oSk*k�ϷN.�$��2��D/��&���"���q�H���SК�*�J����{L�˧�@�þB�.��%����`W�=�p2~(�r;=�����I�dԎݰ�#'*~��]�#/�|Y���T�uU��eky�GC��0eQ�+��g?G���sT����=�n�Z�L�:�Ll������-Y��� ~ � ���Ȇ[���;J�˲����j5i1i}��yl]���x����,�)�Nh�torLqޛ`.A�$ێ>&����f�*��U����ts��F�t(� ��< � ']��c%r�Ok���w�2ɇ�R��%}&����\HZ`����X�De���Bx����߸��W}��@����.;"�NV�6.���
P܌ߖ��:�/k�7]���5�آ��e�c��C�/'�%!n�<�����v��i ��v��`��G(�ra�R����Ʌ-��fc��e����(N��zL��Rߵbo��ĝ���ŵ���n@��3�(�K�VI<�m��.[����w���Q*2R秂���Gҭ��1S���G��"�2<޴���D�������� �R#�!�Q���3	Q0��:�C��7���Ů�;G��w�%>O�:o� _w����UȒ �A ԟ4��6��?.;R��v�Bmc��H�~���� 7_�gӑ�.��M^n����,/����q���+/��{���כ�zw�6�G�Y����~0����U���'dǀ�#ng�͸7��)m�0d/���5 ���'�����Ȗ�-�9���d��-Uz��'fr}��~jDi�*���[fU�o����_x΋g��T%�G��'CB����K��o3��/d5����;�Fw���m�E�Z`�߫��0�|ON��ylN;]����9@�G���8G�_�1���?��Ke7�zJ�����mx��BJ-�2��#��ޛA��h�[��q���F� UH�S��"�Ƽ��4����)��˲	�g�%�fwTX}>����BݷOAh��$�o��NO�K�A����r�Ʃ��A,~
2�7?-Y�?;����%���Z�ُ�+(qd"k�kĹ�Rם�����I���K��Z��5������>����ح��S�7�K��n���x�������d�d����^닂��E�W�,:�HB��fɻsA�)�z�s�W:����;��^`�2���	�)�b�b?����"E��8)�.���:� FO=Ӿ����.�T�!a��ä���@Eώ(H7��93͖�
�ƺi�Z��`��
<�j��5����U��v���M�;�bj\�tUE��si%�w��O�Jd����ǩ�%[�u�S:��RGnan�k���LH�!{����|��]2c�i�x��4N��"�{��+
�=&��R��
<	���<9��j�f�]��AJì��m�O�/i��<��FWVk4)����6�+�Lx>�ѝI愡�å~���,٣��F)&p" K tA��@��.�E�E�go��&����kb����[�Gw1�o����ă����G�BSӷ������C��ɖsmر�uk�W\�^j�~O-�9N��c��aιI����t�MOY��z�^�Fo��ń*�R@Y���q[|q@��y�j����"��W��YA��M=���;ZV����sNQ���kn7uY��]V:,�~�4XV���LHWgQ���IC]�j��)�0s&�"����J)A�K����[	��a�[ӱ�E?`��k1��ė�i��������D�I���*�د'�uH$���/�p[F���ᓠ$��l���]P׸ߩ�[~f^̦�b��E"WW��D�b�I��m��0���x�qU�?���Og��묃��7r�,�벦��Ձ#��v�P�y$��~f�mjܥ �n�t��,�d4�~� Oچ[@�Ѡ~�� �n�U�ގ�-`��%��D�^��ʃ�y�[���q�а黂�_ʓd��!��dR���Ĝ�����>8�f��H5�'� ��dl+r߼zP�O�	U�[p�ƭ�*#���$0�u��Le���B��4*�\�K#c��7"�J4��V�JR"��W��ײ��%j{��O�Br^�?����v����Q�����Z�2��Gxy���I|zԘ�De��!^�B��H���5�h�[�Hl���B�c�
KF6Qf��d'b&T��۸rp��f��G�H��M(�e4"\�-�� �4/"��Y@,6�X��>WA�	���yzh*�#�Swq�N3)��Hɕ~ _hD��ma�%�YH���S�Y��N��r)`9D��R����Q�.�/ez����3��H���F|�A������ot'/f��4#�n�Bԏ�	���Ϋ&	n)}���lH}'54�/��jA��O���ZR�S�2$�B?~�r������F��8l7��yq��646����e2?�e��6��95�Ʉ��q#i��b2'\��T��פ�${+ E@�u]>Ż1F�{��0����f��V}̶6+��fZ�����:���Շ�Oq$٬Py��ծ#1"���X���/����G��!��5�%�6�^�x����@��i�S�h�t�Elo[E��|����168oR]J�B�/f��`:US�Iteá��2����������жW�6%���l�$�X��l����*W�T�� Q�0����I��:P#(Ԩ=c;��mH ��T|�Q�_���|1-�]6���Ţ"�c�L�Dt�[H�>r�[�,��(#	.�h����8e̩�["K�_����U����""A2�y�ꪇ3e���,b��Yzv���u���M_�
T����D.�K �Jh��ќ�>� Aߑ?��?֍��o쌡����ϯ�a�Tդ�Yi�p`PO�:�dS�/���	9�Y4i78��Ǣ}�& �7w
�F	|@��1n�[b��ͧ��ܝG���L_��}����$]xG�u����ҝbh�I$�B>���;Q�%H�81p���IH��<�(���q&�o&��YL����c��E�`N��0�!�xuotpM�[ez]a?jw��60}�:����Ny��?���7��� �M��,�20o��i�g&[GZ��3�f~��v�P��08M���b�����u+�ׯF�$�H�����������~�c��]����C$�||��"s����g�e�ûM���3K�n@u��:ivͳ��L<�l�tT.8��E���V�ޛ��3�_R��\���Ђu�(�C&+&�4�Hd�={+�� w���Hؚ���)Ӯ���'a �K ��S]V�׉E���1�^�'�]>8�����ޟd�q pz<[`u%�gW���^�>��;m��HþX�[ ��z.t7�Q������C�} ��+�Zk��Gi���a�v�1EH?`흁,~�>��Ȍ|^v���^��P2���$)G? �J�9F�������_���@}dUmڕ�m*L+��"O���-ɗfX|[y��Zh�O<���tǈuu�v��Y�Uy�27mt�2�enO&�l��*s,�{�9��U��Ҩ:��,�'y���L�ܗ4���='t���a���.�x'vy�঑C�8`�-�p��xb%�x��_����1y��S�����3H�A�a@M+��M���ˤ0��Bo���g�>]ohU��G��4b_����+\@M��˗-�@��9{���_ͽ�uT�e�W���1�w��$
Ϲ
�j��R���������/�c>G�|;f��o�U#-H`4��7����OC�Lkd��'�{U0&�8 ��3��y�v��ɽ?���Yp-iB�z�z����]�U�/.�	����Ĺړj
�o�9�h�p�����Yzh��k|4���#�͠a(������\C��AE��kn��8�g暵����a�F6n��"����%a�s�.ش�*�WY���*s�n7�&PL|���S���l8o{�,;X�]S�dAW`gG���^>t)k��^��Â����K@g`��!�b����-�����n=`��MrΕqơLB�5cR�0��-k�����^������[�a��zY�V��dY�|�������9��/wP/��o�6�:[��
���6:؜=�9m'k�x�V	�M`�7����<y��̨ �n��Q�v 1�,��m���RT|x����>����_%�Q�JT����~� 7�w��Gb���:��;��bA��p���dQ6a�ly��!����a�%�(#�[aS/�3��M�4�����=���0��᫩V�}�B��ǒ���ϲN�3ũ�Ā��fSߴ�'�+C�I�­�}?�ifg�T�9h���퍸o�H���0W����)��@b>?אm���׎��VA�������o(�Ӎ�%�$�g�v�Ő;��F�H�2��γ_��K���%~!+�QkM��-g�.Q�IE��^�,��h�┕[����T�כ�-�&X�|�Չ�`W����J��@ԸR(��V�y%�eL(���HBj�⢻%�B^�(�� �I�B��+S4b���1���S���[dC(F����������H�ѳ��@D;��m�*SFF�gkL�&b���Ƀ�	��*Y�g"SK3�@1v��<���&<1\�?��%�<�}�/7�@m�C=�"�n`���2f؎�X$��Z��S����!f]�R���_`�R'CY�4����aW����,_>ʇ�2�ht�����I�g���W���i9�v�T����^���(�_���>,�EA�E� �G����� ���	���N�����p]�ћ�c-���M�Dw�e6\G�[�\�}_a��J��ЏYo�@�xs�bD ��5?����Uc_�d7^ΐ�ʁV�����.r;$Bţ�M]����U��DE��tE�ۺI�����B��Š�x����*7q�hf�JrtE�U�@��k�hX�Pb^�w�g�<��j8%E	7�s
*\p��ﯘ�˯��0:L��x#�M;�q2�Qac9���],2�O�	h -���A@W���}�Ds���ǃ�A�q4�n^fI��M�u��5���W�OǙI��()-4�[k��Kք�(��p>���"�"}V�/b�Jk\�U�i��վ��@�3���S�v���:�QFcj��ݥ�տ�!����jO��7Kp�1�jX���ӕ�!��蚍	n:a|�a-�=Ӗo����`0��:��{������o<-�p���Uv$v�;nƒ3��_���5���R�_�:������ �N+����5�X#��/?�ܳq����F�l�X�q��48�Η���]�jt���C|�eЋ�~�G�-��Z �h����r�yw�"3x�Ð����6��Bv&�G^�u	5���/w@���Ɖ6���36�(���\��OZ���*^e����Z���@�8o���Nk��Y)���BG��=�%�g�x�hRRd=���e�fR/u"	q׆�R$�w%r��p���n!0zP,�u^�n�z��Q/{L�̛���]!��s���e���WQ����Y[���f�.��G~M;�+�t�M"%�P����'��<cf����4~º�=���{�uxdO�?�N���Mf��H�MP	�[������&�kz��� �v���l�6\�v._��m�~�Lȹ%Y�ڒt�
�R�x2�pͳ��↱2��7:T�M�V��V���[ :��Cu�ϛ�\:à$�{�A9N�/�����me�"RH����ը���y��&'�RkS�,��[ZLa�7Z�%P ��W�%�/�y9��d]����?�LE?��4:6�{��-b����Y#��-�W��YRr�\��y4��m :G��W�q�<���馐��b2߭��.�X���.L���Q��Z�	:��52��#�U�d��y�5����
%�B]r����*~��K�2�n�f��7b����LH� �!�#L�[x��2��l�8��RC�v0�6�2�]p$�C�|N[���~k�{�1Tt�S�h�*�u�& (rM��p"7z-һ������wM�w=?ST�h�FH�`�q~<�G:,d�p��������'��zd\TA͠N1cm��d�
5\�1
��\���87�Z�g�s�0�ߖ{�����ދ�ꠄ1���c��nӼ���$Ly��S��kC砜XY _�9"_�C�y���]x�)�����c�ֿ�wz����YS�K	�C���j�f�% k��E<(:���������p��b�Bs�����'�t��b��J0��E�h���<,�u�D?��p0B�mBK�Ћ,�Bœk����q�7���ѳ��|[��=�}�����d��?�=:~���n��oT�Ȗ~yͶ�G?�h��&A�]�5�ŵHx����
�=��#Ŭ_�sGK����8��/u���M-n�暴�=�q4����}�8M�"�_L0�I���'�� s�,�H�]�ĵ��x��1�����lƖ2�&�p�a.�it7Z�x2���x\�|{n��K��H�f
��qW��3:��B[o򈬕��g�`�?���ׄ�(�d`�˔��ǁ3θ�\_]JVr|50����sλ�p�ԂY�5�%L�Ta�������~����{��?��a��O#�p.��AzAco�DT��YL,B�s;ꁘ�K��,�g@���՞NG`�˄�;�C$��x Z&L�L��M�y�R]������&��0��D?���|�3#�ݩ4�=�G��W���z�;��;������d��;2u���yj( n�_��%�8R���$����>��gm�	��=���(�L_�����i0`������ ��>A���%OY
̗;8��Q�&Ta�<M����큫��~W��#��������M�@D���	���H~FŘm�J�D�I�\k��Y_ @� ��ؾ�
t����E=��q�֙���l	��X���q8y�T̹�i����Z�.
!/���u#8���gA���s2Ǆd�5{�g���D�P�=ޯ|����n������)�o��N�A�MF͝���iЦ�-=  >;-GV&�լ��%��X\0А}Q��v���OڶC�Aw]�R��ѩ�:o�g�O�@f�*u��m���>��g�(� ��:Ś_|��5b|b������HmSP!�F�Й��i��k��j���Lo���i�YQ��'hJ��"�΍��ZI�k�}v.%v�Y_��Y��7=l0�aq�����o��ԧ"�HG��U�|�:����Թ�6&����\es"���I�>lN��F��>]�V�؞�IA��V�˒�G���/���0�%�
�n�\���ؐ�9��_����w�f�ݵ�0���e����x�.��1��>:�k����F�e�j0��f�=�P���~F���[�Ɩ�(�w��ϱ����w��=�����bͿ��{Z�~��G������z��ނg
�) ��cjn�Uo�(����g��	�<��N'oMUJ��.#ַIVhe[w�P�`�.���ђ?\[�8C�ܛ� i���F?Y̙!�t��Qѕ���=Y������+ףsX�1��ug0�쵿�����i�[=�n=��'⊰�k�Z\ш�Kl�C[s�5�A��-lSQ�œ�R��n�5{^:͈��.)���;;�_��������6�)Dt����_دҟ�_�&!�ot+;���p�rU��Xc�<�:_Qh���5���+Iw
氨����4���aʍ|"~�Ϊ����A�(D���͟W�NFN�nA��������&���`T�p&NC�����&���C��8(��=
��%O*�#��C��z�r
6�s{iA�O��LƓ0sT��/'�H�Ȗ��?�����V�y��Ai��
{�Ym��`�Bi�f� *Rij,�O1(RB������2aA��
�����:��V�r��g��wh%g#kr��^P?wN��ƶm):)��V�B��$il��$qu�.Rő���]x�����Q-jd�ߋi�ZG2�r���Zd��a��~?���9�ď����]�M�`Ԝ�w��:|3�7`�I�z�	5��2���l	�R�w�.*@��&&4����$e��ؽ�3ͯ*`��E��J/�{�<���M칾�b�Q�@W��)�zl�����=Ȍ���#X�cLӟ�v��s6��E�bl'A�b�I󽣬�j������=8_�ؔ>�sv���6� z�#W�l��3{���#�=T�5ƚo��l��d4xq���RƝ*�+���:(�.N
�Tv���J%�=�S�,�o�%U���_HW�-��R2(�"~���'�^��L�Y�� �A.3�	�#��g�r�^["����w��
��;�[^s��d���='�Bb�61*%���S�WY�9}��\�)�x�<�S@I.�-���a�ɹ�����ܒ��=iB��Ю ��^L��+[���A�JcXN\>��	�{�(aV��y\�"s�6��F�XS�?w�ܦ��F�|j����F�F��hk�����U2���s�����
b1aڏ�dYg�������� ��.a�=��lG ѠM�i�q�g)��DA�%r��G��4`��*���Ap�򈋝�v����%E���%���9����l��!���B�Ֆ{ �w4�4�#Q�m�w��7���8���PCS'H
���D��" ��e�܉����w�j�a�m��A��U�)��3��A e7@�$Hy��P�פ������sUl�m�=U�i ����>"Y�h�������� �§��}W9�MR�C��_�k��Ҳ��(l��+�ۥן�ψh�ަxZr��J�}`9�[�Vgx��&�U��5D�CG�j�n���>��\��j�|\�i��cm�מ�T�(�T�/!�����*�YL��b�]���c�l:����ދ�MlQ1��k�B��N��0zȹM�`�'��9!���a[�'
������,/������mKY�Ȝ�m
��z.c�Cp5`f�n�*���wOl2����s�d�,����("�ؗ(�[D�ҝ�ԜI�SBx����6bM<=�Y����酀�]�6)D�t���hм��>�����*�&�1� �M6���m�q���Ú�~剝�Ď[��rx�q���`��IO.�Q��Dу����b�!�]e�d��ˠ�
�?4���z�#����v���e��T���;��sb8VL��g�)�8��{T�l������*3��l0�+�.�}bشCryR;�>x��e�F�C���
4.�(]�vņ���߻��2��r�]ѻ�J�b�K�`H@�ʓ����6s�����bڦ�tp�_z��?^
Bj$�*_p

fe����`q���0��,�G�&1@=J���!��Z�/�~^�И�� s��W�5�U�^����!J���9Ʊ⇉�P]V�H�|�^|���ƈ�\J�B�|K�ǐ[���P�S\/�}?���	p6�468 ����W�s!�O���䎛���S雍�]1^� s�Lv�x�X\�r$��N5������}�QB�m$x� L�;��jg^���d=��*_v~����ʟ�����F�8�0B)z�_�Ҭ�E��3_��Kmjb������9p���t?��&f$&��	ǻSu����<�ÌǛ�'�NCS���>�64@^}?�:�w�o�W�B/j%&��{�S��ވ,�"9��}���}�1gۣt��J������&�;��s$Z�+���!N���-Eg%�<0pl��6|�`ȑ��w��l!��������>�c|v���	0.�@R�Ahu*�D� �8��Ap��2��V�_�Ǹ>��%eE��!�1��ݫ�	Z�&�l�*��,�U�%��-�r��)���M�פ*�^�1x�@��;��a�+�V[����gi4��O�xs��O��,q���C�Cm"^��%�eȊ�AM`#��~�[�2�A���
_�r\=��G�����?vؐXQ�����g�9�8N�(�����:�4��������:��[�:���{��.���p�w!{�DXt�w.6jN$y2��Ǡ��v��Az]4�i4jV�<@��@��+Y��k�q6j��~��QԸ�y�j�(���A�2-M�`����I����,S�[|T������Z��R����-e��mp�@��=:��, �ɊA����8�u�C�F�|$��n�p�����,R2����w������:�{݇<����5?g�.09U'�>����QeT�r�tNG���C }��T �Nd��$����Px^I�XA16,x���HBh2S_�[-i#�/�o3q���i.��{R�� 6+�k2~�
�V�o+����֪��R�P�|[ɾ����4LZ8�9ԡe7��C�d���pZ"�E��-��'��1a�ǩ`���7��"KQ��𸑗��W�0m�A�2�����D���Z��/<y�������[�J�W���IA��(2���\���t�uV�&d�J	ҜL�>b0���-&���hB�,���n*Ӂ���ᚘ��q~�>Ӳ ��"N���ش�t:���P7%�N8����W�W�%0@���	?g����Qj�^��3<M�_�M�D��
�Bt���娇��"T?�
���G���������&��;L�+1/eq�������l-"�j��+~�E��$0R��F�I�a�x��y�sJ�1"�K�=�v��q�hGo>u'�a�������-�=I���� �����=��^_�®D����[nP�������Y������M��l����ePV�ډ�����S �`��3�a`U�����������5���[Mn����j�o;�Z&�W�oZ���2���#��hܚ�,���C g�QdWe�����є�g˝�JP0r�D��<����ḅ,�_W�_�،s{0	f�kƢV��EȔ�� ���ùc���J�WۓX^�W+B�}j��m���k.�K�h���Hc����}�k��~{	�Z�0%Dq����@]ro��Y�rgiM��kv�d�u���fB)���y���F��ð�I)�nu��k�j�a%���k����U\�s��W�I&Gq����̟N�Õ��P��������KD�P2��^����`�&�G�5��a���ߤ��2��K#���]�����h�~{Sn�B��tX�8؟h�ܳ����G�+O��ҝc�d��xt8���L�<+�I������8�$���lS^����H����e��'qax�TPj�J�y��4c�9�	��
~Z�|��2G�������d8����L~j���|��	�`q�ұ���0ك�Wr�+J1}9�i���'ZE�Rp��5hbd � ��{?I�'O:�Ej<�n*��� j���x�����݀\����Qx7)�VE�wD��~�Jb�ؖ�l"��J'��c�%��(o��1�� �A���'��^��B8<`�%�����Yդ�t:�u�ŭ[CyDG��"�b�tr�i�����_�-� �Sm'E%���Ć-�N\K�T�e�#��tz��U�;S���b$)��bF*k�q�w;�.1#Gq������O�k����-��1?R2$;�h"��Ĉa�Jlj���"���_$qF�ŗD���u���L�L���1������D����NN�at�.�ۭ ���2�)�f<ah�l�HF��nz��7�)2��(n�"-�Y��K9���z)Nϣ?�f�(���Z7Ͱ�},W`Ę��q&4}�a��(
W``�Vh���j���]��*D�DGL�p93c�4
;��>��?Ig�\�KZfU:��L�1�+�c��	�H��"��$�QkђI�
��W�W���͜c�MYb��%r��#\�8n�3#�E
4 }A��7"
�޲r�v��y[N���&7fS,6=$(Z���[�G3ܽ�)/cG�E-cc,�"wtʾ�ܡ@�L��� c��]�b�hG����ߌv�Q���܉�?���T��O��*�^�B����_b�x1�Ij�J"�D��L����`�Rm��� � <���(�@��TB�j�%�YQ�Aj!�fK,E`\�k�Ռ���@������ǫ����W�����K����< Ń��/.x��ܫ�$��u_eW�e��(� ��C���R�N�R b.-U�-��������_��
��6�����ȟ0���Q�Tܯ< ǎ��Ż[d�좫f�p����M��B�f��W�?�<o�B��u���Q<��0�ʥ���.���yeS�[����g����'-���q��1o�:ї����1$�4+�a��$|X���z
�����VIh���^�͍o�0B��mQ��j�RW�ǰY<��6�F#Y~9��vc*��>6�aT.���đ_]�S&�l0�:@�`��Gq\�Zu��6�CS0�!�1�b�J�s���S!�������;�>�a�Ӑ������������x5�%�z���/B�����4ͤ��VTn�_U@"��L�Z��13�?a$D~`�WN:b/�QQj(;c�wnY#:*0��e�iXE;���ʫO݀k�wT�/�������<�S����X{,^w߼������	�������{��62�l�u�%=�(@�,�i�#��)����ső��~k7��_2R�|<J��Q��ۗ�9�v�mܛ��/ ��L;*����5�ԳmV���d[�~T��JS��Gg����%q�h����#�+Ä�rc�*��	X���̣XLK{ m���s��5��Ā����`����X��x��*4 ��c/�dP�J���l	���r[.��^ZY�E�g���B&�a�QZ����b�x�0v�Rz�U�³/f�	���v��Le�rމ7�(s��H/��ܯ��m��bt��Z��3J67�bi�N�ɗ@|��m�g'��]���%I��������"`gluSm��߽�Y+�a��>�I�y�;V��z{� ��b�~G;
��R4v
hG�bSF�U�V��e��lɮ+���$�@�������DZ���1��	T�~���+w��[sr�,�u�P�'�7j)��cl2���~���<1�����\�m�ʐB��~���2X�G�	_���e�"Q/C�L�R!24YPg<�Y5�f<U���G(g?� �C�ݥ[��)!Rߠ���fph�"j N7�ձ̱O�����&Jr��2�p\ؙ�'l��3\�%K��Q�*ʜ�ўJ9_�d�Նz�(��*�U�t�g�M�m����	��E��{@_�A�zw���r[���/��1�g���} ��F����"0��Hj""$ɮ��z,��|���f$��wv1��r����� �8^���~L��Hv떱�V9�'��n�(p���݌�=��"�������'7�I�Y)�
��u���s����۟N]9�"��J�,�Y����@�︁Uȿ� Ig�q���]��U��ǘ4$���4q��C7��°����HN�"�G�]���C0�'�c��T�t"������Y�5��� �}�)��5���⇻<6�a�n��o �
f����xHȇj(cN}������󟦨�.4y�^�簰d�#l�!�ݨ���ML���V4��	؅�����%L^�_�z�<M��L�,�~$�N���	�����/v#v�>cck��}m�ZB)�|�1,]`�[0k��!@sA�
i(h���$����W�dCxO��Fd�D��Q}G���K1����@7�\�@������A�Y�t:�'P���z�Di�;ǋN3��#E��z�T@+����y���=`7N������n��ÔJ�2v �<;gG��'�!�W���4k%
l[vH�]�	��L�%���3�>x��k\��|��|TC(��/yD;��nt�	�G������
��5�K��QވA�����@:!⺉��oMLj{��3Ҫ͎����<N�@o�4om����ܢ>��^Q)(�n}�3P>�>H�h`�Mqc��0���b��3i�W�����h�,��+�++�����"�>p{��Y�(d�P�4F����A9��A�����&kz�h��H)j�"sg��ivj:�����i-�ĵ�#NJ`�Or�b�Ђ%U��@��_1�h �w�&��������!�l֊�:�$f$�;����G�k�k����:���9e`��^��q#����m���&�8�y�*:k��֧�,:��_�D��0�I�X�6�T3����O�c�
S%�L���3�<]N5��t�>����ͺ�wO��"ׯJ&A���֚z��k��B[����T5��ÐY�?��8�D?VX�OT]��SS�����&�&=��W�o�s���ؚ��8�*���a����׿���6<^��M��� �䙨���֡.X�'�,����M�\>�A���x��P���eY��*��y�A*DBX�F�0?]���C�3YL ���Q�\k���61s?�� B�R{��s�#��6~"����߰�D��V`�j5 T]�=4���N6��ɨb��6���_a��@
 ���K�����u�iϡ+�tg~b�b!�L�62|�&
�4lwLY���D	�hEC��e/�����7����/���J6��,�*V^����
!���[��F~�%`�+���>�݇�K��'���8���V#�W��.��՗4<P�H�����A��>�87䲱��l�V������]�R� ��x�;t�B<*v@B˃�Ъj[v]Q��B?xD�\��o�i��4����O������2���c"R�v�	�͓�J*6��ppY���X����7���12��B!��E���)Sd,���'!l]�K���"�f�2�B?�����߃- �������)w����cˢ_���>�/��-@�ǳ$�0����!t�3���RZ�s�q��V{L���7䭖Qt%��U�@�(Ҍb�0\�$3HA�� &�=�wb�AE�z��rw���R�ҟ;i�F贴 �s�iu4��[4����'�1qӷ}�N��G&���D O7��hD�:Q$\��鯕�f���g�ƕ/�t1AϭlQ-��]��Fv��a����9s�1*���Հ�^I� nх�߄5<�	�0 H,_,��W��F�I�Q��1Yac�P4�����N߰�x��9�(<Fy�W�VW�S���#>@zA�6A�3Ķ6�z^3=��Sz$c!mR$�{ߏ�i	x��� �`X����1x���v�[4b���U<B`Y7�ؗ�6������|�^�k��"0��^�-���A���fh�Iķ%�Ƒ�ot��3��`G�����;��aZ	[�t��[�R-�����`3�<�Q�g)��mFjϫ�M�x#��U�nZj&��5I�i��o؟���3I1�7�(���Ds`��@C0n��d�:s�P{�U]��^=�"k�k-�' ԣ#Co$R�ػ�OD�c�\|�?hX�%��B��X��	7 [�]�K��IM�į~���fM���a�;�1���~W5(�J�~���k���v�ր�L*�G]U�=�C5�EK�5Ao�D�x|+c{z������X��1�8,��62���ɫ���J.1C�p`����tv��\��t�T9
v�Y���V0��e�;ކ�b�ϛH��8.�F��HS�ʭQX�O��̖�T~�H�Hŗ��I_̤�ZAVq����G	6�$f9�&O���^�dُ��-xH�ʯ�TZ7e�|
褵��Mp,�D��9,��J
���_(�y̕G
�N���A���K<�̇fjSq֞���μXbJ���f��O_i*G�U����QGy2?�ຏ�H�ͽO
*v�<�=�z��k��~a��ዌ�J$���T��<�Z>��Wk���?���TB���2`�y5\N#�pJ�Z��t������ԇ��[9���p8�Կ�N���tr��m>�ӧ�a�yN���
�>��Y�6�&����_���X����Y�ާ�R^ik{X@�+��&E�bנ]�H��yd\���2�kv�8\���r@
�ˑ�X��b��\�&BƂ(����[d���P)K�L��Q��s4(�2x��*æxK�|(�R�
���ҥ'���wYR hm1�Ï��c׊W���O\B�i�]�A'���/ U�I�=tc�=�=�Ͷ���*�����\���lէ(�� cB�|p9#�_�l��n�$W�Z�n�\����0����wcۗT�#�^�*M{'�q�qO�N�"�0�{c!��]g�����vO�����'����i
0nyK1J��t���tNv	tz]l����A�i��2<9:O9&~Yw�m@�Ï��'�����>(�5��vRP��&j��j=�0�Zn���3����I��[�L�w�d1��}	 ����d�#&�)y#W3�h�
�*���K�H#zKH�Ev#�F��}�6��E�%Z6O��.C����D�CS�yǺF�@za�>����;�����K+'>[E��!�\qnG	�q���k��2NtnE��4����5=��Ră3?s(�/h�j��B��*��EAT�|�R����+��?��{�Z;���g��'2"SQ/+L�ų��=�
g�rl�En�Ua&ft�v�wI�T���y����`����m�%<� ��4�'��Z�N!��~m�Kp[[�<������ r�M��L�����1I���]j_A =�h�T���n��O�H�U1T�_�I���2��L3�t~�t%��������%7�%�r�'E`�@o���:��z����M�h���mI�ȢY3�Y�vD��0���!�R	u)���~.���T��H��MAL6��Q���õ����K��U�p)S��p|���(�/@�^������bEQ���bw�[^���0p{�β.C��@r�Js$s_��dN�B� �J��Jw��V8ٔ���E,��h��'_�a��&�a���b��8�n���ibL�Z�މ�y~C����Q!�3�� ��;:�	^��2�������dN�ʸi���=!����;�,����iT�J�R����R����<`S���D�����j@�sd��l�Lr����z��?,Ò�,�_d1L�iͻ\���1αy��G����ڀ+��]��lıx�-LP~��Op1��U
r��˒$ �H�����ԕ�8el+�a���2���G(e��;���5�r���\����_�J*�<9��K�&��V�j�M��������O��k�oP�`'}�ı�T�����C����]��haq�����7(W'H�LV��n�Y����3��8~Q���P{�S�P~*i�`)gRP��w�-�M��,���I-�:J��X��YugE5�����-�Ο�!$ b������i1�"�eߨ/p�3r&o����V�k���K�-5��pCp�N!춗i�w�-pf�y��O��F)�)Q����fjk��r���}����k��{VĪ-;cMnK-g#O���~k�c���d�1	�����~���3rm�#�:�������8,��_�a-����d�J��&p�V�pDP<2Ge��FD��Ү�K��⾱a�Y��@E��Y��\�B3T�ڣ[��ފ���vz�|Г6z��k!���࠺%��J=�����������# ���veµ,,�`9��F~�u����p +��5�(�(0�Fz�%é���':	3�'5�6���_V����ńRv���\�l�ئ?� �(��A?���Կ�����]}��KF����Ȱ��]m(B��e�����?����W���N�����;x���~4��m��ĭ��($�<����U���DH1=e�#�m��'��-E��#/���E��k�)�NS�mt�����\\�#����k�#���=��7	�gI;o�:�3�/+���J_��}���a�f8�:�k��l��(5y�J��7�E�Ԃ'������AKm�?��؀S�&2t\�F�����>��3v��0�G����O<�o�{x�WAu0�]�l����|czH+�� �A�[Σ�{�8�Y/���H����nG���Ԫ_�i$�>��4�n����ۣ�	S'��jf�%�W�ʾJK���q��L�E�H9�~o���H��P?��Z�L��ft^�pn�<�5#J��{~�wSX����>�V�{҉��̔6�9`K�4{�ʷF�BXb��R�8�Jd�]_	��(uh�k;i�h���d-�P�{x�#�Bpk���}^[�G�]���#>�Y���v_������Ly>�a���i��rod;��D�*T�3���>w-�@2H����8�@�?����� ?|hN��vS�d���W,H����w�JA�_s$��+۵���dۘ����ZW�T�]y�U�5ݬ(M���氵��V�i��׌6�xv��c�Xtr��K��|���i��D^nmj"���i��kT* ��j�	�ձٛ]���B\��VnӐ�\�
��Ek�T^; ��)\�f��:T�=���}����q"����"_%�S���~��1��D�ҥG�kb��!�� u���0
2V�d�Y�k?y"���uIM��r���'��A2Eإ�M.Jfy���Y'��B�frZN�Ͱq+�r?$�{/��5��*2\�ߒ$�A����`�&��;e�]'kzO�eu �^+	���D��9�g��|q�s��~��5#Ƿ_���g8��A�i����%�-X`�6W[��t_F�Qbϧc�k������_w�~t�Q|���A�i�Z\]Z�l}�$=bW����&��1K��M)�/Sn!�>lȳ\�~@;|l}9Li�c�& �)u�?D�ũ�N�t�y%���2G"�K���.�����I/	�b�9+%w�F���t����ޞj��Aw# �/��f�w"�%�4�����{b��g	��I� =(�r()���DGPQ+1�4��߻
��]@^~p(����o�v��9u���s}o�G��RZ���X�堥���<N��_]tAi>Dl����S�l�ݽ�\�2��լ�\��D�֟-k �Z�z��-K"aa�F�)��,�p�j��I��q�d���s7�r���;���?h��ʃf\66���䵡��pʶ�@�6�(z����0�7OApN������{�|v�OO����=�b�p(b[g��Ua��^�������ؖ�PT���ӡAE�� ���1�����Qíp���,��`��Ktȝ�A[���O5v���??:��9��a��[��t�Md�r�O3��g�ѩhE]/����X����*��[��+kT@ZB뼣\���LXAo��W<zY��#���V��^f�|��;�8r"�K������z�͞�q���=�0��� �d�"h�M�LDn�,>�厓6�̶Kk[�bt���sޔ������z6���Y�1����+Ċv����ؘ2�,�GM�,DH#g��&�O�#�Ԓ%6���>��ěÝi�%�,�f���/=+�a�wdGH�HC�C��RU�����)\�ɯ'k�X�=�[j5�^�����fw^��X�Uϰ�@`U"g�������N��@}��M�kG�/�B:�BoY�S]K��k��}
v J2d��4����IU��E�	�ʯ��Ui&�	���c��(Ī3KIѽڳ������I�p�Z�B���nt�o:�8��f�i΢A�,+���Pa0�h�l3�1�m\��)��:ڟX!���M�,+�b(�C���W�F��a��ً@��qJ��l��'���f6*�(�,->w��q���G��rN�N�����Ȩ�i�O���~P���©��C����0�Uh�dh`Q4�mjO-)�Y�R[gy��`߹��n!��m��5oO=(�2J�ǙN�*K���ڪN�R�����
K��b����N~���H����������sk��N]��֧1�׿��g�cw�nD�B{^G����fa�0d�[_�Ny���M 
�0ԆR4)$��^�}ױˍ00��e�D.qK� _���*�7ͯg���Z�+�_��b+��q�����T%?!z*&�׷�}�$s\cl�6�s�j��QF�����eS
8�J醈����Y�:�Z>�ă�b��&R&����5��)QK��;9�&��)�(*�-�b?��+nC�~d�:H�O�0�����nGD����7 �;�D%���)z��c:���<���@̕h7�j�~��m��Qxa�h�0�Zt��|0�f:=�1 ��֠���{hd=b)|������Y��e.�g����eW���g1E+6!���{
R'Dْ�p^^6��	�
�,08(8�n�_� -~w�!p�̂ݶ��9��(N>��:�`(�21|�U3�����$� /g�tmb�%ANdH�e����/�6pH�z�7F�ǋ;8�Vmћ�Xb����P!	�\(�us��,خ�Y��T��ћLC��տ����5*#��cx�x�7g�=��v�M1�KdwR�x���e�k[ϧut��;"��qa�.!~k�F�=T�Q�h^	8`[ch��ϛ�>�t����������;N������,�À�]{�Q��O]��4�w�!�� �2��
�1����a)�]�x���V}��ŋ���gNYn��*7���zm��BO���w�� ���θ��]�ȽJl��%�΁O�G!zxO�ȴ-�B��hN��>������b��3�~
Q��{Ol ����+ߜ�qK���L��<ɢ��c�_b(KDy���δ1���^ٙMeC���jJ�:��~ kX΂�|'�������<���bG��b�.]{1<��6�f�=b�g��?��}�w�g6��a����/��zV�`�r�7.�$x$A�NMZ77
������A���������, ē��3H۔�υ�ԇv1�H������KP�G�����2�.-���f}�1���#7P�L@�����������4>>���V��*��?�4�.�.��%�r'���g�R���s���G�X���е�,�)�8*REo3�����f�Yf,b^�Ǔ9)�����^�׳����HI�� �j5�"��w"�<[�n"oq4����5[�V�NC!T.'ѷ4yo�GW�G� ��o�F�.J.�y5@bq�������-�/^E�*�t�t��_<@v��I&�@�s��qV~��e�3��>^!X:�:8I������j���◊��:�9U��h"w�h o�9�@%N�39O���8���W��8P�.�Fr=bJ	�Q�jMj���ӁK!ϭ�	��G�$5�� �Ќ3،F���a]����/�l��YIm']��v����������������,G59�1��j7�y��t6�/�y//�>��w�;��fwid�flV�qr�֛ۄ)5;��}ܹ5h�T���a^��\`�"�n��r09�eC��M���FG���k�l�&���0_v�9!w���Ԝ��|Զ�� ~F7���
v���!۝il�\f�����*��Ǽ�H/�ap=q�7:��r����� �*�4�g/Vh@�>�RAX>��>{g�J7�#(�ߪE^�*0'��[��+����߳,\K.riK|����T]43�2���&����.��!�qΗm(��z�RA�A�6�|c?D+u��6��u!���5���d�f:`äta<�� H�5��3��F;�G��yܵ�j�6;��S!��t��tE��b��|��H�\]%��k��O�b�V	�Z�e���swO;����>��C@��]N��"J�kr��kA�J�/�)03�¡�9%� �F�:kA5�k!�*`q�n�f%���J��s��9:p{�ou�\�v?��h��#h
��j�gߖ��bו���\��+� �f�׮����#t�h�yQ���لp9�F`�<���9�+���[%ⱂF!��[���i��?a"��[-�SP��nke�qd�#;�],��C>̚p4fsoh�fNr#��p<Ҿ}�k�m0yN�;�'�����7��`H����xy߽a�=^��n7U{݆��#��T�^�qMW-ح�@��!�������#��J�"��K���t� �/xz՚�����W�p�+(E�N4M���rޣ5��KA��O��E�ޯ�x�:���z'��0d�#�-�͖��k�✺{;R�#�퀙B�o]͏�&��>�(���F
]g�B�UY-��sB�!�+��h&lC���s��1�Je�V%e�:}-}��z��PY:ܛ���T�av�׉i6W�挹�=8t�Jb�Z݊ݡd�a,y$ �tS�R4��/��6�#	,���p�T�i��HpD���'��_���MU�U%u=��j�u�	�����4ۺ�G�u7�c���X5�)��L���S��)6Q9��M/t�"y'Ʈ��'*��J�!����Q!��hq�uV#���4	�5r���	�5�Ǳ�3���АM�i��!�?�y͐+Mx�P�Q=H�<��[��*�&a�1a+8��}���J���!k�:]U8����W��gآ���@S���y��ه<��\\Q�$6�	z�����0���E�G���Tt��Iny��'���~Xh��\uc��Fs�$m�W���֦3V��UG�jזk��Y�G�'`o�P�4�Q�yG��omC$zS|Ai﫴Y㐡�K�zod�W�����l��U���oA	Tg� �6��[������j��N�����-�#�k�C
	��#���<�S�8X�X����A�J�h��tQ`�(�>����kT���]�p,-_��]j+���D��������+��-�t�	?-.H8���]��}ߚè���<3�O���qRc.� Uk=**r�
宾y��'���d��x|����'/!~7�& �6��g\�Ǫv��{!�^�����3A� ,��8��ށ����]��yD8n��<�����x�5"�@�sMC5z��kCϓ���㜫E\șFP��݉���K�;���������x������f�Y(�;�w�W|������E�6l}��~o&F� ^�@בkץ�6�z��y������q��{��mː;5�a�9���Q-�����y3��q@�Sӓ������uD>�ֆ ��F$�2�=����GG3�5L�˷=`q(L��JϺl��Ė��e��zF�L	v�L���g��7s)Um��$�r���t�2����on��cUlXc���xk�L�bD��?Wڂ�h���_.����b ��z�����q\0o��Om�/m�%X��1D��h��d�����"������n�!NvL��ؙ
��0Z�6S��y#�|�����(H)��u�H��L~��>� �h32}$b71r������|��f�ߘ��>n<�����{�Nk�v���n�Y���!�s�p��~25�s��6��*��� �{WUT��0@�9]�Q�������fO�Kݨ��{���T����^?Ab[Se+y8�O6��/ӽI���6	�k���_����~�{����������Z9�
��	!(Y�h١��%���1*^��~\�ͷ�sAq�o����<l;#"Z�D���X�#�H��s�:�^�'�������6M�@�蝯<��m<\�ry��t
�F�&
��<���P�q��A���
$c.�WOV���.k�Q#��GIu���ߢ�)�+��JB���qhd8��.$ʱNf�I���U	������)2��ͭ���%��t��k8p9מ��Y���@�����qK�=�v���[�5z��h��N���V��.u��A*�ۯG��0�D%"���&�����H��Ժ�����<�4��f�''��H�C�A�	����J�}`!�%�@�)�ܪ ��u$`Pk�(O0oh:���0��9��n����#���#h"\g��EO@�Ge�Vo�����!��ǫȋ�C��^m<�s�6}2���k�H����N}:�E��-��?�J�KE7�4-I��k�?����Q:��*d��z���p̡���-@��$17OP���O/���`g���/��k:��@��r�>:�ʮ�`�����4��Џ]&WB���y«�Q�Փ�13�� "�����I�<.ŭr���P_���W��_�/�5ɵ���4i�Z��Q"�����N���m �qL"ڥ��]<ڣ��gǘ���>*����6^����^�@�i��/��k��yex���<�c>�>Ed߆�����mc)鹾���K<���:ш��a�+�h��������q�����&E�:/}P�ì���?̈́�����kH���۱����@j�)���4<XiON��)��5�v��8��Us�T�:~�¢hb�\�sb�Ab�����旦C3�=��|���$wdnK��A%P&��������gIT��ڼ���e����ʢs̀�suZP1�J��H�;0� {�s$�cH���x�ެ/L��
/�(�=�Û$~�9���+`�%��M<&�֐���3�~�B����<�j	�6@��Gǆ�)<r�a�m>D��E�Lx6Z��ty\V��i�?YP1�u����-7wN����	���[����LD��;9)]��X��+����00��m����/+B�ǘ���8e�ɉz=6��ܒJ�.p��$�Gu��aB>��Y�{��]p׉�IީX���ז��]@�ZOr3e��
O��\Z
*�D�[�����<H�v2���a}�Hz��M��f�)dT��C,X� ���a�^�|a�A'�ݜ*,;���,����H�8�9o\����*�����U׸������/����2I����(nɻ� �����Ֆ5�w&��I��}��A���*��������aJg2u`��Cl��:%���'���G�)A� 2�ODePҟ�<��5���uؐ���ؾ*���'B'���jz�'-�8zNd,���}@mV�Vh��F�/���>��Dn�ˬ�L�A��"�*�~kG��i'��<�O��LG�F��j���Vmu����G�3t�*�t(����D����M`�x\�� '���ٶ�i�P�N 6>!+��1/�R[�Xz���W,��ϙo�m2ڈ$��Y�<�Ӣ�R�+7f0���#W>�uB�v�[W�N�@R�0w�c�/B*f������,�Q��e3��C�w@V:|��6�=�����:w1�*�I������o��E/��W�;��2�������WΔxH�.$E��ސ�R,B,�(��哏���i�������ي饆M��z�R]��kJ.�HS�'GA���)�g�:
��B)���s���s#J5O1�"����\�\%��_�H��� G����v�Ҝ,tfGg�W�!�Ҍ	���}	q�h]� X�M����ϔ:G�����+Bi��w ~y�/�i��
T]���Զ��B���zR�7�P�1�l�Uаx.�@"H�wi�}�� d[�֞�-T�M3���n[T�����h̑�1���r�rfבB���t��=i�~n�P@�N��Yb?��R?�Ʊ�n�hZ�w�fe^���RmR��a�-�N#`]�vu����횒vQsm���A�������Z/>a���{��j�o���^]MR��b���c%r�2GD���"Z2ER�!�bxS��zK�n���Q�@��3��[�٠�K��f{�`�����=��?�^(v�n�.1y�d��ɒz�D<�Aٯ���ܜN�4-���̝yR^��
��4��k<�Y���.c$)7���;�Uy|LF�������~<�6����E�&R<��V�)�j�|�i�OB؃�[}
�W@P���MIK�cbr�v���N��.O-π���r�ί?���]���m#(i$`�ĳ7��'�=� � �3ZH�"n�6S	�ￃ�,����\]$�@`c""��B}x�G�$�e�i�/��h��m�Ge$/*���[g���T�[�����6���h8n�C%�|����Eȕ�;�����5\�M���%%qϣ��6O�>*��!mS���s]������9/�����v���oJF"�j��J�>VdA��2��,C ��������f�W$U
VI(���']��t�/X���p�{�O(?�S��5T��"�NPi�xfBn��!${����j�������B�oz�v����&u����k^�� n_(W̃����Z�5dB|���M�y�g����]Pmc�@d�A�C^��'��݋S�o���h2O�Xq��~e;�`5d�)N6�k���,���e�<�Y�#e֭��#)W6�"�MStѐ��t�M��lq���O���2ڊ;@u��P@��t�6I�=�Z
D1ֽh���OZ�r��Ñ Of��eRx6�B���gV�j�;x��\�)�����<�9߲�Umͅ���,U���	c$t��,��5���J�l�S�怐�R��bH��d̳A�8U���p�p�cXZv�;���Ȼg�Ouh��y���Br��b٘��/.�������;��d�b)��jF�2BZ�C����`��WnL ��Z#['\-�]�E��-�5>$��2�N����%�e���Och�9�7��!aD�Nc��q�"���@e���N�BUn�s�����Gk�w���Ux���p�efP_-�3��{�C�c��H� �6Sh%����kD1R��X,�� V.�6\�j��t�����	��"��T�yxx�zN���Xw�K�5��)��:R#�6x��]jp�c2������r�S~�Y���.�\<��9�7080v 'dq�T��h�:-	T�훎����㄂�y�]���n�U��+�1!!����&��劢��q�+��n���tz+ѹ�ڔzw��q��/*�Z�|�$�w���O����vkCM{��)0Z:!�`�Z��5��l�b�:ۙ�0Uv�}]���ޙO��d�C[�!��9�A��gCb ��rU���j�1t��b]ӊؘ������s�]�u$B�I'l�V/a!�a��,[�0R~�9qWb�+��˥�^Ni.���v��5�}���A)ר���F�?�$�;.<���g��dbV3s�v9�jT��.k6UHP�a�Ď�{�	���p��F}���R�*Zt�dL���f�uo��U�K4o�{z�g�����"�&* j�\�.y�h�_E}M�-�`��۰�$�쮬�T�/��@���"�I��j�
���	�I�7T|�Xc��<�`�X]^E���#l�eq�{�-�H�#���`r�C^ad�������?Ψ<yߎ�����^���h@��V􁼋���jR�f��tǏõ�m*\0��D�c��������5��zs{�hE<��rz6��eC1�@�Ϣe�.ZP������eV8`5'n��������)S�Z֕�
񨑄���o�C]V�,�Um2�2��F�D�'�Ns��)�C�*zK\�R7��῞by�*�z	�����E����K��t(d�.E�pon`�Ey��~�@(7�9�&���#\��Ҋ�#@���s��N�a����[�C�n0���Jʅ���
܋}I6PX$�js����	b"(��y���x[^z6&A{Ǣs)<*w�ħ��tg�3r}�Li(�u9�I�T��x���$���������Z(� ��`�ǝ��Cx"ˣ,qǖ���W��tyD�`IG�M%#�j�e<+}�Y�n��w��h��8Dv��[p��m`�r]G����6�)��ӧ��B@��/
w��M��>0��Wp�`�g�����b���H!��Z�ܩDT"��,���9 5�����SS~&�%O撧���z&��	A���_�'�e��ɳ�zD
��j�.^?f���9=E�����$���� J� ���KJ"K[Z���[�$�Ȇ��W¤v5�#�,�p�@����%����L<��u���e����P#1�'�q�(A��1j��-��1��Q"<+Cg&8�����������gi���Rm�b��0���M�i7���5T��C���Y��G�\*��sNy�4�7�F hp�1B�.*c*�D�QI�2��˥��G^ݳ��r�[n/�M�j1|�I���R����D��#�w@��`��@Z#��j�� `y6*�������6��s0�X�Ͳ�g3d�̜��
+f]��mg>Ei�щ;P""�-��~͉���r[�󩝨,�1�6MR'0����JRN�!��%��`��8����Zۯw����4WS�>��;']�^+�����x�vzɉ3�2RS��%�<
4��{�;l�g�V�9�$��\�+�6�����B>w���I΂���g�Znz 3|�݅�L�{HݣHl���7k��/e�e{!'Y��Q�[����I||�.��  ��S����c�����x~��aכ+��Q����!�^�1h�4��ɠ��}l���v8��eb��tz�sX�v}ߗfY��pM�KJ=bj���}��	��u���nns*<u4Z)6���PaF�/ �s�oN��A��LVzC��V!�� ��Wق���Y�t	l�K!�o��=5O��7���K���i_U�b�P-r��a�x���여��*��~!K, ��!��8�����
��P\��[K�i%<A"�Rk�Zɣi�J���2Mպ�p�o�t�q����4Ӊ�^�����-f�h�����1���_�d���stF��(b)Q'���PS�zRD���j�9#{&>f&��E�G<\ZD��v'V��>���ʬg,E���R+Ǌ�?�O*�����n��%��fYM�R���Uj1F��b�TB��E��F��T��,j��V��x��B�h/�%T�-_��+�%�}ꇁ�M�5|A-m��x3���?7?�+T�=�������� ^a���B��*:;�Bo[�i:E5|�����H~$�g��PJ� �1��x�)�ӷ�݆!I��փ[���Ջ)cgC���d��ʽ���{�CZV�$��.�9V{ƒN^��, ��Y��r�w�  � �6���q����<0%�|��/[��Hi/����26럠�7�hv�yd�=��Y�ox){8��i�>+rҼ�f+��7�@V�y��݂�a���X�WP�ep�:)�egFɽ[����'�ۿ�m��R�q�����1��o���/�I�w�nU��wr��#Ak
9���b�|-��ci�	�hM�)B��G����4��`B�����sք_�G��5]���]^������E~����L�uBQ��̛̰�*vam*)�U �w+��uID�3��`R�<�����ԝ�?
,� ��!Ɍk�v�1<��>W� �&0�L���iW�5`�<@o��Y�#���9rZ䆈�.���J'��!�����]�~��i��-��H<$�be�X:L4�Ģ��[�!�++��s[fRtY Y�	��o��o]���:��>��q�,��!u�۟w�O6�5�C��xb����b[��54�E��������ˁ&�4?'�����-o�"sCu�m��B2��*�;8S��V�G�P��'�Kk�Ó������s��`\�ְ{�f`s����_�ȟ��PBM6���#��O����Q6�9.UPd������w�f�l��I�]F ���o��-kc��%�f)�4�y���d�g����n ���I�)��`��޳.���)�f��GX��P����1r��e�2�4�~�,�y0!ƽ:�Ʉ���q�_x���l�).���|˲?~�bN�� ����9�f[7n�Lf��7<�"������y0u����<t<<��9 �Y��uW���R��-��Rsn_R����n���|0�k�2,P��"��EyU�m�3:ƈ��j���7��YY��|eZ#?�k��$��`�O׹�r�v�⤾p��y�h:5"-Uk�
N_~�藸6P?�Gڲ�ѳe�Syz�z�X�����,w��)��s~�8Wy_a]
QI�b�љȤ���Ft��󨖹�ym_��PIa��A!#=�	�̈p���C�v
r�9!8SB=��Xי�	�݁�L�5�@o��E2 ����}.�,��w�Tf��U�)J�a��}MOt.���{ع^�2�L�+6���>��]�E�#z����@���p}#�.*
̓���a��¯�nI���E�.�_l~��ݞ��4[���:���E:��B���_�����Ľ��p���k��R�i;�33�C��c�[���f�� ��:d3R;�#���~���.���}-�蟗�ބ�ۨ�G?�^r�b�c����ђg���ysY1�fu�o�����w�&���i*i7�6WN@�e���H^�P����<��Qx 5�3V�S�r����8n���6��`U<4F�Z�e����I ߏ��!�,�&�D�Q("!���4�ؑ��I�g��*�f�rg�g�$.-`Ke�N'�%O`�8ydw���k�7,I$ܹ�-�4�m��r>�!��&����@�T��RV	Q�	�'��l{���;���D[f�(�P�h6�c��~���c_eCB������l���x4����(��%.柁�`��!*K��Ia�y}kX�I����
��e�z����q��d�4� H������[n��a���
��i7���5�q�Ng$ܫ=G�GȮT�!��ɗz���� E��ɬ����������7�q)��Ea�<��ȇf�����J����)]�+]SԎ��k F �����3'�����Ա{�i�uB�ǧZ����:KwEgӡ�bϠ�����Z��*u�tj5�Mǒ|��a��)W�U^xp��7�,�Կ��H�9V=��,��4w��4��a#�p���9P���A�X��G+F0�Y4�}d�G�:�r,���ަ��HtL8�����4���6�����k
̱~g�t���{� �eP�����D]��t���9}�Xod{�J�,�r�a��c�Ҡ�����;�OYZgw�l�=��� eA�LyWY�t�L��ow��R����Úb1CS�c̗c�\�霅�!ܕ��'Ӥi]�;f����g{��Z���(�w�j�@q^Hn>��BVˣo��@!�Û�3��_�N�s�F�/��=�D��P]�!hh<�L�n6 ��1ѷS�{h�(�pZ_�'V��P?Y�V�P���=��1��iƖc�&n�ʇ)FG5N���x4e���e��-BjM����T(�������?v��i�>C��cLF�J���]�t�;Q�ӶVj����f�Ì�aO r6T� ��շ�Z'���+�m�l^��J�3��	64z	>���(�
�=K�h��!�^�pi'��F�q�6-dw�k�L�i4�ue�%�@�~ƨ}�S��Hi�:�W6��k���."U�C^*M�^.�4�� ��q^��8��Qj�v#R��F��0Y�z���Od	�Q�wpf��@,�[S��E�%G�`/�����Q�H�k3�z~ybE��&�}b�mL؟�$c~q�]6��v�si�p�a-�z�\v-�_V�782jDuƤ�4�y�w~�%>V9���b.�K��A�u�.�AF��L�GK��@�ꊔ&�f3���h*7�휩+��'Q���|�-e������Pf���E8�#����8���e���mF���X�cy�i!��D��BD���k�Ѽ���r2X��Y�5�eD���#cv��w�Z�D��~Y)�rBĆ��)�Z�d�a�#�½2���wCTʲҽ��WȽޏ�0��|�y�K}೾Ce����P2����/���v�f8�"���&0�Iru�C���h���p���&���7��eǃ
��aR�t���A�-�4���ڃ�h�w��v����%�MϜ�Ւ���M��h�	bJ(z�5$k�p�DM*�}h6�7��@��\� �zSͥ�n!�ߛ3��u��F�Zu��E맠6!��6V�L3v���А��܆���_A� *�5�J]׼�ԧg���8�^/L�2�ߧ~����:� B��7��L��A���*?gخ��u;DN�		؋�r{�=\{�NwO��b�@��.�݇�Ȕ?�ZK�<��ri5�����Bս%��~S�O�&�0����
}�px4��F�~0�O��.��$�5A�=`�S���O��V2���QN���WK�byB���z���ɂ�Ew�gc��V��|=������	��Xs'�<���X[^� ]���v0'\�n�h�GrsgX�Y���x���87��^�et��c�����m���qD�'� 9��|,Y���/���Ѯ�������q$��-*��d�}$�~K�F�o�re�3����x���a�W|���[�1�E�M�ԧ�\�v�wΣ!�$�<�:�=���њ�I|�C���l �i�{�f	̺�t#����~�4"}���1�\D�.�$Q#o-'<Q����Z#�L��
� ��5��:���'��T���~́t�\�d�����B�`�M�"
&M��!�HEmf�g�跶Y'6�x2;��6��t�e���3����W�~J��
Z����:��{�O��<=d�c�PgN�#��L�֒H��6�5`�a�4�deY M'��n����q?��v�~ �a�n _ܬʿ���iV���g����qX��#~��	�J���k�9V��b�O����@�Y.��a(�ʉPIp��^Ķ��ѫ*�z��c�T3��=��ʾL[�C�����d4�`�S����-��,��i�J(�&?�� �qx��z�;qx˚o]_z���A�o%Ǘ[�w8Np,{�s��sQ"�F��R����9�ƣ7��יQ�����E�eq�	KH"%<qS:`R��v�px�E�#�X'VBRk����E�<,^����u2hV"s�% � Rpڗ�������"�����	�Oc+�*�%1��m$k�%P
,w�<�\�˃`ćߡ�|�����w}���s�=�zDG��E���z�%1���'��eq��9b�C�	j��1���O�^����E��� ��[�4%���k�fT���ʩ��Z6zU)�����؋h?%�:0~N�ᇸLrW��E�����ZM�����<���*�)nNz�j����(�.�D����nޑ[��d��K�`}]2�P5k�	~�Y��=l8��P_�GH�`�OG�����H��炳��|Ĕ4�o&a n?
�{T�D2�&4�2-����ʸ/=�S'�'>�,U��e��ȵh�%�p4�� �m���vB�dW��:^����GQ�����IOg��`���!�T�I( _%袻�~v�<23��J�gGJ�^`�����VʫX��ԫ-T������u��pf��[��4��NX�<e9�:�x���)�&}�.[`��w���
Caܫ�7�%�G��{��OTP^#0!�uI񟏌?z�~IM�>3�~R J��`�~o��&{ĭp{X��`$��4b�K�NRn+���CGb��_�������d�YG4H+DW\��H�܂4̽�2��)����+�'P���6˪{ G�����_Y~���L��A]�%���I�p���V5��Ɣ�GH�fe��ޔ���J��a�yJ��0�,�0~HZ�2���+���R�heנ_"
Im���� ���Pi���ǂ>�6�ңf�
�tڛd��nJ�"k|b8�����H2�y�n�������;�\ U}��g#4��m2���|錪u5b���5M�k.�w7�2�J|
Y�Ok�N��Ԧ�,V���z�5����&��D�"�̛a5�'�n����#/� ڻ�`xG=���@|���omn�ݹ�םc��qJ0�y�����M���Y��m�璼�����!ݑlܳ���ϭU�)�R%Nμ�}��=�����a��`�=�����&]3��nIW����w�������(�-��f��֫Fʚ��+Ǜ_&��LZp�l(z��((a%��^��c��<�$���j�$2w.�Hq)�T�p9%�*����y�'r��c~k�8�f3@o'l%2�rSs�[=(�ܚ̈́9�H���=�~��`ĝ�{6n(�[ia�D6V�J�Ew�8{T�C��n���B�J/	�"O�2�	(֠S@�Q"�Dt���#+�u8$�Fw��(F��*��S:#8W��u�o,g|�E���ߋ�e��W�T�2I��0�Ҽ�HYu�F��E�i�ŕ�ob����������	?��������!����t�Q0	����2���2<m*��͖����=����r
ZP�����'<KB<��i�s��kn���cm^_?�����Z���L����`���#�lu|PI�:n�-_����si'�^.����Yj�b]:/#q{���HC�������S&���fH��n=kf�^_��}F`]@�<�3���Z0���5����Ϩ8����;)�.�0R"*� P���p�);-�aq����o%���VJ��S�3��{��J���@��q�&��89�=�C5�߭rP���2�m�����&�&Ш,&��U�Q�}a0�� \��L)�mwg]l���*���8�qd�9����_]��sq�Ye�d�6wf��v�v�\Ō��B�s�򥯁9z|�y��'YՅܩ��'��`ւ`4Fg|n�[ڌ�@/U���O��+W&�]x@f�79n~���C��E[�r�3��_��AKCr،Z
�Q�g��MwL���i~r��TSƱ��8�ƙ�g��69Eպ�4��dL#��������i����7�kB7c��T���23��`���kC\��+o�Q7b]IK�8�1C;8\�#s��=��v÷`��GK�	YX���u0v:Za4���#8�-��Y�LL�)Z�/g���wf�&dP���@�>^�ۉ���
��bK������X���52��\��g�csK�ǂ�2��'R|#�N�8���|���%��5�&��
�S���Pq��j�i�&�!�=��F��|��f,�����;��W�?3��sk��|��O/�� J���������x�����3����;V�
?�h��N<��G��o�a�.w(
��$Y��lUA��?�)�C�O�͚5<�k>A=�fPn���|k;�U7Y>��y,��y��ͪ�ȃzmSW�}�f��h4�!��$S�L���ϿCm,��\��I���"Ҭ��D�����˟�<���>@`�gP��j/����Tv�1*��0�0������C���ښ�qW9/?�W�!Оj�a��F-䑾	ku%����#�qi�_���ݢ�I`	��g��i�ûYC埉������7����J��|d:�����&��D�����PI�܋�t��w�7y.�t�0�\��}��cK�UḈW�Z@.�D�%�.w�������\3�g����*�e�σ�U'-:GB
�;D`�7�yȖ��Dű����C�f��%��4��o���f�?��J����8�m�I� Wgvۡ���-����dA�p���~�$S6��2^�aJ[�=by=�>������Q��X�9�n[3R�i�2�Wl�W���$��W�A��
<�"Pc�W�^���yrc>�1�.?�B?�bQB��B\Iځ�](����������Z��>�USD�N���y�~c��$yNM�����
���'df+6����LF^�5)��<.�;e�He]T?��h�=#\:T�L�{a�9���,���R���W�k�<"{��Dך]iCA�c=/�|Fc�W�,��4�Iq���q'���Q��nG��&��zLB�0���ʏ�L�j�Q������+kJ�}��4�f���v�z\�j�,�V�EK�dQ����!������/h&F�2�?���7�,���!�>�k�3�HzuTc�OXF7�J �U6��67EK?��'�R~�������Vr�e��LI,����Zt�[$x��q����;��n��Հ�3������ƾ,�K�͙[��<m�x�\�r�ߧ3���\�e�y3�Qj��q�I<��M<��Auvf\�g�b묔�}<~�A�l�![�sPO��`����A8��2Rʛ��lO�=�,Ѣ���״n>6)<����n2�Y�&ҋ���O0�0�Z(�t�LX�32�Ө�JҶ��3&�ߕ8�[g�D�	��x�`ӑ�O��_�����it�<��@�M$�K�T��w��N�c�gQ�ȉ���EJ�g�&fo.�
��JfK(E��֮���~�#�zb)�*�.������8
������;��Q]֛��N?��ڃJ��& hR�?;���p�!c�vZ�w�u2�:?P�	��~R+�W����W�"��d�3�=d�>xmW�I�����@�Ҥ����Y��?�ݍ([
���$�s�촫�5kn�;*y���b�T�և���f�j���oD�٫�����@�E�����:�+�����4r�6�l�p~�ߌ-�n�쇧��G�w��>7���t���������k�ӵ
�� ���PT�XRb��uBH���\��+�нE$U��}��+��U[��5�_�e�
%����g�1㮳<)a^���]maOr�����q	�P���� Ɠ�u���N*q�I9�2�A �u��?����F�b�c�R�*@?"g�iAU�j�01�i<em��ȳ��ڮ��-_�D�����7�i��7f6N�+a�E�H�N��O�Wn���|vsp*���4��ꖾ��{#L;b�o�=��2O�����%k��ܑ�׮���G:Ͱ^�Q�������.om���Y����9�����n�4��7$���
��GV$�ޓ�Q��>�p=T�	u��Ί�����y���$��6�'��V[y��T1_a�7S=V���z�z���\���3��IL�	f)P&���U=�3<�4��ئ;��V���ОO!}>��b�P.�����T0�:` �h.������'�4��@]��X}5����� F�1����Z�T���Q>����>�HA�4���t������Z��D��Ao2���#E��W�O.秘b��e��R%i�OU��
(�{���O����EafY|����:�E���15�5�b�d?����d��� FԘA_#�Na��MP9L��������p֔�sXŁ�$�譚/������aFס���v��\�r=�X[�>WZ�O�رb��؉�<K���e�,���ļ���'�sEn��v�(T��I>0$�*�7�|ͦ���Y֦5D.�C��Q�$��a��,���p�BB���vp��庴K��j�k�9m�LXH\�z���ѲiBE��A���B�HQ���9�����\,�%:�92Erm���V���M�6�߲�������]L#JT�Pku�%{����ő��(-twD���.X�;�8Ā��]��Y����/Ptk�Os���Z^U�ax �<��E�\R� ��j1�����Mb�3�������xG�����춱t�Fq��(�i���;���F*�aM�n�2~��EŽ���'�,#��uH���YV"ov@j+R�W�P�?[(�����W�2ȸ��ڹ� ����G���!!T$S�Ǌ�U��+�.�t��0Ѽ־!A���'��|��{;)��x�Wm���0a�9r���(�ʭ��©uJ(NF�[����(��vxV��f�@��<�z�8(������:8rc|o��b8�^���J!�1����K�tdJ ���\@W�vӘ�q���IH~���~�6����a5AhbJl���a~�������uQ�0���p�k�KwK�V�v�7��+��+9�vP�UNK�[L6m���(�cҚ���6$�vE�.�z�#-�c�`0� �gC-�+/b^�:m�r38�z�,�M���,�m�:��x8�%�IyPʅ��f*,�gH(�����@q*�W�bj�I��4y;y��F��mB�Qe������Q��D��V!��E��LU�+ ��+�UOM?U�W�C_W�Gi=�R���}Л�'o�KT�Ҹ�Жa^�����+�ӱ����Z�n�Afv�`v�X;?�µ^��;��<�I���H�E*pQ0��@�X/�����N�j��\�(�{`R�|�i��S�8:�\~Ȳ ��Q�4��q5�k��6H���M�Z���O�+�3h�%jF6�ؙ�V�L@u_���X���ʶ��I3�*��^O�剠	����ekSG@o��j�At�S}���m�|\D|�M��I��Ho��(N��������{�j\cTq��8Q�)�Q_t��4M�C�c�F)}��}�j��#�\��_��6?����n��
�ܛ"��q��K[�B����m���39�$�ҵ���N����g�m��ބ���ZG4����!���Ip9���
�9fh����g�T�9|������#�$ڵ� l��J�\@G��,�|~L��ا0��V[�0q�8��߮�䝴4���9����� �v˸��Gn��j+�,�M.�l�;��t1���}U�l��T1v�xcHRwBطZ�D��
4�ҟt2�Ŕ~hu��������G##��%7�G�%���)��J��/ғ�1���y�?p���Ao(XlB�^���}Y+,w��xG��A�����<�L���
��_c��x�^����^�mx�z4�@�K�W
�S��?��(1�3��V�͞fH�fǖG<�'Of��S �M!��?īK5�B���v��?f$�9�Zp
+q\�o\�)��A#�`	��d^͝���2��d6�>#�u�?���Z��׌����ˊE���q��0�O �p� Z�Ͱ��)���G
��0{�06�f��fN�%�յ�G�"����O�����F�gR�c�%�-�pKr������ƌ�	���h����7/#%�i��VK ��d� '	fN�v��qMG���co�vt@!�L'��~�P�[HЦ��7t<n} ���Y� 4`�ҽ�U$Ƨ:���/�o�.�o�F��	I����¼�BS+�bk��MI�;a�.�|BF������	��_�o�7���_�r[gSDaPj�L��[bih	7��2	р��I�@v�P	޿���B�<0I���C�E��X"8��2bPU_��!1��f�S��sC?�T�kðe>]���7з^�'��t�ui�@)k��_N��2��F~���F�eC�6ծ,�ѱ��'C5���=�S2���즽�G�ך���C4\���fAc��:=wT*oa�C���{82D�ȃ
�'��*9#�05'j���E,�l��4~~n�������(�V����{I|'�����������h���-?{xa�vjV� jىʀ�����np^8����L�+ xs��%F�D�]�s�E26��Z!&8Rb���+�X�Pw�,�����gj�g?�`1��`s�+�h�hH�v���E�FT��n�V��Zڰ#���̄��ŪI��N�z�R ����W�t�?����l�K�g��xej�5�ϵH�0F�:}���6�����߂0�A�}�N�[ b���d�a�Nu'%���8d��QU�$�O(`�.�XÏ�<�_q�߅z����{���C��E�=�	�[�ճ7�-�q%�LW5j:�'#J���O��%��z3\?�|"C=et,�#x�C�kA�A=u=�:��vҝ��,�8�^���.��=���Ne=R��V�kd��jAߎc�,����l���crQ5z���m�Jp�@<7���� ���Ja֖����q�/�)�K���)6�FN����a��Ԓ���U�杶�m�����Iv��'�,iP��4n��9 ����&~�'N����.ѻsy6F�񒾊p�WK:�e%�)p�n�A��-.ک1�޿L��+5��`�M��ge�V@lP�"�Os5��"S�}��Y�y�z�-�|YNj�U�G`���	#�D�
{r�h8)��QkE0����\-n(P-������M8��Қ�ݭ�#�Ę�o^2C� �m�*Vlx�u˷��*����J����1Ol��$*洙� 8b���ޒ �Z?���W#���6�E�4&����.��1�{Ġi�Y�M�s��Pb�+^�p&�s�����J��a����K��ԩ_�w�,�����X�]�E9P�8H��~b�h�Q\�b�B����ʊ9`�nٻ���3m���1�|G��S���G�k"�m���:��<^����J�Y>Qi�6(>����낀�}��ٽ\� ڑx�5NU��{�׋ܥtp���l}�`�l��
3�!pqC��{wl�ivH���C��2T���Vw%ùK�H�+|����J�7&��)���?�k��§e�\9����:.X��c���Z���:K؋�(��,n�^����b>Nx;wz�5V�=�`^o; W"Q���cK�i�P:un��E!dzA�fKW���6�Y(�	���IP���ﻓL�婔��hӓ��-�=��|@���L�U	��PP�ø��S�QG��X����V��ݻ�u�3�\�6[s��89>�8q,�?r��.��бC��i�5��*[�l!�%2 ��9�Y\(/��u��|镛�^��[��_����z�Υ(��2�5�xl�� ��Y��v'��<:�[�����������+z��]gG�خm��\bP��K/�j�;'z�>��rV4~�mY�ӎ�޲&;f���mI�*��l*����k�S���cY�	����l��=~�t����ŗ�4P�����l�"���#[�d��&��&#؅�XEzׅ]�m����]����iIou�faO�U,�i�������c���6�~)� ����܍/�W%V���/3e{�º8�L6±l6H"�����B{�ڋ�8����HX�"e��䶥���Sf�6���d¤��6Dئ��� M�vXB�����h�a�<�u{\aɡ�h�����T����6I�'Jh)P[jȾ$3��%B��#��k�|�x��/FѼ��cZ��[Iv��9>
Zfꋶ�����s�vOD�V*���Os����\��q��G��G%|�E��)��ʥ�5��H2�A`p���I����)'S�Y�q�����8+���Y�V�`�aH�d�S��1�A@�,���po�
�ܢ�c��d}����G�7�_fǥ�1�A�(���8�P
鯝�O�2aӾG����5��ǃF6�x��\��_gJ���$O�l��"��K��.�_P�S����z���i+�E� ��=�]b��!����BИ)�����T+�θ�R��>���,�9���+�9RC�?��s�|������ ��O#�!(�^-?7���ݍ^4�i�8��hfا6�9�?���>	����)Y��E(c�b8-3�Q�^-��s�oB��Wne|��db�!�S=9sAK�J��X�#�)�8W�b�0�v�
B�cν"�olc�.�P��ɶ	��ܬ ƭ�_X
�CʵK����� Ne]��M����`�8�vں�5"��2�,�E�e�RH�n��}r�ֲ�k����:S�=���_~�4c���ϊ�?&M!���V�7ڛ�3o���r!Y��$,���31��hr>�}���+�y0N�O�R/�8�xYJe���f7צ��'�B�s��ȥD#j�N��u�I�"܇J�i��0�U@���fKܑ��.�,R\-�vR �!?z?����Z@[�� 9f����?�Nu�G]]I�
�����n��n-m�!왑�e����C��D�5_���E�,��%S��<���̹��ڋE�Υr���7���D��R��f�\���ƿ���ʹZ�q�3eN��ބ��2�v�����F�:���Y����aϭ���� �զ����������2K�Ы����S���y�-�4&(:�����eN�T�)T�5����+�Oo��>��r�G,f4K|�����
������3��/��w��0١���B�X���.lC��w)N�	�^mo������t�M�R��u�ԧ�yKj��x�2�Eυ_�O�c��~�Ԁ�M��HB��)��fi:��[-��p�5uO�R�l���kfę�Q�..G����.w�'$�Y�\��g�v���p�!��_���-}Iu]�tZQ^o��@�+���O�A���԰;j�[�5�����Y����1�J��z,���u�G]5�1�_I\
�cw${�)A�CS��p�A��Evw�jnG�3;4���5�vYi��/����{E�tP�J��±1� R�<�y��*%�E�����j`f�'A�%�Gk*S!^���A���D#nO>�?r��������9 *���;��L�'~���R ����y��5��_ƴd%����YI`�=��E��+ ����R2_/�O��\�UN�
��U2��쏖�4 "bk�$�.n1S �oHN����B�й�X~�q�*�3�=1��Tb�����]�3��E*El
��D�X)!5�x�2�������\������9V����(g$�h��#�M�5�D�������(�x}pX�4_����\���7� ������k��Y�'��fPR�/�X,�	l�	� B�m]��9a0���QR��$B-���]�Dj%���a\:�_`Ƣ�ѧ�*��y�1Y4>tj���Y���wrA��p����L��5��m0G���*C?.�=��'�)�㓁�A��,�@����L�6m�s�t��`��&d��$f�0�d261o�K�ܷ�"˿uB�n�+�
9	�����M��̋_����*�Y}tFtP����N,� wV(-�l��Țs&^2�շ��
��&�>��F��e}��EX�V��u�n����u|l�|�x���K�^��?L!�
��s��_%CR�3�12�3o[J+C�`����@%�|Q��~�%�h�o�n�t	�t��Dܗ!�|f\�X������~�ߪ�@�8�L8x�9�y#��\��W�#��t(���^����b�4VU{jqpP�i�����P�N�2P���S>���6Ml;&pÃpc_�ɂmV*�h�����ܕ���9�[ 3`�-���y���ag�Ne���\y��pܲ�G{��z���pb�J�G���s�\��i<���s�Ə>�#b��a��_"r߷��Dc�PҪ:C��s�Ѝ�1�����vq|x'WM�?&�D�6-��&�H�"��O0���x�mL?��F}�D3���/���R�³<SDx�"?G�S�G����9L
�U�>({g����Bzjg�\d�+A���g�O�!����F/�Vy!�V�]<m�gR�h� VH�@;yۗ^<�J�Fa
�Wљ��N��7�0��[\��yN�en��� C��# �5����I�8
OQ�mȑ^�y�{F�Ş	�f�*c�o
¸��'兊��a��չ%���+[x���M��z,�U�<Ͱ�!�w�=]�:���� }7ف��L6vD�.���V�,k�$o,�t]�@���Y���\Ú���8[�8ۼpz\�"[�h�ٰ�&��ek����mO���	(3hs�U>�A&O�_u����_����$��=�x-��H]s9�r�ãd�?��1�X��#��.+�-���?77\��xc��
�4�8'�y�HTÇc@ʏ��[z���o�.��e���+���Hh��j���/�K��=h�}�~px������Jѳ���2>*� �FP#�[����A�+�����H�b��eUC0�a��&]����$�NS��AQ4�j�a���M?���� X8��F��Su�v��Q��Ķ���tc�	���FG����{x%Kb�X؈x�h�4Y%��^uz���[��V�V�D����
Olh%��zx_
�o�5�0Je~���}=PO��T!�j�V���F����:Rԙ�WNN� �wVd!�7(&�e˔�$2��T|�I/$p�<��^�}��P�����ʟ(�� C�%�8�ˉ��ѻ.�at���/_y�s��M%���J��7 M��������U���� �>a��J�P!��eP�Z���������JrƝ�Ǡrii�p�*,
���Ǎ�`��st�� �u@1L�����j�l|��)@R[x��[`3�oĜ3������̜hŠ%{D��Q�|�4����.c��u���gۻ����|��mQ7�+�&E�^aTe�9��9h�{�D5j7DMѰq=�7��S�[T{�ٛb�ŭP�7��u���a��H%�{��u�T�D3I[�Z�#L�L^*��hz
'㰸�BiK%_��@����B;e�^$���C�z��ɰ�L�"�����P\�)��P#L�35:�ہĊD�v�|�#�D�v��4�C�h�+��kn�P�)9�YP���OQ���A��b��ғ��!��|-fg)PE߆hk��U$C�AQ�
���D�ަ����a/ (���/����E��[�`�g�h8�Β�_�I(-���[g�%�������)�l�����
�C1^S󻬕J�Y�֍3�b��8�J��z^���_T���*��+�-��A[�h��lvV7bVa��U�o�1����k�'���o�J`M��3�+�#��y�L�\.g�(2��Ƭ56AG�/���9���2��El��k�	�s�d/Jt0O�0�b��Xk�vn�E	��\rZ�����*����C>��F�Ԅ����~���ȏӁ�K���i��4�赞�s(�!.t��^�a���IΛ�1�ҿ�^�t���Z����<�xF��[{��$������� �O���Q̗����7�~��8v?,���w�M�U�M�|C'�� �`��O�s�u��Z�e����]�AS���8b�;[x���&�J{���¿H��kB�C_1��IR/�_,T���Ia�ZW�CQwAdLqr�a_,�!�� �m{��;�#�+Z1��%ṳ�A0��� E�\�A�۶�!m�R!��1&�lɕZ��v���ޔm�%�x��)�A���&�5w��ZK�da�O�8��� �����z�- �ütݥ��~��D��/`��
��jl���JiB�vk���U-�O��W���P�D����i��X
����yn�g�l��g%��!7"�0b�.MkW�-0���?\Ŕ�a�V�a�^p���ʔ�/i��/��.;$�䬋yǎQ�#�}~��'�?9��d����#���h��+>X����@�T-S�▅w
�{�r�	�VdF���LU�a[Q��l΂��G�IGt�Fϴ|F,��'�a��Z!v`vj,�Ƥ��h�a]�D:�j(�:�V�&a#�E��3�����x�d��a��f��k�o����V��`[\�N�y���(��M!T���n��m$q�~sfI�G�������c��l��'QR�V���9�QZp5�m��
GM)��BOåc6A���w3� ��Fb|uRo�;�h�+��H������Q�J��T���~�5�z����6��U��2] �g^F�����UH��A��Wѫ#�\0���
� ;o����Ι�vg�Ҙ�����Sa�;�Y!��d-��A��sT���|�(eϑ�����.�N�iU���.�su����/�u:��9	�'*���xi�a "$$+N����)��(Fa��^�BUuloF,� ���:x<��Δ���M4�&y�� �*������p�vؑ�Ixoi_�L�?� Q<�j�,�0#�.�[����\B��4�b�}gH���#�J�`;$4;���IR��"�vȼR��D��?�l1ȅJFF3O�9���zw��򧴐����@	��sf6�<lN8�Гaʒ�m����''��ۨ���ڽ��4��Ɏ�K�#���qn������plKX�+�K�{��B�>D�H]8�M�&����ٶ�؂�d��7���?��7+��A0��B 9%�~�ɐب���kL�j�>)�C9��^�1Hg%�٘�!>}GÈ��|��W���"�l��"��ɚ���i�k�Q�dva��y�0�f�ӛi�,�����@�=a��ԧҼ��D�j8�� B����~ܰC�c߮W3ci;�j?��k|x?���e�6���)V�N�m��B?����ΟeH�}.8ZxVw'փ��kJ��\��
���6an�S�ٸ�gT�j�`u�H�^O+���3�������q#�!�/C+���[7�Kk9��GTq����PB�*S;�01������P�� 5�q��bOG/�.�NY��A�j#���%�=�ȪW�g�F���C����mg{f�j@3�TMQ �<���dҨs��2�q�oҴ��Gf���X�G��a�4z��3mȺ�%~�O{l�=�K�&A��q���)�ȼ�>��^�h�2g��ܔf#��u��k�J�����j�	aZ��^��Ʃo�д'�A���2h��|ޞDV� ��!����S���h�B���Th��:�X��������e��]�����k#�<���5Ս�e�������R�&��Id> �lV�0���̸Aplq�̇b��1w��a�~�!��9W���3=�S:NU�t1$��h�����彺;���0
���C�#s)�n��X�Y$��L�|z'����qj��؈�%��sڮ�oB̏ި�0b�܇���E\�N1�^Z��&�T �o�e2q�hA;��A��(n�t�!���ʼk�3d�R=-�h/<3��T�a�0$M���N0*���i�`K�~Vt4�.��*�ln���5�� ����8��
���?�l%w�t�x���<�{]���.y���s��K�w��Sy_�ݲgM�0��k�%0j�]Y�GW���'�<��ԥ�śp�H��X�jv�b^Tv�|�^�hd�u��Fz�+���cg=f���'�m{z�� [�|�E$��v��/.��p�\�c.�����6��j����.?�:�(���w�R�v��s쟤)�29�\w/lI �ۈ�a�,�1G��vmVn�z+s�[XҋhGPjR[m�b�VKk��$,��Et5o:V�En�y`��	x��!���z����G焛��%�]���
9�eH�1	Y{�Y��6b��
��ų֢8v�q�hP�C�!�y�RCo�,RY���J`�	o�s�,�z�̱��?x}�:x$4��@d�)U�7�e³�CRSw�Yn��<����H�)G�%�*�:�Ci�����LT,�V�Fj���I�r?"ɠ�{��y�m�_;�q-����؃2���C;�m�<p�W���J�m�4��`�tpѱ����kmgUU��#����w���Ԣ|�SAM��
-U���2�V�s�,ԧ��H5��P��R_�j��pRnɱ@�k��yK���o��6��Ve�\��3�Ϝkw�uF)��U�4��T���j�ߎ��E��U�ԅs��a���b�Uf|JU�����^��o?�d�x;��z3b@�U��20�p���D�ub��9or��p�kO��6֕�(z#�v]�8=����S���A-�Y���	&�����'���'=�o(��"1s(z�a�����:t�7�h��?�ƶ���p\s��=�'�F(�V��;w@1Ki�<<,h�c5�%\�w�x2�3v�
�Տ���8m��[I;����|����*��BI���0�p�e99���F�v ��Y��/jjek�G������7�g�.�+���y�	l����^�T�ZHR:�*k��p��}^OW:BH�_tS։��j;
>!I�2n��G�$��͔;�ɢ}��?͈@��/��VLn�U����C\�r(ܪ�XZ6۝�:&M6e���un��e�3g��������jY�`^ek4��c��y^:����9\��ؐ+��<�M��XX�}愯��\�V������C����_����
�� ҫ@	$/�HfIar����f=@�I zDt��8��������d0(!C����"ǉ./?��^��o�T\Q�m��jE��GE^}d�����m��GR�$I�e�ϡe ��j�P�����';���r7��m8�{��y|�̃kg�zU-�/0��[���x<�3�Kǜ<a�BW
��<f�lCŢ|��T�������~�F��H#�����3�b8��8Z�W�`���5�һC2�g!t/�����4��=�L:$�,	8r��t"s�>׼�֑7���ЎB��IA���ڨ�i����F]-�Э�Ƌa>�[fu�� �I~]�����-k��p��A��/���F��Q�U��e���u�½7�X�n��$��N+
,+�h�V.�X�#�Q8���2�Ғ���>��f�*�o cV#����H��rN��@����im�u�pp[����t��4�c�f�%}�2w*\c�n�Z�Ow8�K��ǆ��|����;
�f����sVq?��-'k�r��Ϲvvl,��Ğ���`��&Bl���MbΜ�Ŝ�	�<�w�b-�m3R�yx� گۈ����������[)�̤�1��O�B�H�`��<ER��Y[��[�μ�L_�Ëi!a�{�'f�$���b��M��������ӭp�k���C���]�ِXd3d�d]�Κ��!\O<E�s'�)N�^�0�m�(b��6�x1��ϲ�����B��#���#�e��zB?�"M����gQ����A&k똪���a���v&L���!�$����Q��\�te���UN]�r0բ��? ��'R�ã2G�01��ʁ�ބ�Sw%'�=[J��d��^g��ge�4f޸_���oq�<f����v��=NqH{��.Uli?�S��/�3�*8/�P�c�zqq7Sɹ�C��fJ�U-q4��n��׀��\}o`�}�&� N�04=�^h�XFusV�7V	���� ������<*)؆�9�L�\m��ʚ�U\]�sǯZL�십���c�^A�O�Xv��}�Bx`�ަ�;!�R�Oi(^�<\�)���b�8�p�?O!���r�.~�+���I%,��@`�[/�`w�QQ��:���%^ �
$F.�����_Ȱ���{�n���Q�b#[��cU�*c1�4�B�T51pn:�6���$��dB�vz�x19��dZ ��Q��U2ǫ
�{T��-��6<�唙I���
bt��~#j���m!�;Kju�nOލZ~<�y��ɇ�!� �u�[@�ښʍ�ф�o=���þZ�˗B�@�����O�Yn���j?�9�\(T�F�dD���u0�;���%|�+�����׍Xm����`9��#>�|a�i��1���NHv�l��;���1�`W
�Hꬷʔ�W� ��r�l^MsRm���wI�1Ő������AV��GQ����Mg3x��j�,{�p�D(���t |��7�T����.R�����?��0���5�����-��1[B�Ro�� N�T���`��h�-�I��G�T��\:5љ��s�h[��٤FxTһ�g��"�^� (��V�N�����7�������И-��X��{����D3�4�ۙߗ���Y+����!�7䔿��ھ5��I�>t\�$�`d*����w9=+���f��B�v���Ou�*~�׃���F%���� �Twa�dr�'��A�N�ۊ#�����dA8ݣ%溴=�RGoF���PZ�w�n'�Q:N�z|A��Xc��f�*u�H>�υJ��gi�[Q�� �ꆰ�v!5���B�AC��.����5FGߍ-�EE��t������d���ۗfp:r��ԧ�5nS�ש/��]+q�z����*��g64Xi�ZC�6uBI�-�T�;�L�â�s����귂ی�L�Ff�MzKD����T�h4�b�q<�7�h�MHu\�.�y�*^�\w��������d���Q�5u�I^
G�<��k�]"�a	�����S����|E8�g��a�0Β�n˲�R�!rtE���j� �֍�A�1뼫�2�Y���g9#��=�Tu׭��M<a���vs'�_%�W�&`��{}�.��-���R38�k	������1���t㸶yή>r{XF�����UCW�|��T�\��{u�Nʍ�+.\yQ]J��Z�d��2 �՟���q��ehU�]W��+�+��=�__�H�&Z��\�,�����Y�p��'P��؞���{��E���TΦ��/c�"��o���*J�Q��l���:<����
8��	o���3�`��w<j��4یh3���gB��������"��-cLʯ���U��M��2Bcr�h��X�X��d���G-!�]H�W�8�S�w�XqF���k���a%O�ŋ��V���f+0:E~(��9o١ٌ�I�C4�'����ݶ��ݩ��n�(�)^Ʀ�;[QS�JT^�� y�f��@??��63ժ��p'#���\C�>ܜ�S|�RR<�'�r�/z�|��Q2��U�⢔/h��p�"ݰ�hB���=�~K�?�I���k����d�)[� ���^����|�4�)畠���[�v�wG�����80�q�R�*r�۲�
J]"��*�s�-Z����]�l��	HK����UR��6�"�֘^�s@����G��Q�g��d����蘋�{:��p���h �� �|�]h;]��ʯ{��Ͳs�׷q��
����b���E;H����X��R�3���r���ϳ�8v�w���-4��hT�*쾨9>ds�UF=Č|IRo� �5$@w�J���}r2��ޗ�n�D�7�T;�9��Ѷ'�9�$P�H�.�W�pVXoX-�S�	�ݵ�M�B�MJ.?�oe�f�9W��4S���ފm�'g�p�g�,=�=[���T7���f�h1S4�a2=��rr�Z95�r.�h�� ���j���FTek(��lMv�> �xT���R����I�e
�?��#�C�K��Y���	�YfK�aS�*O�AlNr�3�<m[�W��ӣβY�d/�d���$¡��e���i7��H<����~9|�ݻ��W��T�ge9�T��{hO�!Ј�'��n�"����jT�)�=Q�Q|�4��]���k��L�;0�Ej#��g7�����q��TK'�}B9_��Y�44vL�`�y[�GXMA١-A����_3�M����׮�kލ���pʟ�fFl�m{�ɡz��-dG�ю�+�o����P���`��ś�-���(5���R�C����ϸ�*�� '*)��j�n�R�n��b��9��tˣcb���N�U��]�S�^v�JRg�]O�6�C�IxsYk�
P�M��9����)� �!�&%����(2D��%l��!�ko�D���@:���=��cΰu|T���p@Z$�p�ϑ��q/���ٺ�W�Ǉ�
�3�v�j�pd��W���McN� نihv���|Ńs�x�rU��||�ʾcYRw� ���� �0[�Ï�f�r���<]j^�=t{- ��˨S���\\�&m)"��sv�`�>�3�v����7WX!�P]ꔱ����G�p33����:�]���"#9�W��-1�8F��)�� yOѦH|����toVdn��GV�XQ7�����l��Vq��g���*��n"��d��7�u��D�� V�&ȵ|N%Z�ΎƬKһӏ�b�)��Cp���	H��`g>�RGW�+4�W��^ƀdPa�ޭ{�T.^ V�SJk^, @g�P���O`�v`GJ{)uЀ}�w�fC���b�t#��u�É0�Q��Y�;%kʈd�m��n���*^���AG5a�ӄ���}�����O�P�G˖�N��m�������&���M�|(5AF�[�ڞJ��
}��S�3ZN����_OI51zTỖVêr�б��Gz
BF^�s��ĝ?�bv�U�Wt��B�C�l }�4�d�F���Oj~6�W��"��DW~ 玑�<�JY�\�<1c�$�O���{uhZ���AHO����Y���!<<"��d���ؔ��.��U�v�5�Q+l�(�N�Vr��U0e��_�-�d,A�|�*�Ҝ�Ie�Zz>9A�ܙ�\7f�"���+-_����H��شO�p7�cL5�B�A���cR���0M�Un!Zz�PM�sQ�M>E��D�jL��n�/#%`����{.`�s�����u�I�]�Ǿx��M�c����[|M*[�A@�#G7`f �����w.���Z��C4[�C����	@XتL�q��oיm5)�����yk=CCŤ]�#�T�h/N��� ���Z�����x�{�ۏ��	mSX=�zy�1�����e�N�-�\�vs�+R�^>"�jt������.v41�O|=v�\��#���칾��H$C�#�8��6(�R�EY�����E�?�dޣIYcN%��f-�m�� 횪.I��)��YɄ柖TA)C�j��?@�q�]��f.�p�2���k߾�m�x�Of2��Z��{���~a�=�[%q�硉�&�Xet�pgf�-�ʠFkK�����Y��������xc����I	��?j^�Z��x<z�茳��H�5�0 ����l9��E��]��J|�T3p��W^R5*I6�mQ��ia�����XL�7�S��
x,���S�NWR���h�y(v�oAZ��7�;����cP�٬���x�,?���n� ��9Os�c���;���E@$�a1�o�xyyH����,�/���\h��m�Q+�b`Z�a�����!�c�P#����n0��n/��w6ă��MU�(��Mǣ�"�%�=7�qd���<ZG���4��͒l4�;��H	P��4ʼ�x������a8������A%D��:�n��F��v����-E�����s���ǭ��K4:n���	�_�����xTZ���n��>!�B5c�� _�
p����O�V�eH��ޡi��o���^۴�� �����bn0��u=d�5�f�HI��]e��ɲ\{���d�,}h>�S��'�@E�,C�~]jEZ(�& Y�����J�f��/,�֥�
��(�ǚK. $`S��=*˧��\�jj�Z�&2���جe@ñܲ-D��ȻdFu,M����:=��AΥ��S��3(;�|�6��c7G�����<�6�yw!w�R���r	F�lGL��Pw,�+`���2�a 3Q%x3y֓P��ѴT��A�!�=i�fɂ��K�&���%���'��ӌ��_c��c��o���EC��p�"�)��q�z`T�*�ΆyMl9�2t���H�ř}�����1�����2��ij�j{����m���0��??�C&�W�K��V�.}����|��z�}b�l;���J�g�=u�\��%������h=�p-�k�a.�;�r;�t�Q��M���Z�Lr�璆�+�&����� >	����J�%`H��g����[���/�%8�>�0�J��n=0{ʨT߹
����.◼�h��ꖑ5MĊN�
R�ܠ�R<�T���?P�%����Ä8g>��KwT��fg��ޝ����y��s��;-�����G��q	$�7f�|���C��	�S����V{���_f�<؃pߒX�+\�t�U__�l�[�n�)��M�N��8���ۍ�x��V�ƸSL[1ߎY9'g�|TM�0Vz����9@+��_2���TǓ��i����=����ȣ�����R�D��˷��hK~-1��Ĥ��y����<�5T�N���Kw��b���&F�@4��]�r���$����V�����ӖvܝEWZZC�;���Г�g!z4}L�,.���=ħ��t���5��s\��deٞ�Ѷ��=����NPA�^�O*�*��lh&�_�ct�i�Z�H�l<!���*����A���"4�Z\��Yڵލ�aZ�z��;�̃�L밲&��c۳$�>,o%>LV2���*����6k�	.��v��v9�;Ág�G���W#��Hm������}(�N��)H�Z�Nlo�ڂ~|U� `yJ ?����AL;u�S<F�E|D�� ��eS"Ї{T>K,Z�(�J�����.��B)?.߄U�$��B�I�PBX2F/C� B�$^\�i6d}E�t�Z_�5C!��cĆ�L
s?�٦��|2�Y��J�&&�E��|C���bG/�i:p��UWi-�u��SF�TK�%�>'�S�(����$��>��6�D�#����`�5�';��K�_&.UWI.�r���ѧ>��i�u���)�f�U���n
�0�T���>#p��C\@5��k�rx����E)��Ɓ��Y������bjB+(g<pI9�/����ܽ��T�#��FIx��і�2`����v��Z.)�sF�����C����d�8A%��#�����5_ýr��z[��L��,i�y�9�=�Ԋ(�f͏�1-Qp���*p�S��q�T�Ԉ��Ғ�(��w�O�ld�y�*��M�<\.���53ꋒu6�>��Q��A��6�%�q�p�ʨ`����~q�o-�=��,�`�ہض����W�L�E@�~+�-^J��Ϊ���k!�ʝ��{�_�{�?�r�1Uy��t��䘛�&�'�,���}���q����Ds~�/
e���1�;B���U�a��$KV%%�&wA��6QˡMH�����֏NpL7��
Smj��P
��=����Hw%]�VI6�"�݁�����I��/P��)/[g�&J2�*�Evť�s	Z(xF}�N"f&�5g��e%��{Ř .��x����%�CL���R V�1�iҘ_)I<#y����G��-�"Y�x���SVC���ު��Y��^�/�}W�ȓ���<��CF��aSay�c���	��%MeZR%�r8�wyL��7n���
s0��V�*��ߓ�#�5����oSG#���Eϲ�������w������<K��aDfDA9��DG	]vr�@kLi7�:#�)�L=+vܐu�̡Q��"a\k[X��D�k��WqGX%����I�V�a^�<��F���]1����r;���+�`����W.�L/u[B2�EI�Ս�M�7F����?�l#Τ	.�0�)V����q|%�s�w��Խ! �����Ƴ��n&p�d�y�:��)�Vڳ0q�;���@�]���$����x�;�����](ӡ�&Fe���'c�
!����T�:B�ԗ��YI�_�+�
�r��s�����9w/?�
�O�Iї�K8Y��Ș�{5+u�G��>��娒|h�o���x{�}p�1L�`(����_f8� ��$s��b�WV��fZ*{�W} /n���d���z !ο�:Gͽ���� i�n�@�2�]��d����
3l�s�%�������=�˗�}R�o'\_�X�ƹ�vŝ��[�����^��O(R��h�I�3A�Y�&�#+/�̖[5y'/d�9c��jX�uZ���F$����#�>��'("�hi��6A�C� Wd��ݐc�h�TI=�\aB`v8ؙcO��mάܼw8�}�*f
�O+Lj�z��0VZ��^��1W]C}cX6�Q����r�nP�����~]�	<���Ʋ�Q=�G��pH�t8�J��xgZb�7J�T"��fE�q�K*����e�[Y��~�< ���(5��s�}��UG#L.3K����&�#��R�\��D�OϿ:���mף� ږw�G�Q��u��?�pxS���ݝ��T׎9�/��`h�/�Q{�J-�J|�R��J �����i�����9��O��Ȝ'>�P�c��%j�{M�dȕݴXrl�����`|�n��НC0�����-S�F�_8^G���`�
��׌ج=��騸�뉭��,�ѹ�$T����P*Sf��H�zݝ[� bam���B�����G��C3�]�1�|�҆����] ]ݕ`����.�fz썼�	ڎ�ը>�5��F#�b���=��v��c9"�b�+�7�h���8��T����S���=(�ޟ�K�ݳA���c�8)�����3S򨹥w����t���I�&bL��^�+5�����9҇3oX�P����J�z�-���>;v^g���*�c��ţ����_��#�!��nI�\r#�S���AK�q�I�Y�Oϧ�"�,l���V���z���s�Ǭ$5!n��9̚�M`V)筨��n�����͋-.l�@��$Ǿ&��V��c����6?��C�-��HF���&u�-J�л�z�a3�N�آȦ h���'d��B�Z�R,��F�����#Rv
��<�N '��:�/��B�s�%U���7`_1ӑ#K}V�_ۦ6Ԁ �	�ڴ����I��]}��X�i�S��d�P�~�Iv �(�s�	"q󵴙ݗ8)�E�ӗB��>��^�z������	PV�G�S7O�) ��7�6� �}����4��r�m��KY9�Z��(�b9Ꜫ6�J���U��߉��'��V�/�Դj��r��5a��>Oi]bX�Cs���Z؅���
�B���3{5���Y��̃�m�q��j�n�<Н&^��n�Z�2�y�2��ɱ�̨����#�4��/���L>�:z���n�����ٲh#?�&�<c�m�|
��)�(�s��2~�^*���^�F���t	C�(V"��?]L�j������!���Cv�mU������L�,͵m�z(jy�ID�m�1�ߛ�p�\?�4��@tU��? |��@g��})�$�X��O��lu&YJC���2�q?L;2Q8��f�>n�u��0vMHy��=�y�n�jTz$=���L(�$�����?�wX=*S�d�̴�Ƽ�D�����c��u����ib���ɋ��g�;�{�q�!y���a��ɼ�nFI"�Er��r蒚���3*�n��d�<1��6-h�Gu:c�f���	�h+p�-&S.�U����aM,�Wb�|���vF�^�O<���m����n�6�x]ūc����FM�:^\�;����U��b�.n]�
m��Z3S�^!��h<����Q��q�fn�k�_s>���"�L'��[�|E�@;\�!=��vK#8�z�g!C�4Q��߾�x��O������Q�Ŵ��T𰔵��K\��|��&JX4"eJ`a�۱��T��yq���d�)5���K>��'����X�=`n�T�#���U�NY�^����-N�rG�y�v�npEb^F�;���j�@aU�s9�.}��(*����3k��ŋ93sŞ�����&�x0��h����Yڡ���gF����_��(��3��oɧ�k��!.������k�(km����C/r5�by��K��7�'�ޡ<�v��>-b4������}5hoS[��t��ܷ4�G@Ȃ4 L8�>z���z�%|��P���`P��v�4DR�����EQx2XY&]�o^�,���S)-( 
��6���͘L!���%���+�o���G/��-�t&�^i\�,3�����(���MQS,��c��3Ζ�ǚ��٣��<�.��ZX�x`
�91orPm�'E�T����p�����%�2S��ն,�Bwٕ�y���$�����9�����	��G���,]��G��6}L�p�vez�wI#�bK�o�}����(�,�?ъ����10������qP)k�+�$�JS��+�mn������{�B��c/F���Q]���B/�_']79�v
*������*��A�]���d�����Rx�!ٚ˴��ș��u�P�	W�A�20�4w����^�Z5оQ�O�֬��_BER�Lp�BvM�M�jb��%n��<�S�����-��Z�>3i* p����d����?�����7��Og�kWw)�6ߨ��i�Q��q:o�&̵ʦ|:M�܊\d ȳ*�뢇����6��8�\�Wf�?��^ؘ��h^Gjr����o%�E�{s6(�M	�+���+��~�d��ce=�ԋ��'�棒�ꔥ����@�@�e�����q�_Fi���\~�nƐ�7��8E���L>w/��������B� S;|�-�((����d��N0�3F���%�d�}��K�7�J���?-��������/d���ܢO�&�����);���O�U����-�ع9\�����ʬ�L����E�U��S>,v�B�1�H 	J�@	;&��&+�B�`At].>�:F"��t��S�j죠ѫyX�Z�d������!
Ԫ7��S�#@�HI-��"��~���θ���'pH�㣛a�d�~a����L�w�w��5M�J�3c
�ng�@Y	�l�a��Q�-��u���w��I�
`}�E8A��b�/���׉�ӽA3{Ԑ�S:t�i�V�➊d�o�����T� �.�(B-@��dy���1�+;i炶��p�G�$�\W�x�vs.�G[p͎a
�#r����Q�w;�׆z�`��V�*߰&��k��\�Z���(Kw5���n�f�ఈ�/Ew���σ<'oY���%� ����::�)(��}���L�zĜ���L?�$3�d�&�+��u��^�D�[-{��gqv�Z#��U��c��<R'C>����	�l��%���w�w�����rm� ��>�k%��Ǌ�M��s�K�'ao7@����.�X�S�>���|��1$zg!2�6��X��N�~]:%}�/�C.G���ЁI���=��t��.�:�=�s�{X�S̖+#�ly��Q�u��0|#��r͊����Zy�+�q)cxy���Wd^{Y%�6��sa�?�#���k�����#��ЃTt�7X螿����9���@�,%N�ɟb���KA\F+�K;3���v%�]�Yd��m�8\���
����fC���<�6#�5݇�����Jd1�jL�j]��\&\�W�R�s�c��v��t;�9��.7�JG'G�@���f%���T@�s(Ρ�u��YX+����f��Z�O�N¯���Grz)�#�,M�Q=�fK#Dv T�zcǦ�+^ �h��
܅R�-�*�������w���˗��N�3�g0O�HOÕ�.�Ĺ�L�ys?+���!���kK��k�`�+�����*�OǶ
�/wP
$HV�׼*4�����>���	(� ���3�I� �0��-r'�(���P����|qR���[��N�T�u�qu`����Ath�܇�d��ȇ��$.>_��EvUb�cO쐀l<}�Y���%ò��	m���ѐTN�:oJ�X���;A��B$�X���7��w�}:�^�;(�>��ڳ<\v�$�s,apwG�]���B�	מ����1���Lɒ�(�#�b��f�Ҙ�B�NfG���$��lgD�>�v��dpg8?��$3y,���4�!b8�##Ő)f�w�j�w#�>;�[?����pg�[]�[Jg<���D�WD�d�K-!������Ja����Sr�ެ��&�9�� �tUn
���P��:�X�@a�2� ��Ⱥ�&�����#�zw�߇"�cC:�#����V�������M��7r��� �!���v*(�ojʢk��7L����_��p��^�{��J_HDa ,�T���[C|�}�Ax����`A$�aY��s�����*s��D�6��'��CyI� ���Q�.f�I��������f#�|�Tg�m�t�R��{��Q$r�l�I����׀�Hi�%�n�ȖN��6/�lBݾ�*�K�g����(�p��U��F`��#i�{�
اڮ����<(�&�Q��k��V�����7��a��E�D���L9vQ,�ܾ��D������ق�\_Sal�,L=�}鵱�!'l�%��tY���^�ͳ�@����pJ`⸽T��L�OGY�T�䨡�"�A�<��3����X3�@L>H�����K:��@��Y=�SEH+%� ;�.G��c\�i�Z\�땊�8�P����띞K�����>Q�b�����8l|g4#��<2L������(ȊOv���aV��PHy�����ޖ���w�r�Hè	�	����(� 3�C�c�Q��w;�q�XɺOkTS�bWǴY��查:����q�C�Lm����^� �Do�)����ͩI'��66���EJ
�����4w]�� �gF�$G]Rǀ1�m�O'�W,s�Ŗ��ޗ0����R#2�jk�.p3�8�F[R-{���N{��R�l�o��H����؁"�P��2s�Z|��i̎��[m<[��r�eo]5SrK�(R'��Ë�A�ȰRٜD2���$RCq�؂��7����Lnx��w'�ڹ$3�F�4-pp�]@�9'*���Zn���`Z�0F/�	�;A�����},rܕ�\����F�׷��~������'�[��u�)G�6\�vN�\�3~�{�������G�W10�	B'Y���֎��,� �U�Y�Mx�"f޿ԉ��-8ED��3�y�,[����g�����O����\��F���G��@�00+���j�;�Ԑ 5�t8�e5W��~!��y��RC��n|e��*����֬�Z[H�w��k�l�]� �Tĕ$֞�(����9nm��]�ayA[�t/ �]��,-�UR�ĭ�w�#TRM�R�ˉ��Pt��z�n��c �77==6��Ҹ%T�#�8�4A}�����S��!�d���E���N��n���U���<霒6�~��JD�$��udi>�U���Կ�����Λ?�u+S�wٯ:�5��;�DǄ߶����K��p�\����^�#���A������IdC�J)��2
&�>m�g���iv1(���!H��	��+�\
}����
BV�v��g����Wۺ�B���Ɨ�.a�y�5Ep��r#9�Ⳏ�F<��@|�'��b�p7��*�0"}�������վ��m��71��}s�@W��l�~w��Y.�v��L:p������=	��#	����_�c�ޮ>�ajG6�Sc>V��a�����Ѹ�S�7P ��V���\\=�G���㡇ǘ���(}��p�l�ktt8��?_�^Ǭ�����3��9�=���Z�Ü֚����"�el���l~�4��:�a�V����
I���Q�ty`�'fj\��B�ʪ �$���C�$��}�hfv�6j���ޕ����I��ٔ���U��#������]y<���d�@W���&�ί7;M1�͏Wy縑3~���k<2����mU}n��"Ј[@��f¿-��Df�CT!^2�r\)�]\Z�P�fm_�X�K�wk0�x�LH5)~*����8���#�rd��Ҏ���!������kg=W ������pe��65��5>d�oc�w��c��e��Z�O	a���?;H����1"-�Gw6�S�������P�a;U�/GƑ>	h��,;o�h!Os ���nC�C[y��g%5�i
��%��ⱌ3��L� �Q���e ���ʞa��$����{�N���R)md�I����~����}\:uB�(�k�~�
��B�m10Wz�C���7���˪�Ci����@����'jP�?8��y����ԁ�������[�j�w��c�ːG� �a��ll�Z!Zøj~}vO&����o
G��~�b�9ɪ�r��������5�[aSs��c��.����F�u��6i+����&�ľu&bq�x%��|��$�1M��F���h.��j�q=g��Io�i<*d�Ծi��@���	ښic��i)O�Mw�ڼ7֞����ځ�m��f�v�~��A	I|G�|�^��e�u�u��A%�t�vP�I�R���,F-T��z�	�}x���^ �A�u��T��*�;MSw��(Q�'�b��l���Ǔ+��O��[K����]"j�cz�9a��M�0��}��J�y��F�iaUH*1�p���r;�x{��.9h��� ���ؤ�q(R���Z��N#�&!�E�0%T�  ��E�/H��	��n�;���2zi(�!t<�����E���26ݻ��2r��� 8�yC�A��F�k��r4�{CZM�o��������w�z��m�ؽ:�3�O+&3�5�8�yE}͟zUIn����]�Iz5d:6��,����Y'� f����%�����=I���+�P�wKF���읦)I�$F�$�y�D�R	�*�
�CC�xO����c� �����)ůq��HC����=�����8�����N�+�������C-)��3M~�CrI��){��F'�c�d������T��Q�$|���VQ����`*���~���\�n�8z�k9^G��><xu͗z�^8aJy���̝�f����yd͏� ۼ�����a��1�������P�.�V�52���!�W�_���.�����H̋S�$�Pj���Ѽ�Qd%�5�<6�>m�\���)�0bn˥n�~��*c���_\M�����]���f�6��ш�pe��b�b����B�s���<㊤@�%�z������O�a%�Z`��0q|����Xm.��,�[�{�7�,D�.Ӣ��rΣJ����Б���o/ݦ/�Όh@�0n�O{��m6�-�چ\��Y�8�������g�c��R���b��u	0=Kb�%1��m�w�^Z��)�#
�nW�����l�N�?���W��{h��~m��h��|esK{W����=)ĳ�F��8F��NgU13ii��2��L�\4�ç��*s=A]C��˜[�ъ��xkE�U�n�*ca'7�fo:���}pb����ƃ�1��ҝ��%y���~�&�,�(�s��:;���h�Z ^.�A͔��X�+��]w.�wE�|e��2�*��n�K�=�4BzI��a}ph<�Z{��r�N��S�����P�*�QV��\����r}�<�%�.���C~���)�/�@��,� ���тϨFRɩ�Q�w�v�+;���twy�ߏ��$S\cA�+�V �Ǩt����?�*��#�r�%��_;s)�g����H_bյ4��&2z��<�����bx��ٲ��	�mDJ��� ti6O�V��N���A�M[���3Jd*�4}�jJݧ4hn�Ds�?F찉����U)ٔ��VJ�>k�;S�	�b��BS�}/�L��^2�Ѳ�s�����`�Ƕ���/�Q���P��z��'��B�_p���FZũ�^N��L0���}���pWA���K�$����w�]�[$�~��苬��!�j#m�«ԊN"r��(ʌ����J�-��C!n�UgU��%�N���������I{�Ϻ���1&N�[q�Š�,���؀�?9�4/`p�L*�z��t5��V�M�6��M�KL�v`�o�D��qe/5�k�������<�Wb�(�e ]�a`�fcfD����_r�l���)��ܗc���_K���Q��`�Կ�p������&�z��&O�I��5�aD`߷��}< 0��}��p�[
��#������!�8K˞i�˃R����ߤ�E[[|��{�/ (�������p����Z�7��4D0s#*��cm�K� }�I-��ۗ��R��zY;Avv���1��&��"�~${�o�1��wg�s�����&� A�4��@X�?>Ս�;��vl���7+�d!jl�Y�Z�x���h�Ar�o�&���b�(�ʛ[��Ĩ@�$�+����*�4��8	*{,�d�}���$���%K�V]7Ao�6��$����L�JT�w�:�^��� \<1Tq��u*�ߜѸ�i��%:Nu�Ú'� D��';ZM���\�cz���x��3wv�2�������bȴՔ�bԂ�PF�A�ű�9x���m���f��2��p�:����Ѓ]~IN�T_�p7�˩!���@�u_�W��~� ���O&�6g���V[�*]�63��
H�������҂⥷ �� � ��M�B}<)@��[DGn�M��"3�^)�g�Қ�!��Xd��(���
SU���ǧ���q]K7ó��TKIːR�-�]��N"홷���C���q�Z���`߼�' �^ez@.!f)�9fi�~�{��7b�Ҭ�[��'�*��~�u������p��2
�+�)]�]-�+�@STHFq|ɬ�l�GwG�MP���M^����)"u�lE-��S�v�`]���?Y���I k}='��w� c�(O��N�y*y$�̄!/��Y5�lu)aͣ�k&z`%��e9�z]���_��+��i�R�a��{숇�:,���J��H�X�,�n��q��#g�Z�S��Q��/�.�q���P�w�_dyR�dh��l���w��'%OTs��?F��[A\�[p?�}���O@����-xW�zz5q�Pic�������#nfO��p�%C�RK"�v�_ �j����j�^0E4�P�z��k�	!�����Mk�|��ߡ�׍�פ
��l�D�;{�h%�3�׿v�j��e=��}�8fϸ�o�<Ȉq1$�'\�쯶��Z�F�O�i��.��Y�1{��v>C��k�o���`o�c�h��v#�>e٬�i��LHT��� ԊM"�K�7,^�;�X���s�()����G�WQ= ���q�\�����Rd��1pR$Gǭ�'�i�A��@b�8�qN��B����M�-��i�0�sc78�>��G��IQc�iG���I�>���!�m	L���E5�%}^��9[K^�&<6�;�B�fMK�u��]���J�0����,�}Ij�d#YѦ��F�RQ23��`�9i!Xߡ�t� *����?�n<g1Q2¤��˩�U8AQΐ�ol�D�5�Ǆ�r������ [`Z�@��e��K#�;��#1H��-���������x����TT3�Ƨ�X�?z��u���x�V���pg����$���Fc�&�>����\��J��[�[:�l!�p�O.��!��7ȁ����Pÿ�εxn��HozJ�E��H@cO�A`���m`}�ZE�6�#�͓Jǎ�S۹�8�滣�l[����9�7]=;���E�vI�/���v�7�Ϩ�'m?�	$f��\��d��ŵ�O%X����S�d�{{���f%��x�"�5��y�u�R��U�BV��!�L�(��-*�z��nrD�t��w7u4��a8^���U��sb���|��v���g��"db���Zw)�7�7�H�ha��l�$<��2]�Ƿ�}0�V���	��n9��Lm&����0��@�i!I�}0@����u����s�a��~k��tF��D���I�IP^@wsF�y��W��Ĩ�i����F ��O���� t&Ǐ�Kٹ�4�6�w@j'��v	��ѭq5�|�=���E-v+�C"s���j@W�o,��Eow��_��V�%�nt˹��o#�NpŤ'��om߆n����6�{0�E����}��`b���d��}eRH`��bW+���I�;������=kǑx_�i�C9m5�����Ph�����E������]l�|����l_�o�X���o�
۔���.ᯮ��S$)w���=�)�w���$%�ZM��c�w�����'�N�B�D��30j0\S�KD�w��Z������W��/�l�[˷?x�2� Nl�$���W6�5.ʈ�a�+��4(S�b���#_F�Yg"Bq��Q�r��G>�t/��{2��w�W=��`9�L�a�2���Q')��B��=�/'�O%�QXirjD��s�+FY/q��U�̵�X�d_>8	����Z�CA��
`��'�PG�4" ��~+ȯ6��3{i<�Pr��V��O�%�����&���0fX�:`Y��m6���[����S����2�/xN�ʹ;���,�H{�fۑK$��pl�ۛ�P&mCDf��R�\<�-F1GKQ�H;J��4��m��D��ӑ[�I�`_����߁��u�0�De���_#DZ�'��:�Q��2 M
vٲ���/SS�{D?m���v �oleg�(�C�5"���|�rs��R�b}���_w��9:Ғ��8�J�%K����������J^�b�����U�<��������_�Ŷkn�xy���� �5m�%�+$9��b�u� ����|���Jέ7�j��qx�\;�]���w�״Q�Ұ:��3A_��QQd��0�LQ��B[쁣�)[Yo,�ܼF��Y>~�ܕ�>�%fԄ�Ci��p	�w�������c��<q64�Q��&�����-&�X�u^]�m= ��xǘ�"�?��,�ܺvJttƮ�30R!��#r�Gs�ӫK�*���;�s�.���6�m��N׵'@�FC��IHֽ��]�bp��̳4i 84dDфuP^��E�*�"��4�z��x�|��d�M�zr�b���xȇ�N���00�և��I�_��}Z�~�.����	2`�j�'Z\�;{>��X,*~�n�WE���@��&�4��뚻M��Woݨ�ә��mzJ�#���=�Óֹ"�a��������j���w�DFn��F���5��\	�܃��ǯ����x`�����ٕ��7=v�>,�Hэ|��u�
Ԋ(�$�3<��xd��#8�iɾ"��70:�K�Bj�&��SMf��cU#mf�ň�i	U)m��)�Mdb���s���3��C9�@*pFL�f\爆�W<�豰��|�h�1$[j�TW'l�' D�_�V%|��8Z�W�ܙ�����@�
��^�W�膻{2����'SyHZ�hI��6�,go*����i6� ��1���j�6Z����c�C�[c��я85E�W�&+�!���PC�����#+S�뼍�Wq�䐽�\;s� o{�?�mX7��6ΠÄɟH� ��rw���s79�S�"��񫁺�B�����A%���-��,<豚A�_]��J�uf4�8�/�#��$g�@"|3��p�Ş�)+x&���:Y�~Ĵ�����gJg&��=G+C�f]v��.!�P,=q�աfQR�!xJ���@��(B3,�;y6�Y�}~�æ򘃳ߖ��zVtj$���lR�Q˔�,��ʚTM��\�½!��}��`J�h�H�X���[F�XݻO���zQ'�@�/i�D��˵b%@������e�r��g��68���%�E(p��lq�lGYLԱ��Upc� c���&�ϰ�GBk�S �o� E����ü�����a�t��{F9�exި,fH�(��@Pm�\#��Ag9���L�	�М���m�<ֻqs��W��d��o ����bMK���/���``2k�P>(��ߕ�d	�y�p�&���	��84�:��-qBq�iЊ'�Y8��@���Q������R-�u
|��{��,U@��S�)���jy���v!dO�d���:XH8�:�^�-ڤwb�<Q�B��_d�"!�����2�N�܋������m�T�<g���mM!��d��d<���a���>OR,��'�C�A�b�OG�S>yP�C}��e��D,X�7�`����M�vvW��bi���d^v=6����7� ��8��?$=�x��@��hp�Y'�������
��QD�� ��G��0�wFo�>`g��\�X���ǵ-g���DL|�hP�����������pp@a��g+X��j��%A��'�ʧ�������l�5lLҷ'�����?	����-E#��� |N������`�˄g�QQ�;:����:�E�Xu���}�arw.�]��U{��A@��!��6Fsd��p ���i�J�Z8�`a�"���1wZ}�)�LJ�I�N�k����k0��3��SJ̋��pǷ���`Mӟ��^�b��c�ߋ�"Bg�?�z���!�j� _�伵ٌ\t\C^�a���7��
j��Z��AO\F0�y�ߺ�t�5g��t��h/nV���\�ʄ����X^P�u�h�$�<{N��+���6�J�|OԂ߱�<�CY�K;�a���VHҤ.oVȈ���g�d@d+�t���=@���"bS&Ab�0Ajh$����Z��L(,���t*1 ��i�xf��9{����Y��E]�������W���g٦C�ksދ����9+"�5J��W�є�z}�B1@
=fA�T`���7��ۘ�S�H
c��M�ᴤ��NE�x�;����r%�4j�v��d�`C�
%���My����D_�W+�mE_0n��ʣ?K�/��
;���-�F����!enF�z\;E�m�_��P 49bD��G�T%�EI��j�M��45h6�ɑ�*�5�e���ZF��@��?�OoC ���ZK<�S-i�����; �ScS��ve�GkW�e�y]��yy��d���[F�-dfV�E+�~������^H�3R�K��Q�6�t� �Z�Iu�4�;0��K���]&��-��QďwEi�߹�<A�>����jN��9s^L_�x�ٺ�[#�p�2As��B� ��%%��e��+�q���L8�AG�RaM�V����Ϙh}��U{;+�؄���	�$]�0�ל�H�I=p9BmeC��	�||��\�\3�үVNE)c���9��/d��o� �9�KX���zb��tf��>�F��B��F#�5"�>�٠唗CL�2�嚘��~��o
��;P�J�6t��.���(�`�gs��K�ٻ�c�d�Z(� F�s#�OP����l�p_� ��ْ�t�rѳ:��׮���h�`����t���BW|�ܗ�i��{6o(�AP���:<��8�=�-�_�`bw���mY�P�u�J���"�EC���˿3���r�3v���J����\��nZ��v�4�)�wd1��_p��vIzVЀ�\W�O;n:d^�1b+k��懩�zTg�m�Ɉ�ИM��GZ���-��n�;�L����`�̋(��Q��w �vG�'9㰰Q\����u�x�7��Lt��������&���O���d��:T�z��ܝ�=����jխ��kTkd��|�����[�p`ϮU,��`�����胳�i�e3tb�����9�nh�K�{�PSL�O� ���&�����ݔՔӵ p+UGx�h�9�&~8�0��@~�c'�fVG�AR�+��F���n�~'�^�
�K�_6Z_x��Q��ѕv��_�����R[��P	_�"���r���z�;����_�(��׾I���p�sk$�3�O�z��%�#�(4�f$t�|l�K�s��M��6JQ�zŸ��.#ZQ�a���뿁�/����j���u�S�w�t޳o-��Y���Ǔ\�'"%d�|��DU^x���؏f���u�94P�'��|S�W	M�x;�I"����[�a��'jj��Z)�#1����Q�x5:�L��0�#1���!�	�ߜ���F�t�d��iל|�!_�,А����a@������)dYX$q��H+]W5wq`,�D��FP�;<������L���W�_r�w����0��/;+��x6�ȝ�L'��9t"�[^�.���;��?CIU4��5�^�����ao`1=t}����j@dMG^^J���9�Z���J���r��|�hs�����G Ō��E\�Gy�x�Q�LQ�hdqH���,z�M����2$0�R�o*�=���	�>���)&|ߟ��o��D�7�#s̃��#oF!6ڷ�.GJ�v]��2�+a^��ʸ��������N;Q�.�9�]�&0���LU���§X%�1�v��v���"k�E��@o���|�z����V1R�߿���'�ߍnA ��
nhG��ʦ3!M�|۵�P���`!���-*(��c�(3j
[�JN
-�Y�����&��&"�������&�����W�;���W����`�D4A �A72��֗�w��ƅl8!��0��@�ܩ������>p ^�5������[��(��������9�KX��o�E kE��.2F��4�AN��j�Q�*Ier^���?��G}_Q��F�r3�=�����R��ϴF�����+!��<�R�4~lKK^�*Mﱳ�\[�0C��B�g3�\�b��4b���u��+��R�!�>�Zy�T�R�d�^O�t$.�K�@�[�<2�w�����#�L�-E\�/��3jɵ����2�jҺ/�/�[����@� �K |�=�)����q|��Jk�x�"��:��ⴙ\߳���/�_ W�򅤃�zzş�j�`[r�nV��K~ZL�������Y���e侥�����$�j��ns0G ��?����\���=!<z��{T#sEq�t�D��t[ wo�C\����;Uƴh��Z�@-�j�9��3��u"B=9�}u�Wd��R�� 2{����ʺ*�'I|_u�
��7��g��迅#��'�L�4|~0\����e5�g�e}�4��c��a��{1
�*�>-]v��n�R=p�든�h�X[���_��K��ˀ�^��-fH1�ۂW[]�Z	?Q����X�<[���;�d�^3�_S�e��qY��wz���������0i�w��`�g�;T���3z�8G>^>��`\yn�����X獟��sM='�ܭP��{���Ӫ���S˿q���@/��8�C�D��i��%R�Mg�	R~�¡.��%�n[.a�wj�s��Bv?�C�g2h��[VM�d�0P��Z�fFCv˶�뮀����E���;,@��/���y8����A��ʤ6������ Bj�{ׯA�TVF�|�J�F�2_��&ym�o�T'��ܴ:��p��keŇU��DX���"�7'��h	��t)�c��Sy��R7'<|�xć�"{h���X	�e������΅?�FN�׬ �C��1i~�	5�Z�ft�Wa5ۆ�#�/���@qv�8u�2�h���t�)�i�~��W��I�*�p�\����Gb�6;�\��m?F��H�Y�h�ٔS��	:�@N��^�>�� zl���u3d�ɰ@� ½f��S8d#-R�]f{����6�/(jbͧ��i���i]�2� �*���S�݂<���5�m�����V120��S�ݻM��R��	u��]�j�"̸ V+�.��w�XפtL�\w�;�����D=%�_e0`� ��wJ����*,c�b��q����LSV�i�<����odMCg�-��5a���ʣ��7���\�SV�|���D��`��p�J��]���Z��;�N�~-o�)w���d~�a'���b���=�0@Pt(��p:�����b�T�m8U�ϳ����.HVv&o��PL�I醝DI��R��Y[���{��*���bg�D�.��'X���{�
�n��u0v�줣G����5�N?7��!����V�( �;��vǵ��.��1G�h�J��Z6�<�jSד��ғ�lS�+C���J$����2�ß�3X�e�=���0CG`�S�o?��������t��J�Wv-R�g�]r��'��A��6Eih� 	�B/mky7�����_?UG��(�j�.ǥ[���2��S�2cx�rކ�X�Q�*�Y���odM�KYU�>#au��onO�8��=E�s�j~
��:�F�V�Pn6��f�y��IЯ=��e��i��-'��h���@��h�wE"XA[��t�/�'�箺Ȉ����5�Pa E�H�gNF������	���%?��i�1^�g�]����YtZ]�Z,"�aP� p��W��S�KpGxR�Z+��#x��v��A�<��R~���-�'���o��k��J����$o���)�}�Т������r�o)���g���I9!ᛜՒtk�}Ȋ�z�%@R�ҫ�'EKw/��O�C��4��Y�$����H�6��c�!�a=oz�+[��5	��:�1�������N�#�q�Q�3>z=�,>ѕ2�%��˯����e�)['��$f��M4��ɓ�pM��̞��~��/��BO_w�5uP�o�㪢�����仨0��c�V����Or8x`A�aտ{�2T,dث�먪���X2E���R��8���(�y���yP�JI��uef �w�W"�6��$b
Kh��luT�#Y�
m�zY��M��SMN.�/3��z:����I��ETn��9�e��U��l�ZL�(+i��^&��$wv�x������,�P (��ʥ?�-R�&;�k%-������&-�+?�0�E-�����2�XX�[5�T��+��-t��5I�ҥ^���zwpq@Eo���A����˙^�sʝy�v;��:���E�r�(���RwYS���v�..^�f�.��<�0��?AO�Ę���������4�N�&a�>�mփNy}#Ҿ(`��D������mP�M����n�Y��3��`T��1��n�.����V�)��c�؛�TCaw�- ��&�5��# a	ڋͮ�G>q]ȇ�M�F��#��W�}rQM��	-���phՙ��J1��dXۮP�DSqO"j}�W֥:1Y�mp�}�t�����VJ�Vҥ+!�.�+;���\Om������|RK3RZI��P��}l��	9�o�����2�U�Nb3�mم�������\赜�ݹ{k6�ü��Ιj}��S��߶�q���a�P?�8� �$�W�����PU���7F`#��v�o��FqZ17#̇�Oe�1b����%�v@���������Q���c�N�q�i����=�ʻM��:��`>Z��f?�NLJ�2|I���|�ݡٛ�'��~`�*6v}�0�Oٍ!�
zEǓC�Ź��r"��1�R�wm0���+
ӟ�6�ǖI�����1���E�b�+��R�B�4�����g|'�?�X���I�C{�:��.���l����iӸ�D$�X�?2O|a����q9��0K������*?��ʒ���;&��r���E�Fk7�{��&�[-R��|8��0"O�V���5�#�.l�l�w��X ,�a�\]�RY����F�o��~����*3����{��cj�(�,����ё�� ����"4��=�&��VÃ��D.��''\��;�*Ƴ{��`�Pa�X���NbK�����h���4���c�n���������x�έ�����U3}m
g��o���g�Ҿ]�BK +x��A@��U�!���˂��������2����=Q1k�?�]�q(j��iu[)�����H�$����_f�܃z|�� 	ŗW�����Xm�F��`P�GI���S�$Ț��Ŀ��4�O�u���qC%��#�]!�VZ
�C�*��\�4
��cQ�$}�\�"�,�?{�a,���,�_
��a2#�~���E��K�vt�ȁg���@a��Ȁ�������t���=��:I1��=w4���f-��aE3�wUJ�8L�Dɴ�v���fu��$���n%P=��`���_��f}�U�y��:ŷ'���[��:.��C5�X9K��@�,h>�Χi�"*�{6~�_�s���
�ׄ���Yx��h����i񀔂0�o��Vń��0�*�['�4C���l�b�ƥ�U��|�Т
Ĭ�
������Q���VH�!Ǖ����y�zՁf}4Rz�v�]�ij��ԥE���n�r����!>��ͽ4�R�
�]����Q��Uӄٖ<Z�7T�ĵ*�h��(�}F��J�w��h%�oӺU57./�f�>2�ͱ[�u�"���;�l�$�����I����[���R]|>��$5�ܼ����<d���r�q�t |u�~��д���ur~(q�yu�Sc�G>�>NF3Q���u�G�h1M�w7@����۸E҅��5��h�Ņ�b/�������	c>���G �Kk�<ݥk|�抇\=iz̄���6ު~T���*J�Zwg�;�	�,a�D7cі����

w~x�ĩ�ԬF���)���܈�d�.�:���!A'1�,�fz@��v��f�g�T��Oe�x�hF�S�
��*L�i��� 5I�*}��vy���t�c)�GJK	�7�xF&f��	�z%�Q��#���L���1ѽ-��+űP�~8�N�j�|��?l�	2���AN��N��ڵ.�+��i�i̓�3�+���x��4�
�&P��^V�o���������O$*�Ii���"�����i`\=�9|4hF:b�Bc�d�q�H�O��E���� jH�Oй���n9�t� PLF���B��E�"��6���W!���X[�vvv��n��1�2u7qPq�x�qb ��w�Uq�T Z��(��4SXFT�/���lt��:G��;{p�aZ���������ڻ�͸��$Vk0�{�ES.�u-�Ŏ�q�n�i��$�ˣo�I;f�Y�1%�࣪Et�m�ώ�X<��}���� �����Hg�/]H5���Oe2襁�=+��gu�?&:�XC�G��v���%-O�N=��`;(
�����n#0��U�!8��1��[���CM�B��Gov�>d FÙ
��Ěa�|�*į����A�>E��Hj�g@W�u�>)�ۻ4�"*��a%A�ʟ�� 㺤<% �c�q#qb�m�����'"����%&�Ds���T��Жv��3�>��ؚW�V[f&�0Wb�L�\Ϊ}f�QC�"~��$�m���*pJ�U�Y���ط98=�l��;vo
9'�t�;�,p��h�.�
+�ܪ�i�h�����I|խwT+m$���oD����I;I�]aD&S��� ����~`A:C	�u��O�4G�[���H-: �V
��Bd��������̒�U���]�9�S
i��ST�o}xrl*>8J1��z�J �����)?g͑���B!�0���6��R�)����Ll�����-4�"��C�b���?�t�+[{/���ƭ��I}�>~�p�D����.����d���I�Sx���S��ᔼ� �䀣�ڿ��b������%�aW3侅Qk�}!~p���Yo��p�zB���k�����.�P_Hp|֌��&�
����Z�����5���5v��Bi��	���X�Ayv����Ǌ4��P�����H��V��t�F#2�?��Z�&�'���3a�c��F}_?��l@	'�y�����ԉ��a|P��TL���x3�7�qn�%�#���\���S�kAU��?G���KF�Ӑ��'�4��<hƤ�bi��M���>A1����,X�"+�_���1u�quJ%�u�����}�S��q�����Uk�E-��j�Z]�d�K�JM�,n�\�����q�݁e|[�ג�v�=��1m��S/O���KI6zf�d��}	���rf	��(��k�O��{�*dtǊ���z����+���Q��v*�!)� �F�<�x��Q.���Aé 秎��+si��	-�asu�g˼�u$�S�Ć�O��%܇8��z�Π`�f��'J�sK	]����S-��Q��fGQ&�edM��Q���?,]{5�y��(|0��
?9_�n�=.~1z��dJ���㨅W~��m�j�^M "�\�$
Ԣ�m.�7�=���-��A�������![�L@Y��x���\�N��
����Pa�xd��uE��}t���7|�X�J8�~��ʬ2���Y��5Mv��T���*C�@K�:T�m$�q�%a��¡R%�����4�Rwp���g��)ƌ3J{]�r~8�7��?)ż�8.E�<T�,7}[�4�~�G�
�#��� \<zݛ�>y]���ʓs�gU���o(�g~j5��:^��u�)��2���8H���M?v� ơ��WO�Wf��+lԓ�?�Rt������5V����j����*�I{m���n�bn������C�
_�} ���#)��ԏ����&+V�	���>���K1�~=*jus��L������?�"��>�a.V6&O�q��}�VQ��A<DB�w���F�kz�.�e�=,4�;.��@X1܄����m�vP,��%���FJ�z�?G��~��ӡ�����!5�a��iy�^����ǅl4�YƏlw��%o�`�����������)$ݖ�<q�İäZ��.��^��ࠉ�g�B��g��I�	Qw�X`O�F!o(	�B5N�?,́�����..r�3����7;����!q��#{<��d�fkG$�����Զ���6quQ�a-�[�w����V�*��hI���~���?�������=i��NDP���RÊ�4-��}Oe��*�@͐���=L2!Y�k����A����[ܙ�/b��7	�W�ω�ض\��4��늛�=^`��狌
MeI\��@�7E�#]��3�pרn-�K�Z�#�~����Z8�ig,Q�-Mv���%��"sG�~,T�s+x�W�q �F8m�}t��]�D�e���e��d<���u=�d6 �"N=� bנ��i��D��Y��>�aFµ%SNS���E4D�Y��s�
�����f�	j�l�ɨ7�@F�>��bT;�!Xu�4�2&�a#ZP@��c�%�1�^�o�O�K!{�M�w�g7rcϭ�,] ���9�����n�#�ŏ�r��$즙k@(n=�~>'J���@�z��@�ķZ���
=�KΣl`��a|�x�(�����pJ���%��0,LB���}���v}��^M��ԦdUh�R�@�l��cYڼ��D\�Ճk/,�j�ֳ���s@�=C1q�ߟ@V}�$
QC��uǂܮ�Ȼ{��_,��n5[t�r4�G��+p���&v��Mް�8D;&ݙ�<.i�\����͆��C�b�E��X���H��ȸ�iD�4�U=\_�IDn�y12�#��y]�щTĻ4�m�<�ZTB���w�^�D2,n�c�|�A�@t�n�.3��v�A��P��~=X��+�n��W�)j��X��9�v��y�m�ɻ��X��-��p�y����*h��i����J�x��g�ڒȭ�I�V�n_�hK�������i�.J �yZ���F&�0U�0Ȭ2HU��:��7!��?�a�K�)�!�����c��+p�|4����j����wC�������m�[,h�ǚq��A��aJ�$P�k��û��Z^�n��~�8���B�9Y��ZdD�V��S(�@��Dw�=,z�ʪ[�k�0$r��\.$��$f��(��O�Zz�'�. ���y�0�m8�h0����@6���x���I�+C����Cg��i���(*Eatg�]�*�VS0�l����E���4��m>��p����$�p��u�h����kNX�k�p�]'�ee&��j��fv���b��S
���2xL���p����2��)��5K��c��31$�j�c-���f���lgc��� ��Q�~�7�8)u3�T^�$!q���R����m��X�x�V��1?7D����TB��U>��P������i%������W��l[�H�}�����;�bi�Z�g_��D���q�Ufj4��n��F����Sv�h�h� ��WM��x�����"� IK�M)|�}��c�)�RƮYI�	�"w}ɲ�0�,o�߯��K��� �FD�غ-�����Hx��1��=?J�^8V5�{p��|a�p��Ct!7:�� 
������u��@��,��GOU\nT&j�خ�lV���ާ�ϔuD��H�v��\~ڽ�0<�nF��3I�+ⱛ�3V��/��xNw�Xi�4֯#�6����!?|��]�POWE��u�y�W�<�ح����-�y:�)��إ/���.����Cs��
+D�a��oڴ$�җ>?I�{��^����o����Ѿ���A�vw^��t�h�X-��ƌ�;!��DԘ��11��6-;zJug�H���L����Y�q7L���G
n�H��X$���A'�aT7o��0�O�����e���ޫ�$a��'������v�pz-�=��������+�%��>zU��=��>�ěZAc���;��p<|P��ᥕ�7�{��3�Q+�?��ˠ����!Os������ ����������Ά�ŭ/���M�جU��ID!á�>g\}�";���a�	�k� �(bj����@U�o$��΅"ri��Փ���S��;ſ!������s�Ȍ X���M�N�\�����F]�zE���1v*r�z����~h��\���[޶W�䑮����7H��vCeۏ�kĂ,�X'�}T�+�h�����n��]DW~/�+����V�iq�T��o��7]�6�`�-�_MZ��V|8O��s�6!�Nf��k�j�Ƭ��cR�Q8%�&uDx��q��������x3bfRr�%�얒��� 8��o]��R�ԃ���o�����P��O��loec|���3����!த�q
s�k����	�/L�0���Ļ4�g���K"-ϗS�&CM �E��x_ޑj丿2[ح�� �E.�&Y�NO���a���� ��U��]�����POA�'�ԛ��+8._�T��t-��Gv����V�%btk6AÀ����b��ί���Nѕ���
ϊl�1{d'~�1:ۺH�`I`+r�	n����>xc��K�nK\����n�<��p+=�ϣMܨ +�
�����2����/�������b�!�q��${O�I����'�����OX��ߞQ�ŏO��Ad�)��/,ѵ8�Q2�+e	�����`ޑ���Mf˅%�*}D��0���ч��J<���p�v��n^�	Cp��DhԠó5K>^*�zw鵶;6����w�羚o��;�(hW�j��Vx@z0:��������48��a|^p%�)��A�.\��8w��-~rvQôhJ��H�9��l��1��G#���v(d%����R��ǚt*v4MVp@���/Su' ���E��o�@���:���Q[x��4�{a�B�j�de�²?/��K�"��$q�s�c���^�������X�����*4y�!���y�#V�5�v�":D'�u���33�>�.b���?Uq��x/�zB��(�tA�"��aF�ozT"uV������9+��}\�"�{��d�.�����@�X�E�������N��l�˂���Q%���C�D���sL�d�`��������C�1�����H0c���tJ]�����_����D-�z��M�["h�aǢmGLiF�O'����+
��s?ֽ��I@��'�[����Q��R7�#���.�O��+��E:f��9������Tq
��g��V]��D�8�_�6�e]�$Ly
f�<�m��i�>e��.���$Ї���?U4EA�K��隸����\�%�n���m�i�7 `�&�<���O �f���r�fχ�"jZ�F�]���e�� ��$���$%�LBâ05���0UΈ)o
��ׇ�DXt��<VZ��-2��,��@�D��y���r��"��#���[a����Øk�{���5��B������j�*���ʭ��3X��DG�'rj���V$�7V�d�E ں9|��c�S6�����C�\4�=[:�Pޔ$E��?��p��]�kZ�H����e`~z�v�Y�6z|�M�����/\
���g� {�X\ �	�z?�MGR��J^��E�*F�t�X�{S5�% �����Y���3�����u�u��	�8p�χ`�e�<U��g[�,_A�E1�*#}=H���h��eX<�����I؂���ݍ�I�]f
��F h
iX���>�y��N)=�}�%�����U��jخU r�y*!L�����7F9�ޗ�|iئ�
�m����	�B�:w���EF�'/+#'ڋk뜜+�"8ΤP����Y�"�Z_�$;�(��2 ��������an��\2���N'�c�_,����������t��3a��̍�j��6^h��1Bz���ѾѮ ���'BFp
Dn`D�]E�g�����M-k����R��~�hV�F�ߧAaX��]9�o�g�%^o���'<��m���p}�?ި���^��,͑g�^G�FU��@�z4yɗ����X|2�:YR\��Os���(��y6��Eh�!O�D��<k\!�k�Y#|�%����t�B(;^���3��_<�T���M�<�s	,=x�?1/�hgV:%s�n�uʣZ��G=�����!0(�J^�uU�ϗ���~d���(,Fc4q�Eku��[BĒ�-�"�~:��1d�����X��X`�1�����K����������&{�-��8��p�;;����j�(-'1q1" ��^bv�>���&�f0�L�j����W��%�	grP���.<c���;�?x|�g����ć8��&�]��	��F5��;�o_��X1�A�ͩM�4k��>�!������!�Z|�H��!v�p|��u�-�2��� C�X�^j��빎T�wĳ��ؘ.�mWx�j��h�u�}�̓�&�H
(��b�H 9��|�V6�{�J��D��^o��[5/���'E���XN56����#�2{��h9q�c�n����mI[���S�p�1�ɔKZ��Uf���R��8S8c%۟3'?|� /�lL��B��i��˪��>�Q�� �5���'�G)��-��2��~�$8�`��-��k#����q�(v9����.(��;�6��^���PD�H�5�i�/���+��'q(%p۩��
"}]�%����Y�Sv��`��B�M�-"����x6��1K%p��$�=�┤[�r��n�:���_R�M4���EH�3����!�J������߶�(�pƖņ_z>�Qt9�7&/�a�;�"�-9'��d�C=2��':�kp����-,}B�tC'��^ (�\�p��<ٯ�{'�;�����Cη�j�>��\ ���
�.CF�z������s�c�ux���߭{�)����4��:�t�	2�B����;МL�����<�W^)M��s������A���@SjN�ʢ�?u�G빊�H�:(�]�
��3��1W��>D�O��6�Kc ���y��ؖ����h�ꖆ�t�cߍ8/�4��!ԣɆ2qY��ib̂ٹ�����H/,^�(SK�cQ�Ce�EG7lʰf�EX�����Y�JfrX��2_o�<�����}��ݝ���13�Gt,��#"Rv=��4$N[�v�tF<���p�_�?i���Պ��e��*v��:ɾ�O-(�v�$S���#O��I�;�ǅ�4M:� x��[$TѰ�~y���l6����x�RyпV]�}_���S��!��I� ;����|E��n�����k�p'���]�g�΋3~K�O#�Ȗ�S F>P����������m�L��S���/(�����6I�L�g�=~��� ��L|�oHD�����!n%� ��P����зZh���DS1�r�YJZK�"J��������t�:��S���-	{�A��{��w�d�c+y*HU��q�1�^�5k��i�"�q�$�Ui�3����X��F�� �+� Ȯ��.lc�gIgb
�3a�O$�ҙaH&KZz���q��&���uܗ0��y(1, N��/�͙{����0����HVj4���s����
�B�P���7
�"�l��x.�)|�=��-a�B�R]���%��*��j{�b��O��4m�M�#[����(.I�	Md~5���?F٧UK-eX� ���8�,v:&�^�ՀHJP�<t�\ݚ,�e���H*�� �Q�)Uͧ����R7�]`������۫���z��i�)>��w��z{j]+�ē�풆(}�%�~�lw�y)a�,!�F�����̞��Xf+�Ŏd��|�\�F&n6���+Kz�L q�l�x=���r	���S�W�n�}�!�L a<w<ȼ<.�����}C T.�{�׏L�h����`�'U�t�}��I�W�w~&r��O�z�����]rB��TCҠ�d���$�#���u�p�w��Ö�
)>�g��i��d�sd������ܺ=dɥS�߹u� ]\���a˫����o�l�xI�"�����1�ʢ�`�k��r�=�^-ƅ��E��{����a�r�����{4y�������}�*���-IkV�Q�T���!է�-JW���	4�����grK�H�!��{�褵f.}@��q;�yf_kּ���I
hhS%�Ь�o�3X_B��8$�q^�-���7��1�����K�]��ǝ�i���p5�+�6��W|woط�%�M�>��?,�M�ڳ���
&oA�:�����0�OMr��l����B�a)oU���GG$�!� P�TR�'B����
�a!sٹ^ �T��˻.����r���ɣ��n�g'S1�rv�{z��d*{��b[�r&�/qPu$�_�(�`���G����y�J= �f���Ѹ:6&U0�{�aϷ���K�Wm-�T=ag`=���U{ϟ�5���k�f���_{ơ��jLÔ�?"-�`�7���zp2��a����+�'���
`���b{�p5={�I^Z��+�x#d.},������LKg����S�`��oӎ�����_�?o Jl��3���Ƒ�V7d0�q��
����n@�CRڙIDZ���ce�{�ͺK�*xXaF�^@m��̸k��Xj�mö8GE��nF��*���g��5[ۊ���k�S�d����=��h`}A��I�eP�}&g;���֘�σUa�:o;�F�����x��.H����x�̓�����&�(����b9��, h'�6�~�m�`��I�0��^�>,��@���-F��ޜ��9���s=,���ň���-�ÀmSC%f�������HO��.֋��E��T��j&x��q*_�풾P�E����y��q`/��"&ka+`mf+�t�x�����Ӛ}gC=:���3� ]�]@D=;6��M٣��ԟ�fK [�b|��^�1���Ӎ������%���}%9iU��Z[��8�g��>\z����v?�����4l���5��:qw}A%��2�;?-�۸w5ޅ-�hp`TЇ�����߿�������z\1�G����(���qp�{378��:7A��j��Kst��y�z�@�5�4�����uF�~��D�j\;�jڪ}�M�r�
�Ra�ci\���lGɃ}Dw	nQ����	����J��r�L��'������]��:G���J�2����/X-��5���NZ�(-�yc'T���m�0�ڳ�K�RH-�Է@�@>�Y�7�Z|��@e��I��e������v��P�ye7�J��М��	c�#��E��Q
aN�F��1C��W��Ǡ:G���� �)�2���[6���ѭ��z*rZ����Pʤq�c+&�ǕșEݫ�B�^E��b�á�j�8n�4�Fw�`�ʺo��?�AZL�S����������_��������DB�b��Jݡ,?q7LL�GWs/��a�v���+0���[u;�_����\����6�*?�m�p�U���������Nx�=`���k��p/N@A�T5I�V^��Х$�(��E���L��� cz�X��B8���-QJITy��ܜ �G���n!�|�m���*ڽ��/PP�� �0�~,�h�"��p��9��<X"oV��e,o�q1��!A٧0�m.N&)���w9ԁ��"xn���=p1➸�n���_ɾ�����gA�h�qU��|��;��Iƍ�-�љ�b��k��E��!��L�����2)rW"RBU"
�SMW���?�y+]02�y�{L,)i�g�(�J]��K����LC�������S���Q�F�+�i��2�vV��%�~a=�T�%B�_�d��#U�R?��e��2ៃ��jJt�g�`��v�֊M�Ъ��M���x���A�Y.�JS���Q`�m�X��ؓł���v�ɠ�x�8[�G��<݈ΰ���9�G��&햖tz�<���xi�B{th���O8��֑��.d��=Vc.��h��Pt�	�!���W��E�I�P����S���<6��NW��������z �2l�_�� f䙖#�΍����`c�����J�v����1���;�Lr,����">�L r2���Ka��bQ�NA���.FZ;��@72`&��5��E2��D�̽k�2B �������d?�n*�S��1�|�V6J�`}f��Xe�� ID�>�+
6|.gH��T�L�E�\�����ޓsq�-/�?�a�3�ʏ�j��%ӡ5oE6MH����]h�~c����u�k��=���ae�<4��}�(���I�[�Zp�Ҿu����Q��QRa9$�����r!o~~��FY蘏=ShP�h�ۉ� K�&���C\���ː�~�C�*��|O�ROdϓ��D(�� �|Y���(;_�IND�l�����5Z�-`����(���pQob�)��̔Z3*��V"�&���aq-%<�M�/�7�ȃA[D��J�6J�.d�S��������r�A_w�.������;���o���8�-gW��aWf��ҋ�x����F�γ��?H�vdZC�T(��3]�g��-[��}R�?�ڟ�G�;�땾f���m[��b���-�39J�a�%~5�ޱ*x�4�tH�Na&�\���6L5�[���`�nZv����
G!��]�� ��/��<��n_��J{��
�oeRB��Ù��B�ۡ��wn7Xދ�0m��̩�T_���������byrb�k��Ƭ�����*�T[��Gj�/HFݼha��0���D`�P \�3�]bh�`+��S�uR��L8��W�.��k�2Ԟ5@
���(�(΂�l��؛��c�C�<�m� E|��#t���ܻ��iFEO�t�|���݇jҌ6�b��~�3�Aa�Z�n��p�@jV�)_�l��S��(���wf����&_M�L�����aT���n���
\tԪ	̋�����]�Gj1�<�)��T`7�����|��4@����N;�,sg�V���7��A79
U�/��u�*���v�C��i�G	s��1ǌB�b��~�X0�q��9�5B��(^b1�~~��?�ev��9�Kh
�0
�N��� .r�F��w�&S��d ����z$���	p�ֻI,H|���9B��M�-�w��C���*qr~y'g6�c��m�s2������`��&٫2�%=|���xk�a��k?�� �H�oQ�I۪�|�d�&L!_��iGu�IC�H5�j���#�&2�=w��_y1s4�7L�M�Z���#�z7�����p�U����A4�����@
���!�����&t�\ә,v~\��CS�>M�_U�-e7���X̎�����8I�	>��H�;��R+�N�s�<���gǭZ���20*�`��#ڝ�<���'U�,?N��)#?6a{?N��b3>ށ΂�M����|-����I�W��&��,�qߣr����t�PV;��F��R��q�v]�j���rϧ�+1�Pg�//9����)�m*8cr*sz��Ɍ+��Tٟ��d}��Z�Kk���W%����)q���Ⅰ�,��Rz�*nM�]]�RGi�Ռ[G�Κw�8���EuS)sqv��E��Y>���߾O�n�!�y�1�i����k�B��"A&�-A�rh�oy�^���"t\�'���1�-
��$	Hí֢�V�O`�V���Fv�Ȫ2�|K&j����}[��3��Mո^y�X����iש���5�a��~�B�^D��Hc3�9l�����!��^���'l"�d�;�]��s��bL��}PXe/���_�³$�v.�Y`,H�˽�N�����w˻��"�D�Ͽ�u-I"�,�H�$t��S��9��q��df�|������2���S�l��pO�Ӈ/?w9E�l%�kN��ؗO����岜OCl����?�gmx���h��e�"�����{��A3����^m��b�usD����瓤�[�"�6�V'�E6�'�פ�U�p��NΦn���`p���j�X��Ir��@疍^qu�b��[<KrR�2�aJmi�v�;
)���O���("W	�1(�c�<�_���`�O��_������J@Y��r��]S:C0d�j�:�戴�6�$����d��PC~ԛ���Tl�K;�&�7�6p[�+�gmr'�"�n�b�q)�1"�׹�	
�)���Y�Y�@��}P<xp�ʱ�mѿ��놩��XYn).��)�ۺdIT�b�[�rk2�A�$�7�KL��d�F7�
����&��(�������ҽ�zJ�B���zI�O����~d�K�`9b�k�kH�Kɹ��v�h�[rkW���������;]�n@ƃ�#Qoj����S2.�ﱐU?�*ȝ�i����Fn��5����e�'4��G��� �U�e{�L?Gc�Oo�g�K�EV4�sЪ�Y�[�mPc����Ȃ�s�'a>���Һ�1ieX��H���W�z�hN�|Lٻ���L����-�y(#=|��q�L��t��3mE���@m�/�NCy��ˑp�������3��{c����6O��sE_���h����w�-¢�j�.t�� n�U��`�ʬ�ͻ�ӰXQ�3�Y�m��z0c��i�C�X�
���z
��q�7+�����92&����ҹFl{�����$��v>��.����}�#MsBV��o��/g�%�����|qJ����t/Ϭ����8��r�˽��bX<�
�X$�"=�16��
��+ֲb[>��zv���I�?IGE�{��^2
ud���-���'���G��?�Z2!�8/S�I�����<�UDi����x%Πuda�%�"��x���s)dc��_(!����]�(������&i���v�Y��w��@<�͛	'�d�>�y=6t��֌J��i1��i��= 4B]�����.�JC�e��Z���Grk,�܆�ٔ�\u��F+��p�䫴g2V��G�U�
W��δj�r���9�m��g҈G���ˮ���+o���~*�!���f�J9�O\{}�o�Y[~�NI4(?� U�/=��ހꩡ��\����A����g�v2�tXբS �ol(G�\�0­u�L(��>o~&�?f��F-��}��'`�p<�����no���hM�� ��#�����99�@��'��*���ƒg~��v�,ű>�cC����{\Am�&�u�����=3k���'���F�43?̈́A�L���w6e����{���Rr�0Eԇ��$���&*�xp�{4���� HQY���sGd�R1]��ק����� �Y�Ʌ��&�u	�é9􄷍��t�KѩDn8�����q�X�~�+nw���������LauoCLٓ	w�)�?ZZ�҃�q	1y"��h�k�ٟ�~"�����<9��J2J��<*���>��&	癲�bPt�5y
']�9����u���S}����<� �X|$��'�Qn+	�� t9�&a	���t�|��OH�����I÷�@�qG��3�����S"�c.oZ�X��1�Ae$�f6����^w�&�H����"#������+*�q7�QT
D<��C"��!3��.F�E9;M����O�{��o��I�%Â@���d#���	���*�*�Ǣ���������B�{�0y�C��B2m�j���E�h�p�ؖ"������z�'�K��FU��8�9��S�� ���9B���~{Q�7:r�t����Ze@O64��b�Ikהϵ�%�@��iM�ȇ�-l���Q���7��Ȑ-N��J+1-Ҿx/��\H����-��}��^���V���g�¦.s��$l�������4�"���R���������e!ڠ�
�\�Q
Z��O�F����/�����=�pO�Y�Z����=y�j[\��r��̓�G��-U�ewP�5{�|9���W��W��&�egup;�m�#E��S�/\���\�>��=����,�!�$�">M�I���3?�,��b�Ƿm������JV:o�G��`ns�@y�f&3��Kg�:��j���2<X�~y���%һG��S�kΠ���\-_�d��s&�%o�r�5���}�1�v
dNu?�S�Z��uT�T�"QZBk���Fڈw�q�����B#G|��h �] y�'y( �#2�P�'M&El1���ƙ� xG�z�
H&�tI���@��:�aߊ�%�)1el��V�g��W��1"�l�nD��;}X,�4�|0��� J<A�ڎ�gI �b�C
�	�Ri�
pM9-��$G7\����iƦ���9(�q6x�7]>JV���yY��1��E�ZD0�>���#h�?	
�	n��[��E�(A��֕4��y}̚'��ҵ���k`�Cz^��$�Q�T����{ I�Q}��a�{�K2DRJ���5SaI��ת2��(#����,����̎��K[I>�e�ò����J�$��}G�gI�3�<���<{o���<Z�:#Xj!d���T�(z�x����;t���VR��hc������qr�0ݩ���߅d�L�w�\�+H�vz���l���4�HK�j��땳��L�"���fb���s���:��E�(�)��f�Kd�����t��UJ��M/�����fO��N�9A�*�)����R�IH�^Nt�Ҩ���� ̫�!R�ߎ�T����������\�#�2u�q�7�\�Rb�����m������u�pP��G�8�q�-�_&��%�_��em�i�C�	a�\�5ĲID�dk���CLJM�����չ�|���Ԓ|leӺ��!�[4�J���7K��l䁤�y>�	>3	҈A*/٨�-�s�w|𩔰��[w���ʷxʜ�y0j�N�%�U�B�b���D-2�K�g�<T���6b�9X�c��'`"��'i�D�pI��)���aT7˩Dg�����Q�m���=90.�}`a���eO�W���Wq.�H2Q輟�������N~a�>EV��	��v����b�8Z�x,�g[�]���,�/�1>¥���!P�*�9�B��0����� �|�%C_Κ���e�4���йW�?�q�->�8�}X,&I�I3[4V��/�Z���w���.ۖ�����~���[�
 hy�2ɼ5VQ�����6�߯� 9���_:忬����zJOg�OPC��nl���Ȃ����$zw��*⡐]�3�[��
���6�1�� ����^���"tS((ב����;��G�����S7E�.���Lg��r��C��Ӫ��S˒6{�� ��1%��Kb��S���#�	�l@�x������w �qv%���^Af�u-�h�i�p�+h\m�� ��.2�]�b��y��'oR�LhBz�S��VH�?�����f���<a���a���������y�t�S�������u�Y>�L��U5pQ��Ѵ9 	w!q&To������kf�x씞�����Ҝ�xGNO��/����QZ<�H���RgsRd{~ #Q3*7f:Ry����6i��!�g�:�w�02��(-��@�kWJ�2Y�_P�R�Z�%��E��C�Y���@W+d�&@A�US�۴���>��cGlF�)��Z���n�6��>�\��pAi> q*���\It��sۑ��M�@s2P���d����e�Yg��opg9�B�]�A�o*ᷭA�ޗ}�$e97��q8�l��{�$5��?��^`u�ߙEK��l����(
��,���Pix�ײ�â��5��;��
�
� L *CȄ����������$���CTM�|Q�ڟ�L�{�Z|��������x��MǍ�C6�n�A���?l&���[�nQ#�56'���hI��l��+�OUE��kջ� ��c���P�M/��l���/��U�A|V��dT����Q��#�=�����
q"xqF,��.��Q,�#=i�5x�&�F���e���s�@��Xrv-�p�U�$-h���l0����b���'bS��f8�.e?d~3�og���r��J��Q
�R珊U�{Z����53dj�;)��oW��O����}��Q1��T	J��i���i�V'�%�G(�{cYK�0$��
B�����$�ë�s�@v����H���vjL.�*���8���0�i�����XvV9�4�_���~��fRrf��6~+> �N�/	Ǿ��:�|�&��YaҒ�i]@uޚ�B��)�صL�R�8�!K¿��R���Uu)�=1,�\#{��Ƒ�_ܧ�-s���&���>����Љ���cZɼ�� F��C%� ��&Nʹ��Ʒ�dm|VI�8V�M��n��a��E˯�9��W�pr}�/�y��a��2��#*
��,���<]�Е}:g=8�iw�g���WZ����-�s2(@"̃IF�m7��m��ʸǛ`�nP���UV�X�ņ���u[Y2�=i?�ί�����UЌ�`�с	w>�.��G��@�s���̶�_�=,����vm�~�Ym��铟��E��
q�V�C����#y:<W��e��B���kxX����<'�L����
+��]����HJ�ƅf�{z�O�mD3A���odd��h���{���;U)��v��z�#�$��.�r�_ TZ<�w�%g�� M{.���+-�����A`��2��#>�V���������ړK��Jz���Yb*���s�N>rP4=�-�;Щ��g�@�^G�w*�]� !/���Ved��b�������ٗ;�L��+)�1dӟ@�y���>ˌz�+|�R������d���l�cD��x0|��SܨΠ�$�P����ߝ�`�e�_�-zf����|��c*k��4у��=qRLp�<�K�����W'�PJ�����	mqɞ�&�EV�>􎭕��t�ƞJ�%k���U�/� 4V�����I���y�G�`
�](M@V�Eq;�c�9�<9��8O.$]|
�ڣi�c�!1���_>�NX���:����aq�f��"{�?���z�Y�ǀ�Ib�0

�@5�]�)�m�RH'��m��r��#lS�-y�6b��C���|K�2k?�N�F�χ�����%S�*�rw��[B�4���^��4��}55=�a�%�
�}�8c0[.Q�������ҝ�mU͑��3.>q�N��&�1X%���|c/�jڗG��L$��"6 ��+��(�o����n���W����-��ʘ*G'c��Y�ܧ,��Om��bW�E���g�w�A(����c��2�)���"�K:۬�va��5�w� �����|�},c	}3�56,%~�.������-J�x��_�,�؆Fe�^��N)��v�u���ߚ�z�+ @~<߈[���ұ(��)}!5�d�l��^(c}�=xJ8�Bд�(h��gVD���7O�?�>���h�b��ۤw(Q��6���TGp�$fP��/�	VD���a�S��7��:�<�ɁAnbA-E[s��e\�O��/׾�x���B2)^��L��x�H­��*�,T<�y�U�U�a ��Mu�*$���$ps������ä�f��y�
����X�ꣂ��2�T^������a�~3B�R��LD��[��)�5c[������OYfx�㑂l[,�ϣ���l��U�F�f��7���-2�����G�����~k;�uf�U��!��������}ǌ�rNH����@񢥙0H��ڮՠ�)Ǜ����^�r�[�)��6N	��[���-���uᕁ��kKd�&��>��_0��e���/C�d[\��1d�B%�e'���1΋��+(A��sեq|a�.n�C	r�B\ޑ,m�)�4�����mn]��p�^�-�)�/�.�c���#'R���s�|R>R���ӣ�|T�@ۜ����:o�o�Ol��F��H����>�˶%iT�C��M.�Ҏ���C�����DtO�U��s�{8${v����k�Ɛ���f�l�����Q���U�)��u~U�<�0�6�K �(�h��[�3#ap��qRPf �����x���]-^��34��;�i�K1���ެ�SNR>�|�}A��&	�
\a?)��$Ԉ�|���SǍ�
��GЕ�
n�8|�Z%4��ru/׷{��}^���h����.���m��`��ξ(�.���R���P�&�{��j�]W^씍||���赍�ܞ�#/�[6�먱��=݈�M��|?)��|u��S`ۄp"�\�����5�"[�y����ʊ&������ٸGY�Ԙ��[H\��U�z�*.)�A�ig�4]LE��uM�Ű�i1#���D�i`pgJ��}=H�7�%CE�� ��d�i�R��CkaW�H���]GWznJ���+�����)�W4�6-,��=����lG%��2���^#����+��*D�k�F�8)��;��J#�]��*:�ȃ�5��σNM���.;z��rփ^D�e5ğ�͏�Gr�i(��St��W⯚+�x���3�Sw2� ��c�8(���k`��}7Kc{�g�V�"�Mo��ၿ�Q�\6�,��Xb�+a��m����Z�i8�wd��Z���t��[�'�܀'�����<)��YC�X p�����v(}�W��G��y����א�[�����O�)&2o-�Z���$���H�4�}���9_�˽֭��͒%��Z]UL������8�2�ǻ�'��ۅ�O�uT�[�4$*!�I��5��q2��w6|���;&0~��r�v.-�.pR�G�(d�FG[^����JG �w�ɓR@nk�e��X0�kޖܾq/�k'0�]�����r��8�YP��i<=r�������4Ũ䌣r�W�<bΡE��;jS��U�b��ԉZ<��Z��7\�Ւ����(񱳯B�p�{�X�{o�d�W�]�ߪ�9@p��_�
 ��9����m�VLj��a7,��'3�W�.7�D$�PuQfE_��0���UG�ϸ��6�������M}kHt	p�-X�J�T�UV�6�ٍqUj��f�92��%��O]<�ڏe�!SVK'4�r87�=���{��5-�O��Ǝ �0V8��v�LRN�:5������<7��^�_�M�噚���wyO���3'L�}���]Hӳ�(��)�����F���|\9ĎnK�#m��t��+��/9o�;f��)��#��fL"��pBr o��@8�M�M��--���_�T��8e�_�YP>�&O����0�n��!)��F+<#�H;����4�`A�R`&Bo�5@O,�q�Tq�3��8
>�x-�!p�8E,��Ag�i9���xsG�2���� "��6N�`���;��q1s�i�+\���(O�u�����q!o���aj�j�k޴رRF�P�a�U�PJ�:�f�k���K�MfѮ҄������SvF�{�� �$�	�큸xZnxy��F�2� �#�	9wM*��[��B}'�BD���-y��C���9� _t�V��^N�����AS���#rգ�(1S�۟]�j!ǃ���נ��l�S���6���TT~+�É<2�=����8O+[�����FP���`��E�8"-wzr&4�����lLf�#l���0hDd�f����
�s;������A�^��BV��t�|�L���#��*�2�����+�5UA��(���� ,U��9�Y�Bҁ��q�������p3�I�;P��f����3�/@���|�f@"���[ǐ�3�|�8��g���� eWU�/(d���K��:�5�0��u�	�'�:�b3هp��4O�����?r!��=�N$�Oi�5�}��xʮKL��z�x"��g����%�Ax���,���s���!�!jں�Ǔ^����7=����P)h����H(����|wr���|�"MI��W��C�('D��P�j���x��Y'F�A�{#�Ϗ�Au`��r�����n��ɮ~�$������x�?�;�x�H�/=xŷ߰]_<JF2�x�L�D=�z'�o��L��)���
4���KTJu�A�h���$�5�4�$������/��cઙ+��,�XTb��_���S��8�o@YsO������,��m���Av�}�#g fW�kWj��` 3�/﷡���a�}���[zG"^�>�ن%�4�����3C����hI"Aȝ�Æ����2�gd��m�T0G���9�������{9�f�x/�X���^�ªR��R6do�{K�Z�Mjz�y�<��z��0�G��6U�)H'�����ޤt?�W(C\��A}���~k��l��]� 4e�^(�#iPx����L=�:�E��"!���A'���C�����M���d�G4pK�53{��J�.3���Te>��k���w���ΎT�V�a��/�7���S�rM��+Τ�u��޺&Nybz�h����&5���,�09;��~t�JF̒�H����pEer5����v��X6|ɬ���]���9���G���xST>��fk�T�I!����}=.�X�89uA�;1�I����������M�&�2��(~��5-1���l٢����'���(���u>ȇ�a��BP%�naGk��[�컖ԍяM;)�o��8)|̐˗���#�\�n�ʠ[7%�$s���g�%<lZ��'!���69����$����`�8X����k,�oHDX�l
��#��_�a���12��'& ww�Cs�����R��Q��������{]��Ⱥ<�	��?��~A��YΌ;P'2��w��*R��/Sd�P��U���)�!����Y���Շ Ԁ��	=�h����w��M	���������y��l�q��C	�P�� ��ᠧ���Cǫe�24"c���֖��^+NB��)l��o�&wi�)�an�-��9�i���� �y,��������o���:�Y!�%�>�֗�*�sD��_��q�E��O����5E�83�gp'A�Ml�W�Ϝ(�
�@��
�v��Å] yb#xT��ր����ml�=�/d�M�Z[��|J=6@j���P�%�ڷ�0��)x&_�@�=����P+�*7�07c���~pu�L��d8��i�1k�c4M��z[��������Jy�F�1� �
W�ʘ�ћE1"����nU�;���e�^�H����d�^V{0�Z]P��],�E�$�d
�(m �I�
�40U�ٱ��!�3[�F밿�S��)����VMQ�+Q-�9p*�N;/��E��V��eW��&;��l @��=}䰿���CC�cF��'�X���>	e|l�=��8 ,�忟�*�J�{�g�C�
�{��ZT(�	�{|���=J?&�֬]��A���{�.t�y<k���t/�Xn� ��=�qxxö��Q����ju���i8��qk�4�չp����JY�E���\R��z�KlK����")�p҅�����я�{o~B�����G%���glT�����g�
3�堇GEc�ro��㯹_Ӕ^}&��v�CxD�Yf1�7�yE��Dɋө2��M�ZW�R����o3On��3�_�EF��=��ވ]v�ՌDۆN�gG���Ji�*{��Oq��U��c�I]N���G�j���pcEE4���&�@�y����J��D������V !1>�\���Y��:=���3|E$ɘ��0
~�Yҟ�1+r���A��G`�ԋG���%):�3���ʼs�������-�a?'���a&�0��R�80���OmR����ޞi�`X�Yg[U��f��B �	dh�L���T����+}㣣@�w�x��=��\}�hY���{���XtBTR%K�"F5�ƃ�%Z�Ba����)�����U0���	b����D��%f�%r��TO�k�κpá�=GhC��B�s�4��T�5E�����lǆ/)dfً�|�K~����pg�`_R�}�!�!��!�b��NC���{{�d��m�(�`��hZ&���+j �o�F���<�������!M���ދ�MA���Rz(��1��mH,�?�%]�u�/4�~A����t2���)'JH�2�[F���M�gz�`e_^Atk� Z��GQ�hH��'�,�L�T���<^���P�y�x��8ۭ�8/�z��ظ����1N�p�qCw�y؍�4+15k��u�4���<=����?j�T+�,T�#�Gwm����v��Y߯ل��-�a���`���������˚�@����.Ba�Ǯ$�j�n�'P��pS� ��ft�В3�9_8��?V�T���"�hw���U���tv��k�����lױ��b�k��֓�=�m�s$P�VJ�	��� ��8���9�?��cUAto�i>RN�ע3O ��F���B�%�|��Z�����Ta�vD�l�`�H*%�+��09����1Z_�g�~hy-q @�J�c�{�E������7��Ơ����,�����$_���3-w�!,��K~�6$���O���G�C�*��ᓹ����9��Fu�``jy����2�\���Qɒ�@T�I��P.ޥ����,Kbn~�N2�`q*I�b�@PؾC�ɪT���X�Or�u��D�/���k� 
	x����]���eAbAl�����|����y����@?��B�z�~���Ѻn ؅)�$[)[�Z��t�yh�R_�s"��a�I�m���Q*��t���NY��g��p�x��in����2d�������� Xc�����H_�h��P�K���-c���}�f��ⵠ���ZId�6�Ζ��)m�rl����3'��B���"��Pc�8b�"�:�ZC�mo��L��0���Ǎ�Y%3E!�~]���T�2�2������͋�?��rh9Fsv�w"���с�!�k'��dVF
����^��ˑX}�G���r>�d��P���$s�E���x܋��8�Rc�V ��r,�k�W���.�,�;�����6�U�����_,>f���e�S�bx"�v����Tz�Հ�ɔ�&��aww����<~�Z����Mk�'7�=�zhܧח�ڹ�������k� !(/��H6@.	�r��Ȧc�%[q��?�n�Ј�@���6?]�Z��q�>�ц�?�\��RՁ�w�a�	=Z�0x�#��]B3?���U4X��-�k��-[�\��`�\j*b�����@Ďo�򋛓��)����]eP����o���\{���\����L/W4gT��_p�$Ή�[�������ǿ�˺vGP�X"S���:��j�h3Y-۷A4���^�hp�ɇ��^᩷�(�"�����;�]�h;� �́i?Q�wY�R��t��b�?A8���	U��f�]p��0S0�;��){ԍ��)��ha�@��2ɿN�S��B�>(d�yv�����/0ѳ�) ��4�������M���Sϫ�xl{�x��;�0,� �;��$CD��*N���<-�+g�h�+��*A�ਡ$��e�o䟚-�	54�C�F�������!y�~x��B���_�4�啃���|k�g:��O$�g���K������2j�1 ��:I�2�.#<E��B���ȱ�Ǉ"��=j�	�c\��O��O���צ�6��;'��j;r:�e���cOmWs�x㓆�|b܁�Vݙ碷��֋;\r^�t5�aM�_���ec�w����5�i}62��C�/��e�쪵�T�?�����2��ϯ��ӑliJ��n�E����fj�\�f%݊ �w���&�����˥����/Z�ח��~�ٖЎEJfCi�?�����2���U����hEp��TC㷚Lh���HC�>p-��1t�=���lG����AƉ�~�֟P�V�� C{p��B35t�WX���(�l��3�����CяW�<t��x_�Tur�ίU������*I���_�㭭*�"�R��l:^�����&z�o7\�*�D�5����6����#7��L�8�nLo����3X���q���驫�w�EL���zV�l�3Qg `̰�2I}PYōM�z`��'I
9j1g��5�a2�0�Y^�P�̇C@��Z��i	mv��r����<Q������d���}��/�����.'�+��ߺ6�������K�+R��y�@����gr+zѓζu����SF�g��_��X��^�A�w9�Q�z�%�`&�(��M�~���;e1ϙ�Z1WeBĶw�҂g�ά�n־��E5�L:�[fb����M�i.@�ހ@lg��,�Q����Cpz-�����o�w�<I�Έ/ �R)���+V8��A]J,N�r�d�,.j����A�/�
�_�$ۚ����#CKǡ�y�XF_��>��v�睸P������2��7˳�Y�l�L��ޤ\�Vk;����7���D�T��	���w	�ˡ�Oļ��Z1_~%��5{P��!�R]|�A�c�i9��]�>of��jI�0^ҕ'q�}����D8�iu�4�$���A͍�wD�,-%m.���JB�<K����T�r��	��g��:C���M �n��g����!�'3���M�T7q����"V3��k7�T_�������}	/5d^D�1��y~=�����&�����U �"�f��x��������_Yk;89�F ^cG�(6�VE�ɨ�[�`���q�����(lb�v]܌�m�]�]a,��N�[�����ʡ��.h@ ���ceWg	z�æ)�ʳ.	�;HkYW8�D3E�L����-n֡'�*.Sb}�8�,�0���:��<oG�G8�C�FdRvvḆB1�-����r/]p��(`��p�6������q�Cx��m>k���C�bf�{^��E�R��`Qr�>;w��`�^��7���o~�!�=���̂��p�֨g�b�{S��=,3O��D� _��**����P�sM��v!�Yɛ3�v}�)����8{��p?�� ����� �6C�b]��pJW��U#��_��0Ch�\R2���#4����:w�q�)9<��~%|nv"Y[���4q(�����@�2W�c ��Q�ݹ���6s5�>'u�F�+��;���� 6"��6�6����)��N�z�7�.�n�2�q�A�|/8,�|:ēi��xZ/�\�an�ľ ��'���?9��0X�k��SآD>��A.�h��X�����9{c6�6�l���:ƘQ�l�/�r�ז+�m��$Vc\�ᔭ��E��k�P|&�]� D� {(T�]�:�IbCs�z�+�����0�}s)c��_�	��~�����Xw��vri&�o�[+� �g�����ZX��+����]�ݠ�������6A�l�ui]��l�^T�F\n����.3������ 4���H�R����늝���ׅG�/,R�,�Dw����< �i2D��|��$�~���Cά�X<��a1A�u�3ߌ��7���F�&'�����+�\;��{E��o�hfK���H`Pw�@�6U�#'�0��y'�����h%�y{�q�胱�W�&s��ft�}�(����}�뒵��r��`$.W&����UC����5G��2�_�7�=���!�b��>E~���_l�n3
���4����|ϥ�,����v�ɅZj�V��O�[�f<���	�?a%A34h��	�@���N�u�T5�5�A����_[�:��m)���u=ޓ�`:n�%,z��2q�Ҩ�KSC��C�=��5�~%�ğ��Ѳs�]y����檬W�qT��5���c�$2H?�p�p�k��óB���G[G"TV$D%��]��=��i��
k���9P�ً�X#<���
��d�!|Tl|�@�������wy�J�0��pF��@�$��<shR�{�K4��!�����<�j�>���o��2E��+}e��&w6��vuNX�����vm�A��as&	������i��|Ԥ��U@6o#���v���m~�%XX�b9�]J���l���BHH(u�gd�$u�mR�Y\���`���	ϼT����T�V�Q�R&���F�IA�B�xz�Rcq�����Ż_�V�ޔ��|h���ޡ`�X==�j���eTBC����A�n�]U�t[<%gN�H�����j3�0O
Ü/���ߪ��P��F��B�e-UA�z�V�X�1�Z�%��]�FR@��]5��dn3o�1akU�c~�:#bj_�ݞw�P{�]U�
�����ͣ%/z�Kн�z�!��ٖ�870�k<�(7-�`0���r]�F��șG�\�c�k�1�1�^jt)k��u�,�.�R���M�)PI��:T�zbJA0�-/
\R�}��@<�#-��ce[P�G쏟F879!n������g8�Q](h$OTYZ������Z�i��F#Ào}��7`SF�z��O������W���� D�҅C�3��o�Ʌ�(�R��k�3*c���|&�*�J�x8��yTX@MƐ��;����i!i�����w�!�s)��m$�&Q��D�*�.Id�%ϓ)	�'�>�,j�k;8d��H��l�^���_VE+�s`�C+������<�Vr�9{���'�����|�[�ڋ��s�w�9s�2t��<K�!�.��R.&�P�>'�V��!��w��6������`�d;fs�$`�0�� �$��a��?�#�қ�R�O�u�����%nM��ʀ,Y/�.=�@�爆�x]�.�K (�8Ŋ�/��f�!(�C�~�J�w�J��9D�;U�1��ٞ�`qW��,(1�������O���>&{����� �o�#�(��?�u�I9��3����|�%�o�dܞ"YJw[��lPW|�2���'����g�l��\�a!�H1W�n˞ˌ<�oc�#Y�K�ĉ�!"4C�J�U�\yO�N]7���v�9���R�;�Ek�M;{�?��o�u!�G��qO�O�S��I,�m��qmt\2#����T�&]p]��
��r�#�ãu��n�g:懮o�	�{�6Ԫ�<��!��Hva")e>���D��8��#��b��#I��xe�k�ª~hȒD
#��1�%�dN��Y�6,�mP�`�'�;��w��k"�) \�.���ɶ��#\i�H2�C��(�\0)e�����W�^�6�![���aT�8�A<dk̈́ɫ{����Q����T�]������{"1?U>���&h ���-�0><����O�� ?��X�l;uQ��%��
i��m|H_���{<&���s:�ߝ�򱂨��w�AY"iR�6\�pF�xE�J�����~���_먹�A4:?{��g�є�[{�F������7�:���'�3p>��-&T����]]��ὀ��1ʆ,"�N�	��]����Vmk �e���F�ԻH�v���t�Ǣi8��"�w���57�[��6����7�����	?��e@^I�����x��Fvd�L9��J���%y���t�!���̣oG�)�Ɛ���,dhAr��)��ԅ�]�*�h�����nwS��:E��l��M o���B��{�v~!"9��[��M�TCr��poI���"*
6(�5\�M���K�Z�xQ��c
�<dP�����R{��V���
��i�}A�3�_��o�+��)��f��.�Ũ�6q��/9L����ҟ�۳�4T���'��ѱ/��s_d���[�R��
�O�1�6����WVR٥�u^�~�'v_Ik���oi��ٹ:��������#���PΖ�1��Q���y�о
�+-�$������z�{M�%,=�e4�50��wƫ?�o��\�% M�c��w�%�5א���c��}c��vġQK�OHO�ͧ��+��g��Q!/�5�nz���� 	���{W���|h$�#�`Ex�܆�!�ZՋ���x� u[�����Ϥp@w�u�-nE�%X��d1`a���	�}h�F�U�f<�4��1ߥX~k�p�P%sq@�3HnJW��t[]c��po`)S�t,	�8�N�����^�!��8��L�*6�	�b��c/E��oSl" '`���Wd1�pR����u����t��62�/�ScJ�B�=�u�i?����v�XhbNp�a��
&9���+�@�	�D]����g*C��$8�!F<�t��{9�&ߢ��,F��U?����9�R8��1�H^��%::�Aq����m�Q!v(M9AiX�Ρ�V<�[*��>�=�r� ^��&[x�=��ur6!�I�9��tZİLb4<b�^cO�[o���Z������ȿ�-1x,b�<� ^>�ޭ����3[
�q��h�x�ˏ��_{#��8eQ�'���-�$�Ԉ���ٽ��  ���'�0��y7<��/�6�I_!�J�R�A)�⼺^m ~cЧ��$�ڂ��g'�B�3�e��N���·�րL7%�,� ���"H+.���U�ղmm^�-	=C�)��+��'65\�0��N��9�Ɵ�0���:�lSl���6EQ;��_ �q�2�Vy���_���=ٱœ+�ڂze�bYfxs���S��L^F�w�Nf��Ε�I�F���p�$Z����8m�iH~�>W�8��?�ǻ�89�_z�%!�L7�{�$Yj�c0��a_PQ'>ˮrS�!��.�;e �:�����p=�i28)�я��J��K���8g@��(s�BCw2���"J_�]hj'wlk�/��d�T�X̩�=RLL�qz��X�b��"��4���qV�D �T��!2�Y�\3�2�2��i����bƟ.�{f���oU��"n���<?�E�&7��Ά�Xxe��)����ȷ�WJ2�P���4��͐��\)�~�v�c�a� "�[�+��o�!��'a6��@�_�8Tv��u�v�C"��H��./T�}��+����}��e�"C>�sѥ��ݾ��L�f+�f��h�G4$5���~�A#��s�٥���.6{���2�!`�7��n~����Ï�5��P a[5 DY?��g���hiõ���΀W�~�� ��б(���e��n���݉�j��
=�5�>J�s���̜��{����nB.��d~��o��ʙ�*RU�X��r��Pv�{ �B�����.Ϯx���T�
�z6��C��$�V$240]Z�����RMۅ������X%Q}vM��5�G	�@:�í��N.�;
�k7��4�6i'�zl�էE�x>�dd\�Lkt_��G�QR�+:�/��'J��f�� W8o �ty�Gw�DJ��B�hP<���T�"��Q�����ng6|��G� `�,E�K3���eF^���`ĥr��=�N������9W�+t}���Y�f(����� �Ř�N#D�gO�0cꭳ�9�'ݑw6���s��#�[�+Cҳ��T��P-���za�R��Q^�F��o��oݓ�ć
��3.��Q°�&�/Ant)����7
,X��'T��߲>�y6������jR`�4���.v����t��-�Y'��z�P4���T&G{��=�$�p�qo�n.s�Ch�g�~6¸��'(\ݢB���B�LI�M�1!i��p�r��+���E]��6�)�7�����]^��s@lR�@�Ѫ��P�9��}/��>�_lDX^�=���C��2mm�k�
��K���!KZ��=DgE�t�!B(��!1a.���h2-������LF��Ғb���	��f���Ǻ����!Ͷ�'�yqs�Yr�)E"Z p���ZK1�2����T�{7���YH�zw���NDJ�t�h� <�X�L��42�K/��Z���S0KJk@�{���fC��7���v�Ss��9h"�ϖkr%���F�pQq𥶏�~n�'f<�9\n�a`t����`_E�[�1��Ar�1#6y��i����j�84Q���i���X�P6��ɩ�d+Ƥ0|�K��rK�s�6����?I.7a��E$�5w>�Ux�؅�K�f6O��\n��Sv�����A2̑�.R�YwkCύS8GAp���aJ�l�r��d�u�Gq��JW�J,�?m��	����s ��FTP7�� M�=�]��&�����&�y�A���9Q�^�˰�����z���|d�;��l).j���I��M��+�&&��.�/����{)@�b���8�u[��b�Sn��s�K>�?w/`zV�o�3ar6"ڣ���:���a�S�-'_1N��)�D�D�%��L~6"ž#�āg��5�Vl�}s2��w���Gh	���@�,s��ϣ&.���Wu<o�k������a΁���_^��>����4=w�g|��܆?}��'0VJ� Cm�/��&,�*;;gw�D)ѭ�(�*�۷�x��tݽO:��]td¼
�r9�G�I����k�f�s��C͋���+�;�:��&B� O�P�a)g�sǤȁL$9���]O�>vT�<M���|�Di	sೃ��#�9�McB�Y�g���R���������/�؍�"����+�`{��L�W׏��Nt�'c���6��3Gw׊�,�~�����ogu\6~U��[�N>y��}�t�n3�Qp�	�t-���ނ��`^�"�]�"�L)�3䂛�b[�C�����}r�F" ��2XM~G1'���`)G��_�<[��?FN1$��
��� /���F�OVW��p���Z./�{�%����PD�B�!�������A5E��I�C��`bEt$�UD2��yE*���<I�b=����R�fǷU�d�c��#C°�X�`&69e�n?��s�E�/�R
�	�sk\��?S�h�,���<��@�Z���y��$��/Pnyn�.��Z�aM|v��ц?{�G�!IK�a[�^�l$�K����X8�Ӡz�����e
����pc�j��K�V�X���g�7�C��V}�3i���i�k��S>� ��뉰�#�������x<k׉��:���)	0�������Ӈ�:�b�3�V˨̵	7�__�K.��l�F)ʋ�m��$<�ã�jZ	�إّ�D�'��pK��T�O���:�����#�ñ*j�9	������_ ���E�<\HV}��r˦/��V.y���@HF��ō�,wٴF7R�s���|s�k��X�i"�M���gv��6�-IԼ:�dJ�U��dJ5UGC�s�Qڊ��ũ�	�1Yz�FiOk2y�~��A��ׂ�K#���9\u�S'��Cܕw�pgG\�r�!�����pw��Y�R0�Q��k0����ֱ+�
t���"/�O���{!�zHo��P��m+�j�y�|=�`��k�m"�g��c���iB���(�+U���̖���� L�G"�^��yn�ᾝ.��T����׀��\�l
�v��ۡ	�dl��"�R�x5�zj�%�|Q.p��$6�}����d҃����T�;�(�T�a�.W&��hT=P+b����,����䮴����\Zֻ��ʝ���t!m.���ɋ{�$�w	�nB�=��@�\`�d���ҏ�S�
 �C�5��ჽw��E7_  ����!�\F��X�̵��-_��=�H�\ki�_�c��^Z��]�6���w-�)����$m�i�&��򴚇�et	�V4�o�Q.���Od �/~g�^7����t�A���H�Wq����4)B����L� �s|]�?��|��*���� ��e?N�	�dcO:Ϭ[CEy��ٿ�;�����b�v|��:�]wn�۴m~#�z�q$@|�'���75�)x��k���\͛�I��q����Z�En���.�ģ�zܞ�]o��>�m���U�p�^j<���EV\n����Z13���M�lK5����ʻ��Iq�Q�A���r����!��{5��>�\�.9=ގ�����$K.RŊ�̡ڝ�b�������cs��Ԡ`z	%N�t�E(�� ��ň'�8Z��0��E�:�a����^g�T<�9���'��8*��օ;#�K~m� ju����ى`�j�JL�T�S��L���	����(�0nA@����3=����j|����M#黦^v��tf����p$9ڬ�ڥ���� �nN8�f~���x>�C��~�ي��o,r�J�<�dR���O���J!A���]9�d���
C�9��?�-D_�t�(��/��HØN|[�v�7c+#��B�ЭJԿ%�b��(������}p�cN�5�7_N������R���0T�u��@��$�6,�-=i����f¡~݃�1C��m�U�n�����91��&�N��T�9;�(���wQ��sm�6ͳ>{t(�6Z�l{��<<�s�ށC�;�s���/�D{��=�<��v3��TG~>W$Eh󫺱��ԍ ����<���'���RD��E}�X�l���a%�X�@�k�y��\�'��B�����Έ�0:�k�����k�����D�YT�p�s�|���0>ڶ���fͮ��U���*w6�)�����L4L�\xIQc��,$���Z���5�g)EH;������+Q�u�V�ݕ���)b�����d�8���(��:v���[tX���kR{�#��903S���x�7���v�G������!(9Yd�	/Y��ї#���ӫ����v���aE.aj�Ӹ�A����	�4�M��VA2��&V�`=u+el�;N"�G�1�zx%��G�`��g ʕ���{�!����Hdd��qї2��7���%��Ok@��A��l�s���)����s�h��ˇm��Ϧ���}�s�pB�-,ŵZ[�4�^D��8sG�#�.��`�a� E�@�%}c�O�54QB4�1�w`�wb��=��^~;f��i��_�� M	@���o@���W��7�w�j�ܯ�]xu7�L�Z٘�G�F)D��Qd�x��MQ�!�j��Y4)M�7<��?�������࢘��xك�쟳8�"�B��$%��޽�(�E^ٯ�VCD(6 �t�qg����]|E	+"�:6�,Dg-�ٴ��(��0ʫ��w�`�<��d�qA[��5K�eb������
�JfB��0pO�4������;�H�wT��>����r3g�.2�0�P�3�u��Z�)�L�4mmz�-�S��l{V�㼮>M��	a��Y��u��u�+�ۿޚĮIxӅuv�+73Zn=k�*�f�#d���/��ع��KxK!�ɱM�K�+3Te�:����P����~�^���7ő��ۤxك!=_�˿��k]��̧�����1�1ʤ�}��jۋ5��L���=Վ>2R�6V.5���:{qa��K�x6�a��������*LX!?��e�L]X����`��o�^-��ŗG��\R�fA���L�]7�G>�R1�ɜ���H����DL��#�y�䒬1��F7���CPs�� ��BYu�|��
D/����f��b���ĵ%0a�D�	яaf
xuo)���������K�ub�s!������Z��H��Q�ٯ5����vƆ��Of�JE��DB���?,��^�Rζ�����X�!O��j�1���ȝk� �sW��60�d��YZ��x1;�Y�7�z3C�#^C��"�����1>��>P�еT��F5={B��Q��Jɥ���ٝ60���Y��!�Uըr��xn�9M�G��DK� �F@��sU��RMBSD��֐������gD�T� vd�;Ԡw>^�sRTB����ڳ4�q��_�l���e�u�'�#���.�Р|Lk�.�X�q'LvfD���G�~Ց�8�C����J�+K7aU��@3���뫫��g.Tk&��ޗ�Q�Wh(���ß��m3����it��i�ؤ[�� �&��&�3S���4�M�N�>!83z�ַ�CODAJ�����H4�d�7ӟ{�]d��4S�C�oP��}��H�{dO��;���,R@<$��1륤'��JEC�錸D��B�*�N��/�61��ID�bW�쥤R�q�ϸ!�q~�𢦍(j���m�/���/�R��$���Cx)#��m�S��q(H?q$���������3�� ��?�1R�a7��P���Y��\y@��z5폼V�	�$M�ܜ]�Ϋ��� �u��MR�n���G���+����0­��/*̗��-)Z7��|�	&�����2GǘL��&R0l�H�\�K�䮲g��S��hI�j���l�|��S����[���¦�Xl���+�Ё�#�O��)�"b2���
���ƯBᰄ<'��֐Y��P��&��-ܬ�UZ�����J���*�!AMA�Վm
�C?ǽR��P���uQ��i�(0��暺�~�Y���� �y/k,��Vx�:�����i����a�(pxd�p�(z�I�Y��0��
v�^E�,�)&y[�lƻ�f���ȫb6�*ڥ�1δ�/oB�mK���,�j����Xj�9��4��u�ܜ��m�Y����&�Sh[l�X��oIA���a��+�#�J�j��&Mdt���g?M����"zVbB{�z������SU��O"�X@� �%����E�q���(��ix�u��X쏡3B�a�Ͽ�����q��ٸ���f����NH)0s*(��p�p&^����v��3���ޥݎhG��M�W��63Q�,e��j�b�0��|�:\��%�M�`�J:���V���T��±S��jrY��	��9����ׯ����H�.oxs��Š~20�4?���Z+; (��[.V�O�a�8C
�BU��E�+��Q���S�!?�"2�)i� ���<5,����%��F�.�zg'6��i�h�Dq���Lm
V/9�(v���/���.�����]��s��<�R=�A��C�¤!��f�҃UB@����J�(h;���
F�i�|�}�'_q`��_��<xH�L�&_��*Eq��o5��"�V�_�A���5~φ�OJ�P����T��G�C��2~+>�HDzHw�����~�����ՙ�*[}A#�^�.�D=TP�𴬑v��TP:��;ܜ�ia�����3�Qƚ^g 1��f]��(��*�:��ӆv�`s�w��۳2 V���3-��4�6A~��F���~��N�*�-	H�Qb�eT�q����dl{FM@��.��6��1�_��p�	���^�F�m��UM�G(	��r���Mt��GA��]c��I�-��#PQ9�t�F �e+$NS�ثZձ������|+z������~X
�"��#�vdX{���q�M7f���C� -��Ӧ�X��,B�o�0��
4 Z&(�.0���f�g5=K�+��.=`'�U�<K��B�ݠ�>w����ps�� �����{S��*m�m�m%CM�Ud�q����^@Ε̒,V���yj�ˢ���А����oL8oN7���L�Q�.���l��Oj��II�.��Ҷ�ɍ<r�J�B��^BB(��4�A���$�.gޢ�>�m��y�b�8�����p�8��K�_w��b�A��ٔ������C���*�v_;5���єg� ��K$��%#�:�;�x����u~��!���ε�=�3&���Q��-l��qN���Zm2�z&��~�8�4���:p�\u���T�?�i:S=��\.IxL��"�@�`[U�銩E���l����m�� R`��{���EIޞA�I��e#�K�x��8��$C��RJ�kq�|1�f���ϥ���\�ݵ��O���}�D��.X�{`c��Q�,pIv����n�vxx�4%B{�%�l[%h��;���߉#*{�~H�cɐH�K�ں �E'�~GF��f�{8~����£N&$������-x*	����b\����K���џ�8�_\���Of'�ME��mZA��g��&��ɇܚ�z*7�I�G&����l/-�A����.�"ﮂ��d��������]�^߰Շ�++d�y[{��P0��P����*��T�5�Qo,�ߥ�I�w,�<��!�ꞔ{H?5���U���+'X���3e1��v�!�Ʒ�x]���{�U?@Z᪞RoQG*��L� ���Ȯ�pk��)�c�]�Z��O�2b�Ӄ�A�XP�������>�J�������18fkc�D]��ͮ��	H�|,WZȂ�A5$j��$J��\�OqbSh��ѩ�\�D1�R���pc_
�t|��<
��sV������㜯��B�<���J�m$�J/�[��i1�ph7<����f�kCrʦ���f�������i�*�luۤ~�j�
�@j>��PW,�oO��a�8w��6�-� �����;��vM?�4�l���$�b.���xa[�.�ck˰�=)9���μn�`T��7����	�;&�r?B68��Pku�T����nhςG$���`n�,?��\t����HL���Ke�IҘ��z���5���p��Jv+5p��#�Vܡ� �X��'��]�6ԷrM��.��*OE��0lm�s��v҈R�����u1n��nX�.��쓍=�����oǋ�?�r��?�:��5��U���1����>[ј���MG�6�j$Q�M�Ee�f�����(�1��W����6�iM�L��ߣ���b'9�S_-J�^=���� ����;8�z���})IBz�aA*�f?$R�)7�4�f�O��9a��+�O�k�~i/9��#~%���(�̰�Zȓ�r�)�R�4nS�@�I�qdv�]Z��=_l��_VX��ѣwG^�p��@��u��1�8����~j3�\������7� P��M�J�^�"��fy�}�#�)c�|�Cny�=�m�S��j%��ܡk 3���֓�@��5_-�F-^��9|w1��PȒu������,��Ǘ��WL����PY���_]}ן�#��8�MM�k��q/>�*�P%�r����1�ǂ��������Z�ᕑ�"'�˵�D�����{e���G��{�RC�%���D)�%�����Z�͙�7jj��BS5����"�M�Λ�i����lP�z�4�ޛw��\}���-��[h��@�h�KOz�P��\sџ6�C���H�K�oX2K)r}| /Bח�6�]�ƌ�(`<���>0���T�-�.C&�Mi'؍��,bS��G�����K 6C��c������1�{���a�$Ÿ7*�m:-$M>:w�8w%�C�C��a:xÚ6r?,�"�,H�1 ���ڟ��%�#�t�w�K��9�G����3��~|��;ר6�]6�G\�����c�2AH���ʒ�S���6�4�|������-	u�˭���H3$�v0-�0�f�U�@k�<��؛� ��I��U ��XBPE���Lը;�sޚ�.���B�C��ωҀ��c#!�փ6��#w�Yy�ڥ3����o�J�"s�8��q�{�.7�o �x���B���T��4�/ݻ�:(�������ء���g	�_�]Is4I�{OZ �����̅�Ez�/1�-�Pz9��m_����=�ȧl�go���Dc�����(��q+�����a\w�;!|��;��86�;�N\�I����bɊ���.O�Ռ�^�zi�w��9J��fT[�����&D�is=��������;7���d¾G;0���!��x}���� #�p��{@Y�cc��p��/�xL�ƍ4u�fM��M��ӭ5y*���RF�|��z���PM�ԗ]S�����8�H�}�|�5hQ�Um�<2S!p�'J_��G~�K�d�o��
�"��P+־�X,���X�]ڷ����Czm�A�}Z�<�����r�Xb���.ϑ�tU�z��uy:���UٱzI[�go���J�ʊ��a����h4��}�d0`�A_@XK/�����q�I��! ��8e�ʶnz������lZu>�P �&l�~ŕ��C0��$��}�t#~[���4;����?z�����9�j�#�V�o(�Y���MLӬ�B��y���Z��Q������|�"����j�m*R*Q��.F��:RI7��s�E�TC��@����>�bض���k�����&����Ӵ.��3�]����`8y�&�(�=У`Aj�]+���>,4�C�]<zJO��<�uގ^��K����bu�{���� ����FЌ(h?��OR�F�j��Qē#���L�J�����j���nz�m�f�WDC�]��	�����Ai��}��Wjg�%S5J�&�A�S,�?�]��1�����Ъ˷I�o��MZ��]v��hZ��ޖVSRK��o�I���m9��߆���H	�}�H�r��GBYt+��`�4DR�F�������&��J@p�[&���a� t̵L���=��
}���C�1��<^e}��<��Q]�{�@�!�c�еx�0g�I����a��<b7�{T'����n�<R�k��L6,\�;I~p�V�\K�j�
�7�����yUh�߯&�H�;<�M�S�c]�ޚ;�%�i�y<F��Y�]�.�:^�3	����?�b�d`јH��B�c/?�Γ�Ҿ�T�R�qL�zZ�ъ����6��K�y��`S�ֳ1��\��.���B'F'<�O�$nvB��Zb� 1�h��
,!��'�͝�]��vGU�����y�#�Zn�vw�cIN��P0�x�M�
�^���6����q�c�'o^�P��a�#d���-�Z��$݊]�!�L��f8�:���}��X��%ޠ�p�=v�$e�G�k8}#%� q��_Ix�O����:yxh"��v�-�V9��'�&�Ǣ���HJa�H>����ѭ�� ô%dA5�d��6{��3u�d�V����*���s�C�v$�!9q:�Τ�, Bgf���ԧ��%��Oc@�,lt��~�K��C���v�a'��!#���l��&�/<�:��p$��eފM����+)�5��?-�#:I��+ ��"����
�]��´尘�7���e+t��y��^��=�����Kn�v~ĸ�� ��y�#ޠ�]������-�����e����ݜ6���Ξ�OXy�jZB)X��giLl�Xm��DD��9���l*��z1�\߂8R1Qy�?aVҥ�g��u��>e��l��?����@�'�v�U�*t��o�h��tF�������C}_]��;z���e�^Z�F�|�����ڑ�T:R|Zr�DOop=��?i��ׇ�V�}�U�֝`X�%2>bL]V���E��cK
K��h*rB�uL���{�d�v���[Cϒn��Fώ\�8��U�R�C�oR����<���~��<��9'քg��I�+7 �<&�E�Rcav�&>"���1�n0G�:Z�h�	��{py��dr��k�u�?���SeZ0|��Z��9��>g�5bϴ�zquY�Aѿ6j41��h2/xh�YVqr[a�[��f�_]�u~U݃
a^��XXYb�����h����ٰxkO0��Js�m	�B#���_���ڛ\f�4���E��ꮵ>8ɥr�@��x~&@��"��7�r�lZ���^ܴ4���@75rU�x8u�!�!&�($em>M5 �B��m�
͞��)���#�S�&�U�#l9�"����'DB�a9W�K���:���<άIr�v�+���@a.Eǃ����+��'Oxʐ�87�R�LК�Zۢ?�c=�vE"�i���=�6�8I��JbR�f�	]��˾v�u^��� 	OKP��p��3u�'(R�Ȫ����k۳W�J�ZG�I��J�]�e��_I��K �	1���(T��0LQQ֊P����Y)�����s��[�z#���ꐾ����$	X����4� Qws_@?ҔD�*"�G���I��v�w.t#�o�8�e#F�=h��.�*�P=E�fɆ��Z��\G!6(J���>l�ZC[J�  �>8��.Z���l�j�먡J�_fz���ֱa��a􋭢��x��IB�Z$[�G�O��>�g�2
�jN̹�C6�"�]��� ��}|�=�|h��L	��  >M���.���X#�jS��K���t�A�����O5j�}L8�Z��zuL��m"QI����Fxz4���������XS�����w�~��_��.��0�����TW~GI�1�C9	�NA4����®���j�f�Y�-�9�uD4+ ���]�-�A;�|���F9����V��+I�IlԱ��'��G|�0bڒ<��PL����]�-����s+%P��hwf�^*�MD�1�m三�0?[�ySB��d�|�B��Ӑf��P~�]�o��Ӆ��e��+8�ԏ���Uw�jJd��d�W���Y.+�/�g"Gߢ�:��Z�����^P9�O�H �����p�0�j��.}[�JK����<�T�=��C(^}���H&�Ahh���FD�� �C�������+��x[���d�\4@ |B	A�'��[~�LH�^���
<�ǃ-cϜ�d��4�L�H9Z���솶�C��e������#m�W�cgɶ c����V�*5βO'H��뷏`bT<" R����h�SGʗP���7�'�3n����k��`D�[�g��
�}[�~����Ԙ���PB��J��&2�"G�u���%���%�/���_�C���g.�E�P|��'�l
��e�J�0.�,O�����4tk�3��Ь&��[n��A��F�ַ6�杍�y�Ș��]��ocu��G.Kut�<�(%P4��i`Z�阮ϝm�*���I7ˁz��N/��3O�|�����f�Ȟ���BC�d`T��o_�B��D�hj��c ���Nh��Y�,��e|V�=%��t� G���{gB)�W�	�E���x�_Ʌ���j�|����*���w�H�7��ȈbZ��MKW<��K�R��nG�g%���Ʒl0H�&�Ϻli::������w��"�,��4A���i�2L_�
9��zX�z��4�\7:�6O��b��S���BǁTa�ZY����aR `5h�9��<�ۈ��+��#��[4�'��x�TbD�n�E��^w���Qw�ҙr���Ш�h#pap�V� W�^�q�=�k�����-���{�u|/�Fc�%O�D��V�ʻk�4�`I���g*M#� ��ld�>�w��c���J�i#x�L3�_R	e��p�x�>��ۼϔ��T⒰�~n��wp�8�����pk�2�:˄�hu]�n��aa)�I`` �S�˗�8~YFsA�[��s����~���vI�,Y7�&{����[()�)ޢJE�Q�;��ݸ=k�%����k����cf~�){&��	RM�#9���Wx�>.�]\�Nr��������1���j�@ ���Uف�t:_:IO�D�c�}�kL{L���$z [�y��^��ps�"���ɹ;X�xc��f�hv;Y?Cm����01r��Q2#����R/'�<��	ߺ�סN�+�#�NQ�ۿ�총AnF1 j[�_�c��U6�U�q��~���c$;˞�CK!&?�� [޽��H:�H&�0����9^V���h������W
�����s}���(�}�L�qf@-)��"j_3����-���f
_iY:�
�z��V��R�a��_�n�D�CH�78dVf�u�.I4������F��&�%���l�PM`Iޘg��|{�tF6��� ��.��xEV+d��h����{�vӀ �8�Q2�����:�HK�<�*�F�>�/���4Y�z���z�{��>�:��A�b*�c�"�-Ȯ�/���u�\O
2?��e�L��>��*e���;t4��c�`�0A=��b\��3���\߭�>�":A�+�?�ժ��a�2���_M3��5#4���+)hj݄�Mݜ%Ɋ��/AW?22�P�תq��3����4�_�5��R���2�=�y�����x�!���G�V��!�C�M�mK�SZ���Kn|��̿���A�N-���v��m�/޻� ���?��lS>��*D��Mf�L˖%�d4�6��
�$j�����7=��b�� ��(�;��&�YRwp��Yt&���#j����y��磼Ǜ:�^$�t|e�� ��
=�ĥv�b@���S�����i�AB����f���C�	�<���\�T�wD�	��j��&W��[����L	3 {{M˴�ḕ�K��"9,�5<Y��&�BP�i�Rd��_7���n�59fh�h��:vF���tݩ�G!P�]Ә�7�SR����>U�L������j��Xʌ�����;�Qs�H�m,�����t:\Qݸ�����ƗwwI�JN46��X�y������S7t
��Da>/hlo3K
�D
3UL��i��.�'5e��^5#���>�}�c�FA�pq��=�1�
�L��7�cA�Y�K e1jp/Hc�祔{B����WU��� �s.M�Q9U�[X�� ��X��ϩ�"AmPt#���4g+BBUB��K�qX�"k\l�[~>�$A�!��e��%�j�?�`��zM�������񀚛�iC�|�C�B�@p�j��u�UH�񔡬k�-�(BF����d$�=�{�.��/\:��<����;����B�zO4Hg�j=��o���\��JJK�u�#jM�����o�a?�:��I_�ٵ�ݭ˖j�X
u�[**�F�qDso�!AIC�`��em}c0���`2~4S�M�ʮς��O��������e;Y�o_��"�|�����H]M�t�NÏG��=��g��_\�L����0|W�?�ud&�$�r��#T��%�+�F�褜%��RJ{�?V���P�7_�&��vo�h�0b�Y���\P*�����lq�a�NJJM�_�ϑP	G-�e�q��T�*����h;\{V�&�{��������e@��3�� �˴���ݩR��	���2��u�һ�:'#n&��ĩ�^.�bS��u���`���xNes�������Sz������5,�M�o�G �q�7�`(��{�*U��v�������J�,���JuU"�3R)"/�.,T�����gǠ��9��$�ezu6�~Ŷ�sU<\�9���/��kA�f���]�Z�eh��a��Um�E�kw~��*�n��#6��{f r��Y=�D>�_�o>�m2�	��ؤ>��N�n�,�{�yw�F��	$���r��3��35�R��M%5C��Т��3-�NdgƼ�*iȤ���ˉ7���9��9����%�_hi��c	&��R�l�"���K�����b�:�#s9�7���
�+,�^���Q�>��q*����m��h���F}��n4q�[e=����i�h�=�d[+z���c�'����m<L?O��0��T�*��F����Y\�q��zE��
2s���>�̉O�z%�WU���P��<^a��#���W-	����+����g��% ���~h�����o�6_�8]�F�2{r���{�G�d����1!!�F�F>���{	��d��.����2S>��'_i�)�s"▰ &~J�3����)�~/�:�\�6���
�wX]C�u߳�B:q�Y��C�a��=�,ƚ�!�-�ɽ=K����|���)���(��}�fS^z��%T�`i���3:�r?�S:Xg�G�]��zSl�{D�:�:��_��옣/ng�ɐv���P��7��$�M�i�e��'![�R]�b����Q�b�.?1�R�l�������H] *u;C�5��-�P+���A#j��C�g�����v����3N��� G V9u���m>�쮿��|S��+1��8��X����'����ۘ4�{�K$��x�̛�Qj��`���W����@��X��F6j�5v]^���
���>$��u_�w��|�t�<U��u~����v��a��#��^ܷ��SL<M�B�w��FGy���{��T��%��C�M�l��zL�.���
��G7�	��S@C&Kz��԰����gr\��=���cy)��	8v����,��,�F�	ii*a+t���y���9��.e+N��h�E�s�\I����C�{�"n���2�0��*\�/��7�C�����(ū�$��2O�y]����5O������s�?���H�(�
���d���v�E��DJKh���Ա'1 �0fO�~=�����^�����0.��+�4��K/�1Tdb�+:T<%3<�G��]�y|p�ɡ��)l���ZR��;~ٵ<��tI]�o�6>.f�ϭ%��T����>Zc�;K�P`� )��*��詊g&B"�_����NQO�?T�$R<���*z���b���
�XYڴ�N�OS��,�5v���L- ��ZQCqlʕ֡�{���B8����Ġ���Z�Րie� ���{Q6kU�V�v����3u��Z3��#�˞��(����ߡ���+	nR�'J��N�F��ʙ��r@(a&��=]�m��7rmF�⣩Ԡ�\��ۣKZ�ݣ0l�r'������A��}yF �����6��	r��g\��/x��o5��bs�5� ߼�Ō�?E�-JO����Z���ٖOFq��]�m��Y&ۅ,\ʷǷ]�^_�l�6Z<�TF��u��8>���2�"F8Ml���X���r �q������������M.�����w���?*v^_f��Н�r=P�3���Iý�,1!v��(���c�fp�f���1��B~��W.�ॱ�AtM�Q�e��ټ�ڀ�c>\�|z�Ȱ��[m�j7M+J���� '�U������	��H>ե�>�Vֶ�Y˗�ZY8�p�!$.֩Li2��&(�A�;�k�z��aȗۘ�{�fR�¡"���i;� �:A��T����%�Fʿ��?ftN^Y����V6_��R���˄U���EC����T����f���HO�y�2a O
joX����y�(��#(�Lϊ=�d�CW�j|y�qo�\��(����G�U�8KJ�}d�m*O"�?��[���32�D,�ԁ��)e� ����2����m���\��p�,(���-��T���#��l�	s�/��������^��ӆ�M�7$}���Q�wۿ��͵?Yxk �Н��0��`�6Y�E��.�����QQ[_1~���L��섂�JP&Ł��9�)���Gj����ZW
�U�.�M��jG���j"��`@�e�[X)�.�5q����c��
Bb�2��]icߏ��]i��~FN)�,J$U{V@���r4�D��!�Jk��E�.[*� ���ߙ�f��=�p2BEmA�wH��c��M���B<����-��	0��c�����w�x
_�8K�pS����PH|�7]#��c_7-�W��\c�Y%�RKAU�ɟb]�^\��P������d�%��չ=����o�4�y��:�^�w����hm�JE&�*t�LJ���a�#P���[l 7�G'v�Zm��"�z�9vQ%��#�yf�i7���p�<Hd�;�E��$��%j�N�u2[ �{rT�3��ПSr@���b����.���U����,Φ����o��)]���CJ���� ��s��8
�	a����9��Z@2�
�sY-O8s[�}J�`CĊ���-�U�ut ��/]S�&u�I��픰B��́8l���G�םP$Jޘ&4�%� ��ΘJ��oPB�6��w$2E[�#�<c�����PE�>9�c�����.�VKG�L
�@�6�ivU:� ����R�ɓ�MH���� �[��s�iၔ8��~�ɤ� Q���ɷt^j.k�GD�֑�w1.�=&Jr�~n���~@�u0Ys���=I����"x��+y���mi�`��at�T*ᜌ��>bG6ґ���ύ��k-j�eF�U����
�S\���� A�B���K�Η��0�y;`}Hy���r1MBDzL��0iS�Ӏ@.a^�5��6�X%����	;*������-�Z�<��Q.[�Y��������-�j'��	>1t�Υ�z�O2��nS��Hn�#�T���^w��kå�a9��]��D�F�(�peX�n��
����D�`�qR��iJ��14C��瀝�dD��Z�#k,�/�8�xIU ���C�s��	�T�"z��>4�
���]X����r�k�G ��ֆ�����c�@�^�^S�V��c@oҫ;�Ԥ<uD̎���?̞�����SSg�vK�?Ċ��p i��'��odM�lKƏ���F�/���<n�	g�w���{�9�ہ�BF�>�����v�����El)���!J�~r�.�3f*p��w
'C[9�l����i�J�|��H�� �'�v6�z*'�B<� nF+��4,v���:;v95�h���K;G�����f�t@����iD-%�P���j�>g?�[1Y$B��\]�;���L?��Օ�ۙJ�P�2ĲT�ԩ�G�{���͒�G�.�%�:�ya~Q��sc���1���VR�i�5�V���n�!���|���'�׋1��Z�H�\��z�p<���Y+?(}N��U,�[�1ۨ�*��.&hHH�� ���i�ܾK��u'�0x�.�2uc���M��o��d��[l�Z����ƍ��M��G��&�`:�o88��(�\�|�#�*���x���C��k���Fͪ�[�����SB�ʹ�$��I@���e��߁�Xd�z��ÉZT�X�ۑA3(�t� ��3��PWB�r��}Og��P����Pe�d������|�����i������M��nb5�Q'������>�L1�1F/?hn�MT�x5�]�KT:����I����P��&��縈F|�Ɍ-X���o�Q�Hc�<,z�rRY���J�$�g�sR־>Kx�j��:�_�z������w���g�L�	���m��q"Ȯ��6�U�V��v��돶ڮ����9*u9L��\� �ƪ��u ���|��C���NK�*��R2��ޝ{��ʋ(u��S���`"�(�Ï��.W�T��tԀ��7vЬg�cx����&I'���6!�� ��|$�ٟ��L͕��ْ��MvDы˶ɾ��f����<l��R��+���\p.Uq��u��x����&�^��x�Y$\�O3�����{����Â?�s p_S��|�D��/S���80�43N���݉-��Gb�<��#_�dMhQI���D%;6��B����Y�-�ar���'e��q�D"_��f����qr�ӽv��
��V�)�����k����]DT�j
aA�$���!'HҷO��)&w���J�5�U�b�G����$cƨ�앋�5|f+/�Q
@�x�]\z�M�u��|F�
�&�_y1%��@�V���ʗد/o��L:�Q��;�Gbw�Z��Ѷ���Z���7f���]V��������Y@8��n������<�z����f���U�F優_�������oM���E�U���ªK�����.�����auZ�d=�2Y6�5�w(�A��>N�P�����CP^�p�,�D~���"��,�Z#c���nK#&<���ؑW�`+h�N��Þo�28+�RA��Qvb3�*y�������^!��X3X���RM�~�& ����A���*?�Y�W-����
zP�9�KM0��h���N� ��Ҥ�D�PO���R�%�S.���b�"�L���]�B�>�yPo�M�냹�G}?|���i[��۶��� `��B3�uG�����xx"��	q�di\��,z��7�gV+�j�J����5O4-	)�������gΈ�Ԑ���V����|�!�9��$Cm#����x�õ� �*wO��T�>?���H�(I[Z-L�j��*&�'�>0���: 2<�۶{���64�
��Y���u�S�G��z!U�`�ͷ�m�<!�-�1v��`�d�P�2�]Q�(���K��i0#�
!�:�''�!YHc�bt�+Ii�O�)�5�@�� -gG��(�R�4�F$�@��A�� ��d�^j  �`�T��2�X��>��\�%d��H�l�l`�6yhT��,�ӴG$�����OKMZ;��kW�r�݀C���8ܥZ�@�e�1����y �JO~� q�M_Cx-K�)4CdN�3��{|�R�.�����f���u��Y�u�S�	���@3?q�_��q�A
��}��ߙ��qӆ���*3=�zU�(�H&/��K1�N2f�ap�����%
�+c���uߓ5�	�,��?%�/�
��z�����|Ý����%��IϨ���'��&�1�)��i.|0|�`�s���n��d��{��*�"M�(�aOҝV;�O���Luo��2QJ�x��8�˧��w-���r^��;�D��jج�l��:�#�r�j�#����Q��.|a���S�k>IH$�EQ�U#��0�̍(�� x�M�8�>xڕ�D��Ƞ'���>��U��6��->�}��g}���(h�:�uJ�hG�y���`
[��x[������D�FI?;��%�Mz-wUv6e�±؈��TW����:ǻ}��i+�o�����ݨ���N��;<R$�/�q�uH%�Ҷ�^���%��G<�J�Z@�S�ڲ�x�w7��?z	9
�@��`Kȼ��.�^�[��Y�0<T_ɔ��ۖ�(S��E��#)s�-��߼�b1��^��O��"���Ba�x��%�~�$�q���r1� �t����`��h�Iƕ��k�����,���1Ђ}Qō��[3��I���a)n�br�y���N��R���>��!mm`�7��_=�a}����3"G��c4&$'w��dG~T��p��G�oj��)����d�����)�0�iZS�j~�'�;�������R�~�y�z��ҧ\;��f���4=�4/@+A��gn<�o߫8��U�_�ht5)T(��`���	h�\����11jhY��r�	�f�X����xԵ�r8��<C%d��K�Qm̉(�a>YC�����YtN���g�4a��3q������-Z�8�si���RpE=W���ֲY��%6�r��H���qoAv���Cj�Eby�j�Q
B���M04�@(�ښ��tY�%��tBk��¼���g���&]Or>����ۿp�� �~v�mCv��h9U0�T�ɰ���e��ҹL�J#q�~��+��;_|K�E"�w�����G�3�|�\����Lb�g�V���9�� �� ��"ʩwH�p�@ ܆f��yI���v)��)�ՠ�)e���C��T�7�eE��hO�R���Ne���2���h�Vh��|4����01ƂS�++^��Qs 
E�
y��F�A�,��h�g���j����]��'��ߍ}�c��kr"�	u$�٭����>�����J��#���b�j���cA�K&�/������J4�b��#d�(����r��bwQ)���
p.��qt����0�|x��Mg���I����g��/�P�\ZtJ��fޑ��Ԯ��
>ٗ�U��ƭ���gJ� R[r{���c�������c�%����[�G�:h��5�uÁe6w#�N�B�4�vV�oP�����u�Dfr�`��I<�0v����?j�'k�#�����<�t[�M�]f��ү�;��O-Z��X<Y��z�� ���O�IɄ���+P� E�D[.���Vy7��(�:�M��s�D�w<�z�̤~ӗ��9��j�e��0�l���o7$ M�FM	2z	/
��AG2��\S&S؆/tY�IM7���J�D��T������x�܁�)+2�-��b��u3ڦ�w`�"��"�~`�>I�^�#賄�zA�s����5�~�@���ҍ[ĸ)�P���
R�E}Y�d��;��5k\J�*�E(1;��sJJ�A1�iV�h�!��̺�4�z4�u۴�p7�%8-cn��E���5��#w��A��`\�x���M�(�� 	>>����'5��@�״c� @3����x�/I�	c�P#�]�r��B��I3��s��gm@#H�^>��Zd�9B^=�:2�� �B["뚎��B+�<-�5��FA�'�
9�"�W�\�ʻ��y�h���ī�dG�B��x"�j��F<h��0��8�6?o��u��eT�i��!B"�V��y�1�K&���X��$d�i�`��=���HL�b��;k�R�5�7g CS�I���?���HCWmd��fP�HO[�����D"�R}�X�`$0 �>%H��F�ZD����S������uJY��m�ѝzX���Z'��򾴒�"'���������a)8�5	�(j�@���d�k #�س'ﺙ��g2�*�f+��Q�$�n�շ����4�s��|��!tk`��R.�]?�N�.��8�)��B{��+]�D�ɘh��B�~�vgZ빵�r
g,����/�z�ZG ���)���h������59yx�V�����U�r�v�s�Id9�ѳvo?��q�7?�Z�֞�������3�X��I ������q)d�w�]��V��C
*$�k;^�T�#�e���U��/�x��hz����D�5�k��x���+���s�'��QQ��T>�5l�D���5��7��W�D�,�Ul�4�W�b��
��@��濚�;��j�l�����O�ù��^���l���z~����Q�w52Y��/��51�����ݭ�x�)[o�Gt�3d6K'>�i�m����Q�y\����ne{7W-�.`0�nz�OJQ�3<O�
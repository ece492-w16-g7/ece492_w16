��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d��p89��N������Dacf�o��!$��Y���*�#�`b�[2������T��Y�c��iN��iO4���7�xDF��������ʽH�_�l��2�ȿ!^vX����6�n ��]���,a��)�F$�IN��)��v���i�]��x{'7��H"Gp\��.V9���|���:�#�R����`���<Z(�|�4l�o&�hwM=�������Τ�@X��Ś�z��Vz�5v�.�+��d��I�0��t�{�[S��=m����eE�A:5��4=R��G��G��`�`M�E5��|<+�x��s⹸_�tx�R|l���&�:@,�ZRv�{wNз��4�zs ~�Z�
��0��`�.q���qT����ڎ1�Bn]�l�df�>�M]-�°��t�f��.Fo����5�?LbY<Vj(���K��=�
�ht2d�Uz㣢z|DC&�����c����h~��Oy�0���2���?�x:�u]L��#�ݷ�u_�y��d�f�jZ�[Q��2�y�����mxMu4�LV�+X<�CE�/�ۡ��A:J��^U���(l�V�W��٣�Ao�X;;��@�l� �M����H��p��]0�xKJU��ݗ�x�L��̄,�3�IW�
�G��슡�������]����@X[��5�I��Qt?D��x��O�53�>���G$o�X����׍�Њy�Z�8�4)8(;9�@��]��X�~�[ W����&�>CO��[	!��_��x�5��	�zB���N�&�LG����D������^~�UՔ-�Q�����q>L���r�I�<IC��-"�.��f��$L�S%��f���b�dr�V�{�X��q֒��F�Uх�z���MC�h8S}4p�}J������ �ϐ^�CP�h���Xsf^M�3�W��i��
��"wg�I��)��)�#����g�4��+yQl:5��b\��=z�0TF�����i�c�7S����q��J]$�[��l6k����IЊT�T�g��ߗ�Y�	p�����w
*/Z#�O�>��@m9��7�ϕ���L�-:�Yȧ�D����~�8���]{I��/8Y2bM���Sp�U��O*u�c�[bLJ���LT9��Wa�x9�o��=q�Y�4�9����Q�LN��֠!e��!S�E@��i-�!�w�����y�	�
^@��A$�F��")�8�$�bn�n���"cO\�\p��C*��yuv~�<9OS���_L?@�ҧ�{���;����L��t�p�>�#�C���Օi=���0�Q6�[���,b�a�&ěkŢ����T�skT�j/�/����H��-�L0Кi7�%�x�s�`w+�f*F�����p@a����!0J��:���C&��c��۝���#�8
�;O��nr)����	���HѼ^<�F��:aV����,������$��CV�u�hu�Y���=(�;�\��������Gփ*���7w5h�.�(���1@ƃ��K�O��
6 K��J/��>�PZ���X�M<�#���e����}	p��r1���f`��ܒ_>�L(g<��%��g�~�ݙ�UK��	Pm�v�R�#&N�� M�_]� r�,>����}sז
 �c�������B�G���?�N�'^!�W�g�-6<-"&�c���JZ�g�*��/5��G4�zD��f�E�w��[�v��n9h�$ꖧ�a�U�C���}��S��� 1��Қs8A�F�����*y	��Y?��b��9@��Z�sb������랰pD���θ��p\���1|-�XL��,8�뢱!�	P��GG�0�����O��@��{�O!D|�Y7A�yw%��ۚ�]�L�mѮ0�ד_��tZ���CG+�Xh�������}2���q��S�� W���E�י-{+���v���H ��qޚ��K��#�E�{o]�����sW��ڨ�<��P
�s�� �˄@���E���]͘�n���&�
�N��
sy�!i��R��LE	e��:�X��sPII\��]5�>��Zh��ט�77"B(e�=�,%��ާS�_CE]������К1x��;ѼH6�D)��"Mlu�zm=�UhD����v�|���?���A��0�#�z�J.�Af��O>���wE���}��1��3��5��� �����/�+m��p�֋��5�#���Іp�?9��4TL�î�ǩ��
�{A�C��<ɔ��3m7LǾ�m��Є�IY譋��D=^xq$ӇD��2뗄�%�'`]��>J]�No\g5�����Yq��l�s�iQ2H�;9������zV�;ح&3ȸ@��!� �f^ ���}!�KaK7�'�r	���S�ɩY��Q��KP� @��P����Ii�Q��}����<Re<"�%K���N�-Ȃ�6Î�ς8��MТ{��@�FM1p��X���ʡ�qu�R�Ϋe�y���}���z������f��@U��ʹ�~.>yN��G�eU�[��
�5/�W��O�~lL�����b�9f���{W}Њ@��KTT{x``�A߫�`>�ZX��`��DӺ�s�����(�������j7t�Fx�~^��J<Z�¥1膇������$���/Q1>y�x��&�B_��b��w�43Z�|�sj�cU��\��\�u�A4�e
�(��?f܀��^��'zRCb,/���ԧ�'on�IjKY^��FMZ��Z�
����f�o	m��� ���4�Ww� ��!�Ⱦ�����l��"ԔԱ.w�h@:A���D ���,`�?@0u��%$;��qP��IqEFO����	�/�mL�*<��m�����/�Aq��YZ̡ԓc���4Ḵp��Tg/�/Tx�>��P��m����cAh�|Ō�l�=�o8����}.��Eø5����g/.���g���5�	�~bi�מ��ѳ���t:(B+\B\@������aP�õ� ѯ�C/N�U���L�E���C/�t �eJ��ǂC�O��ro�3 �-[)E���<�q�+���l��J�������̏�#ݐ�U�9m��	D��t��Y<�I����b�t��P�F����D	�AW4�V'ϧ���⣓Or�Z�I�B�kL�KyxwU�����%:��p�����xT��PA<�ԕ�e
�G��fP�]dR��r��ުL#��"О�
ڏ�>.q��%��"���,��uC�Á�yDxF_��;�3 �da�ء����/Z�ӔpX���6s}�y��ש��.r9����jcϹ.K�4yT�� \�pk���I�X�I�.�	�_�Dԃd��H��n��)����:��>����Ķ�Qu��u�YGn���9�ւr�!_��,��� �̭��
��!�W�6G����@$1i�o|�pV�9��qj���Lg0�
:&�#K_�D3²��uk�h�ә��Yf7�soCh1�	]W��ب�8���2=1E#?�W,2:�'�y�Ň!4_Eƹ{��P�t,� ��
�ai�Mj�,8
�,Uý�������C���P�H5`_�����IC�)���P:	�@?�");n4��|U,������EJЯ*+�VظН1�g;���jV	�ѡ%~ٟ���k��5�J���*>������o8������2����7.��Ʉ��z��:��/Do���I\J ���hAq�edyO���8qAS���&�G��d�M�P�f@�}�I7�o�֯{�+���,M�D�S2�65BTE+��,;����:����{A]4��+�G�n��Oq[�¢��n�����ױ�F�)+Ns�(���3��y��ks�M�^�������0 gj��s��	&EK�3���c� ���i�)�IE��=��^	���]�(|���Zb@6����&�?-�K�ܗ��y���~����z0y&*�B�X���7&� �%ܼk���V��&� p��ˁq��u�ysA��V��c����c;�̄�]�Gw�!(�����vgAm���0�4?��(JW6!,	f���b���Q[>����n�$hezP�yk�m�H�- �
���}�$%����רBgu�؏�����gx�'9�M����a#��aH��0�/.Pj&v���j�	��i""�p��$���cɇb�^13|=��K��g~F�3��e�v� {�<�������%XO5�Q��Mo�X%��%�*�3Ҭ��NH�/�ַR���\j�|�}����2�;]+i�B��:Aiow�{�i��[P��L>������PhLBVC�� �c}c�V��7/�-��ur�8<eDܸ��TV��vTr8��bj?��� �����5�SaD+O��J�:�\2�U��}]�ȫ�HK�*��-/�?���]8�%��UW1�L��>��BZ�V�����?�R�Y����W�*y��>��V0`��j��,m󏟙��,r�����`2O,7yO���>�X�E\�.���T Pǭ���	F�o*ʑn�=B�4{Y��5����\~���`J���N�i��sި& t�j���*�ce��״1FيS�}2�����E"��.޴���i,�%%&��y��YH���R�沃gE����4�pe�4J?����f�����2��<�d��-��P�q7�l�$`�c�YH��x�2_r���׹��xlx�����<�^�"���ȿ�u�c}ٞ��%k.>���R���]M�c���̣�Hp�z!唯5�*���S�aF�!ޛ�C��8CL��Jn�;��
��A��=�����d��pP|�zO�v��Ƌ'q��:�	t*�ZrB�RA��(���h�7O,y��-�]�$r�+��z�c�9w?g(�t��6	����� ,�rh�Ԃ�r��0[�.�0��tf���-U>��N��3{��ˆ���p�x��ǟbad��.�w�D�r�0����y��\a��GR���3L�����)�1W]����w❈;<����eH��������]S��?@C9�7X�$b��yMQͫf��.����Jm`�ن^&v�Fe�������mSΐ�Z@W 2��§�җ���T��6Q8�순�(jz;C�� N,�#�&hܦ�7!5ߦ����M� �t(�V���׿�j!������U"3ً���x�Oƺ��G9S�k�d�9��k.�;��)��h%]�B���=�7�r��W:{�z^���U#��XuF�u��)�N��z�q[�5�7~��9�(�D�"nk]G�54^�M�p�	��o�')>�r�s�&V`T�/w�QE��7?���V��လp�CJZ����l ���k,_dAή�^~|�	o�)�
�1=�Ji�t�j顢#�,���V�]͜z2��T��O'��<�M����+e+������/b�CX7ÿɵ i����ٱI?�]7��BI�N��%b��kh^JB���N�������i5b�i9�k�T�=�@�E��N�@Z�~�P�:\CR�S
����@!i�cz'�1�q��D�(��t���11��"�B���Mgp��t�<�#y��kٔ4���N��g�)J���T�U_P� z�"��g+a�r��a60뺼�m���8��_��������@b�Zy,H:h�t�Oq!��g�,pwo�{s���R���Y�'�2��������^h��ߓ���T�`��u ��Ni?�4��Keܰ��Y	�π��`�C�-��~�ut�QH��X�t�v�fX�Z_��'P-��-�p�����c5ǥa����n��-�'
MOx��|�n�=Ng۾tͪY�=- �;6�!C��&��07��\	�c'�Xyt~�șP��i(l�6�M�(s��[A��֫�y�\.��x�h�S�7 }�jq.n��t��gK�a|�V�w�RJ"%qP��J��D�~�):�*��A�,��k���ܕ_7ƿ�<��O���vY�B��n�����/��e��H�f�Zk�l�����^X
_��B���X\��%x��^Y��{\�[�BI3T�B���ѳF.�, �o�#&� �DX͍���;���t݇����~�i��fhI�������-N�:1?n�W��
����+��>Q̳J��M�L�Ơi�2�����Y"�zj	z �/�s�p���h��χqz�Y�`_�,h$b ̕ʄm���T��7E�Q�MJ�}�;B���4Ġxn��*������Ig�f�������O*(C�q0���9B��9�W� 5��7@�T��y"�G@�jq\X���c��+�vN�(�OI�0|SY�i ��o�������7na�h�\u��_�H�Yl�G���0�PU�����a�r+zĨ��gy��#�E��[��	\&��'
dq|��k�e0JM�u��	���LԒ�"&���AI�#��겨�]W��G]J�]&���_���(�R`)zٲ�@<bJ1�Zۛ�I=�&�Q<��3^z��xEX~��a�3V�a�a��
��>�_��},zCg; ��B��ccd� ��y�1��|��F9��}-�G[�����G�L7�"�S5�Uz{�7 T��.}Lf�Z��-]~�l-�oM�%3k�.?K��Jh�����&��M���=�9`�C��2���Iz�\6K�|���@$����������x�Z<�}�@.��#ߣ>�!�TA�ˢ���7Չ�s��h�9��Ɓ����΁�X��#�`6wdő�H~�T�B������i��>�ﴅ��=l�(�CM?��q�����[���'*�ڵ���I4a�%x*49�"%v��ب�4�Q�0�sot��W�!����$��|��x��پ�H��SP{Ө1T�MILW�^B�~�`�*婥�/���p�����-���=�I�����!Q�&�r�"¾���Vt}&o�50�PQ��@<�'��ۓ� ƅ9��m�J���R�f�0�jQ���������	r��ϿO}(�#�)T�[l�BI��*֤B�OM�Y�֣R��W �f;� ���DQ)�v���$��a"�'��qk6�u�74��T9��"�["h[����m3݀u�T-,s�Q�Ij_��4.}�)���j��1�������W�ƌx;�����J�z0���^/9����n0�A������֐pHs@�4��2�Yk��"��[�{T0G�J�S�p�/�(qQ5���Y1$3Jj��� Uj�����U��y3���F=��#D|
ۃݺ�ࡪ�W؍��]yխ�r�v��r�x���ퟛ0W]k���, ¥����9�iZ���gCM���Av�xئr��Ì�"p?XQв�3����J�S�tF/��@��#�o��
��3�>�fBc��g�����ǝ,3��b:���� +V�z@�	�W�n�����ˀ���X�sάVg�bP�~�Z�?���c{�7��1��a�NW.Ӈai��^Ç�'���|��_�F��RziO��:�����<43�L9����c�dr�l�>=�57;��$[)�T���&�F�2�
�G��j)���y���,��@��Fej�'�p�"b]��喍?�M](�u_�V�2Q�a��r;|��	
��ʇ��	8�(�yI��mv�����==kH[���&� �K����<���l\\�jq��ߢ�=�#��&(<9��M�o-�� ����'*��v�|�]����X�*�w��;d�놐E��O�>�gp�g^	�|�[h��Y8�)�R?-���-jr��\�2�� �Ȉ���n="�1J$�d辆e^�-�e����n��Q��<>�� �RF��q�k��,�K~�Ps�t�ilO�����O乘����m5�a��KSi�ȷ5j�����E��@�mb�i��^0���tC*�g��s���h��5@�9N�h��\8B2�!�8�pIH>�{o�U@l�#x�݌&ŗ;"��g؞�bX�����ɠ��9U�r��~�k������1�M�s���a�a��)��|��7��`�wo��;��!j��䯮q�u�1�c�R���u�pC�� ���g��Qy��a��z ��{/���G7�PF�聎�qr/��P�* ���UBnYn꣊������j!s(3�2,b�5<H�Rג�!���c�Һ�Ν�HmS	.T�~�\�X�ޫ;@�tҝ��VK��C��Sf����d�s����n<V�
K���K��J&�5F��j2Nw��n`
������^���R@ԣ,�M��gIPǸ$�i�,{�8�jv��]�7��3[�߁n���[����vd��N��(�!%�	���"���U����t,�{d�� �>IM�w\޲���Q�AXlNH�_C���7zZyq��?�y6�w�*87E��� �ϯ�^ؗ��3�Ǫ�6��$UU+����/� �)��IQ�������C� ����Cm/F#��U��$��{Y&�f�|���j<u�S/θ�l P���p���b|u�va�b*�Mn�Q����|ג���$;�!�����U���fcc��j�a����fG��"��r�k{󆹩=EN�~ߕQ�S;w*��~RM<*�p�RdxTLE�c�o��f�������?l��AUw>�%1�jY�)OC��+D:���<���S�B��]�L���ɿ��a�ã�(e#7k(���B��2����d= �df"�9�Y�t��s�g�g�>�+��d{wU�+~:y�Rq��0��{*�C_=��7{��U<9@�`<�"��z��%�c,y�|��z7+�ˀiܞ�.b��y�T'�����T�Rj����������c�z���	�t�~Mu�)z��P�jYs�.j.��[v#��ʩ�({� ���Xy9M;��!XRb��L����뢌��j
>�� ֿy�俽��&A�$a��؜W���n�^+�k�/p�3�fM^~��!�Im�41����&��*,�rŀ�
������E EW��#k��aZR�+9�o�rϨ��3'�@���Np�f����1q��)��������_�B�V��Ss�'�辟UsĔ8�%��:
��ʷ��B̾,�U�-;�d��8�6���B���:��+`[��1����T�Uo}z�c�I��3��Hͦ��`21$S��b"����G�y�xR*� kWz���1R��0li���G��$���2o�AA}��өˤz�2nk�z��J)��_s�B� �d�r1��95��rC!y��}g��/c�E�B�2����0N ���J	nV�w���Xv���%<z�]�����)���m�����):C?�`�������x.(�z;�=�o_�O�pe�;�!�b����f{ɀf��D/��04��#��6L'��Y^λ�	O9�ǛF(���s#D��h��[��k�D�B�I���1�	o]���4����*κ���������g�d_
���Z4d
6p�Yc2aE�.Z�~WB\Ŏ�!K�إ"���{�:2�1��t��u)-�_w�|�V��T�i�Q����)徲&FHr�{'ɐb��1r���èf�����P�!��6Z��{�;���c���h�h��lS vu��t�+#E�K�6:;N��lux\h?�� Bj�ɏ'd��8Mg�%a��T{y���J��7���MdP�e�F�>+��n�͠�t��� �
�pn�����k�;Y�hu9���H��[�"G�����ݫ�t��L��G0ҷ�L���7��d��L�u��H/X)?7��6�6]:
6�0�z�������<ֹ���$�WL��#��e������a�8n��f���Yc�MBx�3��("�Z�l��DC���t����D_s)���Ky6*Dk��6�n�I��G7�=QQ�尃0���W�j<�pة��֕�����0-7 ��O����0?9���˨[�T}?�W6c��"��O8�T���Uli�������l1v������N�Z�~�Ylo�Fe�%���M��H�H%���ݣ����*J��N�j�Ox+�3Iw�_�I���1�Q4h�T]4�jDv�l:��4}�5�<`�S�`K2x�5APe$�,�R�o��bE�z����O�+�^/a}8�����"%�P��x�D����'�|Z�K]~�@�w\�#}���	�#�]1q���FVcڂbb�8���YeOn������<ŋ<�%l�zg�Jzx� m��F�r��U,Q�.�td�
���aC]e�}�y��$s�X'��+�WV��|�����Ek�u�h�v�p��<��Ä�lB嗎������>���-A�k���7sh}O{��d�{j�=w���FZR�G�V%��OoPw�μ gμC��B8�[�b�9_i�SR�S���C��BT˰T�N�L)v�ѳ��\d�����L�~O�:��|��8yc���_�!�4�_��	k���N`�/���	�^`{ڰ�ĭOډ���]J`^q��m����}�����\+�V�v��͙��#��'F,h#B4��y|US��Y��Պf����E�&ߣ�>������VS4J	-�q:�ٍa+��T�G\�����W��h��׾l+�8�1:q~}�βɥ�P�=G�J���������o %��i��P�#ΕTe6�$��b���}����z
���v�Ďu�W�4��+PJ�Nc`�*�@*fg:�ހهu��Ø��&"�H�y��c�wA���w�:�&��Z(�lbU��S��<="=Q%'���.!d�,��f����+f���C���2����SwKk��/�Ң^�[_vh6,��'[i\R��	p�޽�����xl^-WDZ2r�0*�V��m�L�ü��F��Q�ӇX�Z�3�dM�C�I����z/�kbeO��_!�'-�k�CS�$�����\�����1�����`0��@�Zv֝�9�֗�ʾݎ`���9��A`�T�@z���*�a�!����ODс���%�C�Xt[���R��N'LKwEc:j�*��80��k
a���wĠ/�̈��2�j�f)�c|#R�E�[���s]9L3�DϤm�ţ��a�z����?b�;%��؀��B�MWR
�B^�����[p��*C���E��B8�2��
�ၷ�ǆ��s�g�5<%�m�v2!ZI�!�1cD�� e�A�aq4�!��}đ�q#{��Hw��}'�E���5�x�&�_}X2��胵�'ء�� {˓葷u	�)��@QAn��g�0��D}��>��B��W'�Y&���B�h#���xq�ՆP���ҳ�N��O���y���ħBr�l�]�%Gj�R���g��� ���"�^����XV���1ug^�Yﮛ�̢�y���}�T�9m�F��D�$�	��%�ޖǓǶ�v)��a͊��H5�#��@�K���j���@�%f,�1��y� {�)��ك3E��c�sD��=%=�Ӳ������2�v��'?�������N�a5~��0�'���Q���\�徇�� J�)\�C9*=��S���9�K��σ��$�'�W�.���?��'����@%#�t1��9�G����T!�
B[�Q��2y�&���ܐ�OF4�D��Q�V���]
��-�)WF	-#�0r�5���*r�P<-�&��P��t��H@�V��UR4��s�/���/�q����8�A���C���"��\�JO�f�f���y�Z$��x9���@)Y�54���.wW�Q���)����QZ¡;p������\�Q'��W�_`P-��!YEq��ͬ3l�Z����3b8\���%��H�5�b���0kI)F2�z��К�Pvr�F�K��/|�~+�l��Y�iD�7�P�k�J�/���R��x�G^��s�����$�h	�0	Հ�k�Bf]�D��7F]ƶhh�Z��n��P}Z~UOKn�f�jQ�w�J�U|��w���ޣk�~j���q:!q����}N�2(-�S�2odC��4U�b������5ssC� -aa�8��5`�L���#�5/L��![�h(��a��2��a�&���]�c�>+�9#���/3�@���a ǝ��M7ؒ���ƣj�wA�~A�>�KYM��Sq�8,b:��I^djU�����B�;�1��W��v�=1k��_���K�9t��Ʒ6˴��S��Q~*��|H�Ę�(��$AP�>��2�z�NS����?;K!�2y�m���q�V��+�tʂC7��u�n����b
Z�ʅ\�K��.mLO�~�f�!
�I��_)GD�	��w.f�C�Od�^oyO��H@�1�#�QH0��on�C�tۀ9/������-��O��|q3���(��(� ���\���L�L��~�� X�J]��+�8\6�w����MM?�<�B��3�~��!��?���+
8�*����BNǁ�D�"��!�#��j��眮
��$.s

��"I3?�f�r~h5����<*k�cV����D��<U�^��MEY��ZW4~��>A*X.=�D������9_L�^dn䃹!{�=��o�'̯˸�[K'56[�3J�@�qb/�����ݷ�S}��f)�:ږCBpK
��w��\��-���2�E{�nk=���ߟ>�D�>����izG�@�g�+�����iYx��ٱ�3?Z�-�#�-�m�������i)��+����%��?+v�V�����ϖ�r���.2�9���0��X��5�U�{,aف��Q��bj�e�h�f"����6ϩd^E?%���Z�*�]�6�C����;�� �)����(�].Yc����޼f�!�!Y�XaKcd?�B������n�{ș�~Hc^��5�|U�Ù��m�x�qa���Al���_�Bg�.*CC�V�EF�G��D��}MC�J��x9��d�.�~U�<�A���p���ר�ԡmXo;l� �.�3,�D!�C�ϳ^�\e:�A6g���ܭ��L�#�����F��]1��d�&na���'�s�Mގˏ�-�����Ɨ�1��<��4�%t��?�:��W�	��~���5���-%
���G���z�����g'*�$	|Җ}KL�2�#J�G$���A��K��� ����?�\Li�rj�C)E0`����]��{�G��;F�{S��0F�)�g
��Y��[��rJ�*'�����g��Z�\�凓���c��.'����y�>'D^��1��c{ka���.���?�叢�A��V�rs>�4���h��*����&MOfޘQNq�KaN�u��#���+�Z�|�@`�"��n;�u����/�ǋx��=�+ hD/A�R�P3���)�ұ�����]���'�{�<Zl�=���nGj{B_��J2>`��{���Q��黱��@��C�"~f�U�[�
�z�I�k-��50	���Xz/<�<����#77� �0M�-V�[L��@1t��x�1�o�%�p����N�ssho�@q2���!�5�3��O^���=���`3�^�F_�����G�gZ�F�c5r]�%�|�5R۳���u���oΣ���%�6�a���3�4;�O�әs[�ɻJ��W��N��ߙ��#/E;)C'(�2
 x�dW�	sF>����& g=p'�ҿj*@az�dM6+ś��w%��W�K��[7�da�����Opg�����8/R� cO�
�i�$h���M�CsC��M�?���gC$J�_��ߝc�����Փ������YǛ&��N{�E57�d�>\4��r��d�6}��GH�əub�}� V��92�|mx����:H2Ue5:DQr��Vǣ��P��U�N����cx\Qwo�-ئ@�&S��)��W,�EР������JzS��~�>C5M���v��L�|e�Yf��nr���Ys>� w�
=1MO�?�sڳ�y�S������W�)�X�j�G M�,&��-A}��s>�{�S�7!��*��M�*��Z��֪�9��16X/�"��[�Ct��_�����Ef�;7؝F����Ы�[��H�2��y{#������Q���������@�(m�yO8���H#����b;��+��ٵ0�TZ׶.��d�q���{��iWdT�NuL��K�<���e�2A��q�`wm�[���1y��:��?�������/fD��)��`w�>�S�	u���\y���`�I�88����͵o��N�.ko�졯�\c�c��>Z�d�KTL4�GC�H��S�����pH9��Tn�DI��
q���mcb=����8�KSG��g]�QQ���H��z;`� ��8��ZpT�� ��\?a�5.��A��.v�X�6�j��+j�������A�� ��A��^в�����o��}s,�>�P��X"c�a��MƓHj
���s��0'� ����v盍h��Ċ�n#q�Rϰ�P��k���X�Z�uk>]<�Bǲ��L2��.��T���<ފ$��� R���aN��έڱ�Uj�6�A�i������Ml�ױ����_�m��5k?��w�0[�i:�[c�:duM�E��xs<χ�ܶ�5*R�w
�Fܮ4���8|��\��,*��%�1��e��#;FGQ�"mB|�s�C�
g�0���IB� V�(�V,r'Ⰴ��I�
�e�0���u���t
�!�@7U�)�� Q�yu�l��i��w�x�O�֨!��,��f�������?�#j;F9w\c�l6��R�?������U�7�S�P�x����4��[�����5�,QO_r�ף3)����(S�)mþ�G�^�*�"%��J��� �dWS�\�rD�ɭ!'�����c�0� ��!�������ޖ���(d�]�v9�DJ:��QJ6�2���U*#�:ᜯ
��_ៅ��ޜ�eM���y��9��~P�q�D�r��]a��H�ۍ7m����r���ŀ՘��]���[mk�;`�'m�ds��`>u��Gt�cj�{�G}����)g>�0�oLHw�zt�-�xG�m��(�`�%��]��
#�-}��sK�\��6�5�^̌%�iG�����.��1ϡ7�S�)2���9�j�,^����\க-�8+�(v��,���ԜnWx��^Ț?T�u�S�L���?ϭ~o�z�����h�����7#�KTA`���NS_/�^�E��g���RQ�!ڎ���R�����.�6�c���pT��eWdN)�*���{�=��/<<��k����|V4�� Dվ�]d_9)+7c5ޗ��3��"��Sr'v�զ�/���i��oɼ��J�Q|���d���|8��r���:!�-?�]��㦼���L��ZRht��i��9�9 ���Ӥ�-�jhʯ8��&u�#�P�B�P�Z���W�Zn��`}P�ˋJ)��n0+�z�'�(QK�}��C�g	�|�_H�ωR^�F�LYS�-�K��Y��ZIȊ�/��|�}���QP��e��dog��mf	Iю��/CQ:���ͥD�j�8�/�y��s̑�}�j�J�.�P�Yr�*{0hN��d����B2	!�]j����)���c��c!�i�s�rmB�s'zx:����GG{��F��t'�+��]f�KB\�AJ�jҦ�6��iz�
���M/P><c'������K�~Nf@wc˕1�Js�L*H�(�0�J��O�y��(�$�g*S[�c\94�;�@%�[����_�~�+̝�u?͠�"��0HH%e�ۨNr�V���8�� �H+q��h%�
FBp��5}/?�:҆�A ��d��7w�)l�|!���f�Q�.B��������|��ע�>�<!��+F�8+zM	`�._AVPFV��&d���'�k�g�a��_k^o�;��>-�)*ݕ�7��]����G>B4ը}�F�Z�dG7�?�՝"���;9pҗ��~4�f6 ���j959tz}W!�}��{\K:Sc`m�pF����3br�7�9�o�'����4��p�)e}@���9t9���q�i��
@]�=�Aй<���M(($Q8S���!��UZ�@6���������A|������Bý�T�fb�'�'�v���v�u��Ж�Mչ�t(��h�c���;X��	(x�mzb��	(�F�q9L2Q���|��i�t���0[�t��}�����]��U��*<ME�(���B���Q��߆���%|���Cm(0!I94���O��ػ%���=\g�=B05l��dD�&�ܵ���:҆G�Zh0�\�� D6�>t�גa��J��[�s�]˽�6�����s&��t'5
q_��`-����wl9d�*o��%k~�adGrmj2VV�t��0$6�j.�zC	�C����y����[��J�K��EA�Ç���}H��|g��I/�!��[e8���A���vM�
�Ҁ��UӬ1�)I��z���i5ū�A��;&���	0F� �����"ҵ���&{/�o��֚���[آ�,Y������*���ګ�3R};��;XR���+
�� �F�4��w{�	N=���iE:{#9z��J�7�{���!NA ��#ҔM��h"},!��2E�@7�嚎y�*��ĢA	��,ҭK��Ma:�� F��nʀ��tI��j��$�]�Tl�u~y��θV)/hs��O{�����|d����
���i&vUV��'��PP3c��Ta�W�$F`��7�B��=)7+���I�bb�{-p���`�#o�$>x38ߵ'�>?�����Mū�h,p�B�,��`� R�2Wˊ���̃�>u 7bΔ��]��Q�nE:Ŏ'��r�ɘ���:����6�ƢIkuWt�!�dv�����I�&��Q8_��`��`}��4N>��\TU.��>�~����Q\�gOL*m��5��x,<)k��/^��NLO�iEwMp���8,�'<&YhN�2n֍�iw�O�w��$�FX6�A��s�뷠�����|��7���IYXU@j�_�2���	x�Hv���xUF�{�L�TrY�xv�i��R~���:ԟ[���d��io�,J�zˢ�C"/n��jz�0�� �:��/������ˌW���0����p�%�H��$T�]�9�/�@)^l�c?}�к�?~��Իf��u�6G�V���
y����]G�&Ծ�Y3?�*b�N2k����nq����	��+n%��Ch�ɿ���K�R$��܌9�)���ʩ��y��4����@o'��a'[<s�M���W�4R�O����>���g�W�#���,"_��X.�i�Y��V�G��"	{���hG���E+Y��uU&����Ӛ����}�2 V+=��@ru�b�˕����5�xs!6��U�^�i���q�I��Ep�3&#�'n�r�� i��ї�RҸ�(��E�6(����3F����Zj-� [��0x�g�ܱV�m���ke~/�Z'aE����@d�� ���:R�d6yRy���{Y��F�<u+�G�&b�Ķ�-1�A�2G�1$XA�q@�e}�#����0��@��!h� �H��\H�)�?��J$�m���V��ڄ]��x6P�n��wڜ���g�g��ߴ	S�����
?�RO�m;t5�~QD|�#a4�����np,�ųԁ�2�x�F�H������s�І�_4h���v+A�{���!��?����9sF����;�������#��0���f�u�v2��ַjrQ-��k_�I��ĄNS���	�!Bh�I�yKT� ���>ᯂ oU�Z.�1?�w�����I�j��QO���4��L�P �*�l����u��$&v#�:a����'��#1�`�g,x�eXOF��De�O�.-@��+��/I�aN�H���?s%#��+R�lG��6ד�SZ����\u���PU�|� ��ox-��m��u2��%��A��P�E����T��f	�؏����>��]���k���}�7�I��z�ҍa0�V����.V����!�I]��rA%߈�[?�1"k�۲��l��Y28���ND+�K���7�������K��W��L�Vְ*���_}�1o�٠�kL��3���s?���U޵q���a�I �GL�������k���ǽO��X�4;���5Z���=h��I��p��6��i�����B/&2��ѯ���"켸�
>)��o�Y7R��& �?-�F�#>W����,��Gu�Uf��<w���q��� yFY�LjmU�A��bI-ʕ	m���Ĳ���9\̈́3��E���B�Y/X����m�s4=�����lZa/��t��1��t�J�T��\A��KBV	!�_�o�#�So5�B�/�������^��F�\���n��2�X����=耝��jNN�y�=gn����ԁhԔ'1GÐ�
�*�( �+�]�.ia�R��p����$�Z�k�d��J@����Q$8#���e�4�����n
d6���R��1GVX��R��a%r;[)� �������z��N\9��g����n��s��5�e-�<lzPC���X䷆�~��u ��e�[H���,6���ч����тm����\���/<��OAi������UgR���^#h���Zn ya
�m�c���������=(Hh��RW�'�gp屸�>!A��/s�r�9H����T��'�F��lS����?%�0�6x���O"��؂��*(b?:x�F6������ۮ� ���}�F����fx�w�]�ǚ�\	��f��Vj�ϦGd3��7?��V��u���l��@D,�psa��S==�=���x][�L��'������E4���2���v���.�3i;y��g��p������xJ�ڳ����8*�, ��9���Z#b�fd����f>n��{�~���ui ;f�f����(�ozP\����>��d��b�,�R �~��^8��W�Ł�e�����t�ݲ5b1�zд�]x�rr��T �C��sU~�2����v���7�M��x��QF�?Abw=�z.f���{/��&���a jM��bՋ�v�h�]<�<=�7����-\�C���A
+{Z�gO��z�"	ڧ��(*˒�3$��w��=�^)M�Y\g��I6��h���?�\8�l��~�P��������6�+S[���i��&��b�&�հN��h��Mw;x�E��VX0(��
�.���a��*�&���Ա��~���;��5��m���9����R@�����7l���A�SSug�����H/�4���[kQ��0�|�;Ap�h#4�f���E�b�;Y=A��b�ln��f�ߩc�^�J��_s��:�i��Ђ&��V0m�٨��r���_g;��^+��Pa��P,	���E�v�9�M��]E����>t��֍+����p����2��m0b�>�e̓ÁN�ښ$W����\鞓8�L*x��s��U�`��s�Z�pAt�����=�K�}���{�a"@�fl�`�{�������0��&B�Gb��i���,���	� ����u>{��	IG��C�lp�Uvٷ/��W\�cC���7�nf�nN�7���L��!I�"{aɏ�TO�9�$���Ѵ�� ���f@�u���ۿ?]�G��
�IP��_*�O�Lp����?�7LE�y_l����>��i�4r���r��?i��������6&��*L�7M����es� xy0���]9O,I9�cq�?��=;+�]n!Vu��,�R�O-p��5G6�'�'�"_^;�otV,ʬs�ub�b9s��Ҫ��ذ�{��o��r�C@��~.m�}��]ѨW=�g����3�<�`��h���2�t�9A��-�2����m��#�hqf^$RT�DA�NW1��cƮ��*�*��:��LJ2#�5ǋ>i)cpyZд`��湖Ǭ,]̀�ǐx�G;D����U����$i�<-�$��?{�$�P��������3S:�15T���k�1=Db˦�g��?W��3�1y���3��67���Qn%�"�rNƖ3�I=/��u�bV�.�Pgƃ��pα��Bƺ^"�^��X��"�%ޓ����1^�ƫK;l�������鯾a�,��w�4V�""��?��&�k�:�K������q�M��i@�lc��Zʫ�K��B>�~�������;E���GSW��e���V�t|9F3�,a4U�-̄�Q	�O���3�`Q_�@%�fL��+������L"���%/���i u>���g�{𪽶1lQU��-��;2��zu���ǩ���FP�8~���Z3���n�w��������<p�{k-_�������T�"���.����
�װ��
�^x]3�A�O.G�A��s��o` ��2ˇv_�y�[_���e�i�~���k��e���Rt]��c��(?Ã_�Bh�-8���{e_�6� |�v@�m$�2Ud2�_�H�݊|N�-�A����@�(�(G�ط���sT�1dނ����T�sAف���2n����k�I��sC�	��Kb8'2��E���wn��7H[z3��s	�}5�D�}��TUpBz�U�-����	F����J3W�}hl�Y��[Mٯ���~#��QrH��5�/�����K�5���g�j�����c�|:����TP�Cl�ZJylՋ)Q�lo�Ҕ���f�`cm�#�����B��EHd([�-P"䬧��:�s�
��|�QkFp�k]�k=&0eگ���'��j����WU�[l�č2����v�هH��E�}��u��h��>H��M�C+��"N3�W�i�.짟����(�����^@*���)��Зzh���[1������M���{��H� 
��:�N���(K 6�rd�,�yz��
���]�/�"�]�L{�1��7�LJu���t�z[f+�x�.һW
��H��*�J�� �&a�yT�[�{MEzޘnQ��`�w�ݑ�ؕ�h�����0�:��1�w�����%*V�爼ӱӁt#�v��֣\�]֕�x6�@�O�*������\c�Ig��*9��դC��&���P�c�r3�^���W�sL�=zĤ��N��H�K�Q�v7y�(�8Q��)vDqR�9������(��ƙB��\>GM�Ct*c�|mg*\ڿ���tE�gt�#�oj9��r4q�r�X3�a��ډ�o�ԛ�C��2��~��\�3�DRoq�ȏ��=��TY��s*�6n��@��
��BON��ٔ۴�j����KT���p�ҙ�p��~r� ?.�m�`�B�$DP�s���x=�ܒ�����s`f-�ߺH�S��YjME�6e�&��O:��NE�#&�	U�nLqJ��(��ɔ�j-g��4wc�.�z�u���R#'0d�k!���R���n���imF�����X�
3{)M��J`��j���c0��w�d��D�����{���/y�����`�8~�f�<�έ{M=�^��У�����kS�^�[��~b�ɳ��A���t�� �B1ܟ���o���N>����\�~?q-�r.�8sы��	��Vl.f�������y�A�Z���gm�Hޒ��$)b�66�Z��ۓ���zuNM�3��r���lk�[�kK�?�(��<û�Xn�h��8F�L�-�/ʮ�A��#�V���n��s�F?�Q��87Uک�WgS���D;i8ϓ!C1	a�e�A$62��KO	p> �'��{1%�ٯ,JM�����ȷ�P��˘��G�~����������ʼ�I㵖B��2�r���O�7O^�q�����n�l�b}��[D���`�Cu�å�H�BP��S�gdO�'�܆Y��F�����hu2C
/�_��֚�=�D�Ҷ�c�(�5�u��	�ۮ�6�c�;Al G�,��1� 64��r����J��a���~��j��pz��sY%�c&gM��"�@���'�6\4�ᤙ�'�'���s�S
&[p�� " ����Tx����?Z�b�(U0C5�pYT�0gun���0�;ߏS�SN ����n�4R2���%���&��B�&�)O]_	V��G<cl���S>�
��4�w� *\� �,a�˯	�L1u�?Q�w��C,�Ę4�<�q ����Nu��!���p��m��Q���7/7^:��5���C>�i��}�Y�^��^�?�&��;-w�ʨC�Lܘ�Cg曠\
#10�ԍU��s�F���[ŰQX��c�>g��~3W��Y��︡���c7�.���\�fɳ��ҙRM!ta	����Sc��kZ��LR���c��Y�'kiM�_�����媨�����fk���S�!�X<����$�;��Ԁ�X��=>}r�>�NƆN�Q$��پ�!TNU��'VH���%��{e
��&�ٽ��������2R�Ӂ_C��V�8�맦�u�
��8m..I+n"�=S�l0��^NȀ\˫� ���C����a���f	_�Y�� kt:Z�4>]�Z��.����7Ɔ|Cl�9 y"
,~9�2�^��u_k���"f}j�Fp������ǚF �x��2޸�+=���i�A]����n�����յE�.ϻfg��{�Yݰ �6˳�546!�мG�O�z��>;2��'�����+�$wx�ܪp�TGP����v�R�,YK�����=/�����gh?X1��ow���g��
Q�����3�p]
&������D!�������8`�>fI�Ct��&WZ�K�����b�����'�i�m���,eS"���N�� -�ϡ�y��c��U�f4�Ja�m�7�i����<��s۔�ɳ�4&c��j�0A�_ ?��F����dI~EU�f�=����~J�4�N�����ǵs���2�1�W�������l��zN�6	gs 6�d�#��|��j�A�?u� �B����O����~*��Y[Yy�qO!���\�D5��|J~ށhxh����ֵ�_��7��=c˞̉�p�XM�x�/ip�Z����"mI��P��ك�z����_�s�����[~�gS^%�b�"�q*�؛e�\�W�VG��-�? /�����4�hb��c 
@^&E^@�˞�}~�b#�h8��pd��&���lA���uoc2�[8��������s�`W����ٖ�Stn�'4�E��+��R�ƨ�(I?��7,�x�QD@�DTu{�h��k�6�-�!�/��a�a��l����VN?�sRd�K�R�i^���WK��G���N�L����$Q��b-+fgj]oɽ\�&Wݪͽ�X�fZ|v��-��Z����mQ�!�W����U`���է^���YU��P�-}�ֶ��!E�6j��}��Q��H���y󘘢���(�)�C	�cci�H!��4�̅�@�����{�%å�(��� ���E�YX�Ԙu��:��{��p���������o�>5C�UsA��m�6eß��W��ei��HD~�s��8F�|8�|�Az[�͸�<
ċ<$A�6ƾ�u���tH�� ��,~�=}�sj��~���K���7aFn�j�K�%ю��u#�ܰx���qN�/��O탉�U��Cjjᙝ
G�-���xm�"�\!�E�i�x�£X�wiH�*X����c�j�]?/^"�Q���?ӢoT��b�����5�Bٚ�T2��u!g�� ���F��@DkE�H2�+���{�����0 h�N������2ǣ�#qBM�M;�K�C�*c�&�"ҺD!L.��4�6v?� ��j��k��PMG<z�c�w �5�J?��P���m /�%��0͸��{�G��Qo�����a�>�0GT|���e�ag҇/g�
�pL�%	�7gq�m��h6I4���@ӡ���P�rL�W{������a���1F����IY�� �>���z��wA��t�	��%���Z���u��3�4�<����5���xN(#uл`SpL�E"�Og��U�>��l|z�7�����O�p��Y��ΚhjdAkf	���"W�^�w?S|D��b}p,�f��>Ms�đȃ^>[��U����f�O�8�(7�6K^yПJD-�MΆٷU���x&{d�`�n�e��3Wp�p8/�n�+�8�ut�ѐz�Qs��(M*\��tM���ߢu�x�w������(�t�=�6͟Q��;#��D��I=���^aM����3Q;��q��]�Dm��vi'ŏ�삧N���#N���G2���7%k"��?o����������D5~������S�X?��G2q�0�K����ޜ��3�a�����F�j��V���G���Q��Ó��ặ���]hzd���B�>��Swx���x)mƣ#��RT�q�1A���M�r�`�$�#�|h��|'�?w19�K��H~Zk�Yc%O�O��Y�M�b�b�!��!hg��*�"�G�};Ȫ3U��~W�ױ9Ȇ;����ȧעt�	��'[z3$���3�?ބM^�u�kّ�v�+�w�r�A����i�o��	_;��9x�JH�[4�X.]F�y~tKk�g[WL3���a�#<�[��6�b��e�f�&��7f�?"K�k�e$�VO *��d�^1�0p�I��źN���=�<H/"z�[U��ٟ��7J������,@V���P��L���|"Ɩ�)�J`gjIrMi}�Ɏ��~�5:S_�O���o��!�Bk�߂�_�ӚP�Ό��ޑA�ӂrfs�ϖ4���ݫ�rjk4\�ZK��[�H��b)5�2�`�)�J�H"�Hّ���s�fY��b�~�+��n����ܱ^��T�.���?��a�ӊ� &-�{�� Dɬ^�"���Q��\���#���	�ϫ3þ��ڦ���7��>K�w�����.-�o5C�?��ֶ�ʪa}�9`�$|��7xb���,���X��.��gi��EL��"o�<�ԣ(E�6_ހ"�b��`��{�ڌG��v�=��F�0�Y�0��ƛ[�c��I�mi5E~T���fe�@��K�-�e�3
[ E^����W�ptӃ��e9��0ɿ��t��ɽ����7�eW3��Q�;ح�'�������7$�s?�$V���@���r���Ǔ��f_�h[?/����t4�'xP�$`D%�R���`�Ј�5Et߰��շn%F[L5nE�	�����:��SCT���إ��.4~ׁ�$���G� {�ګ��v�z�X�>z�ޭ0�|��4�w����y[�<<�:��]���&B��+
��3��乼�u��,u�W�=�e�d��mN�%�(�L4��n ��?i���)b�.�~R-���a��b�L���������E����9I�M5��!�i��	���Tűb#:Ǭe�)Nж�	�	5$쪟��J�
魈���BV�������8le�>wJ�z^G�Ve���[�]6��4�1�嚵ǘ�n���܆=�%�N�&�>�p��G2�4���P?w�ώ�t-��:^K���vl?H���%�H�-v�E��-����8��2k�$�.ݲ.��f�^��I4��4�-�r��)o�e3�qW鐂h�Qc���q\l֩����Q��w2�	��Pۻ��PZ}}�]M&�SNw�})�ۀ�;��ͥ�(�l�O5�/�!a�/�I���l�o��m��a&��sS<e�2U�P|`��#��N�nx@͕$��XE��_pqH>$�����']p7($I�}�9�;�*g�"r�1����:@;��H��{a�1����k5��i�"�i�����������to��<��V�>�����X���}~�ˉ�Um4�73&�(/a5�5/	��%���`�TT��NnK(Ԍt����5Ȕ"�nv]�WW!w��l�t��m�-87���ǋz��0�4������	����g�~xjk�����6�6���a������1d�P��j�Im~��W��� �W{�p��K6z)_� f��RCf���=�Y�1C4_%�t�+���x��v��,+ކ�1����qT��V�p���Aa4**]o�8�K���`���T�ԛ��NfE�� ��,���b���5��R�Lv��5�{pj;��5*��	|p���p-��h}	�g�8��@��a�!��ɧ7ib��a���a@g-��]�A�3ϟ������G�vC#=v8ZDyޠ"��$�-��T�A~Q��b���d+b-�`~D�:E"Tr�4ƒ�` �E��Q�^P-�"��&�A�\;ʿ�81}�n�7pO�
%��@�~��.��
�G5ET�n�3��Q]���s�5[���Q��������C���[a�;4 bey�zr
'X'��!{u�!�[��Gc;�[���������O�4�dfO%6���Ʊ�f�W͂����'�	�e�㠷��4�2��!W���<���'�5�Ҭ���5Y,���g�������١��a�gO�k�ME>!��{.�'IkZΰ̌�,�z��>UT�������`H�o����G}T��,�?z�6�SԗYS��g�j��|�ih��m?��S�	?�1���lh�.�ڊ�+�܂����aj��`���=E&N8ﱐ'k�vǰ�b���u3��H��s��%��N%���Y
�(��7�w0��l=:�;�D%��8��U�i��҄�փ�� ǟ �h�򺽼%rol�[�k�#@��q������ǭ ��b2��تI������A����D�3�#�~>�d_~7To�z50�y&��m[/���d�"���\VB���: ^i��%n�����J��ل�*]���_�/�+�ǹ��K��|J�'��0�������6=�2�r�ě�%�i���[�`�Y�%䝪�5�0���fh��8w�}�:&%�;�hx1�L4��]���u�$����C����H��m/1�
�iܙn��%�,�i���I*r�n&�A�v��#�͋� m�v��Kg�0�9�W�ʤ�(���rۃa�BHV�y�4�T�|�׸�Zd�!E����r�� '����7ƴsȫ:AI_$*c��/�	0_���:�=�Mj�aX-$�݂A�v����@�<T�i�Ff�t��V�d����?q�vr�J���E?�7������P$w�������!�����џmK���I@���§Q�x��qs�������(O��|�s�w �3m\Ye-6l���3?ٳ��l#�R���B���뉗t�'=k8/���s!�b�p�n�MGWA�ȴ���4�i
���I)�X��h;���ң�<�Il(R@�Mxҍ��NEG���[�A���!��	A��X�|(�I��� Sn��oL\K, -<kG"��3M?�����竳�5�Vt��ހ�����0�8$�_�;�Kɮ����R+!��rqWĪ;�tl����o���b+��ɳ�O�r�5`?�ʜ>������C���W�*�ۿ��5S�A�S�36��������=�E����i!g^N��a�ݮ�FV��ڦXo��D�Yp��E��n{�͋gJ�N�O�H�&��c1!pPHD�!+�m�5�*ڛU��_�C$�wq�+7`(
-�T'@ ��%kӎel�PCE�0{�;n�X(C�J\���	��&J���\{4}q�ca����OTp񑕓�KB۶�N��`ALҵ8��Lr��@�
N�&��jr%t-;�Z�psezaZl�(r��
���sf�����(|�<q.ɂC���}��!���%���T.�� �hb]hys��Џ.4�"�~Ʈgi� 2e�-��"��>[P\����$]�N߃���/V��R����v�q��]B1�����3����D�b�3h�Z�A�#QV�H0\L�����">v9/��E|�y���І����Ruj����Z�[��`r`�����%�n��me!��6���'��b��i>�<<�м
�;�8�Wu��KTτ�
���a훔���!�D�:�
��4xMd��5��QHe�;�3����)�\+��Z� ��_��c��>B1�I����uX0�.ca���EY�c��ag�d��}@�����g0iǉ��ڡr���]H$�hfY�<�-�����p̀�g��W�/Z�Qu�d��>,��p�z��Fב�	��%�����7�3 ~B��&+����o����z�B��1m��7y.�N�KgG⸠�Uݕֺ��:=�ۮ�=��>9l7r(P����B��A$�v��:�g*�/:k�3Y�L�P^���i�Ktba�����j���Q�����OkJ|�щ2FF�X��V��x�z�jy�n��� �%�Q`�ED?4��㕕���o�^���sglDIuR��p}��e�J��V��ӌUrU:-�Z" ���v�q�|bv��G`�XF�<��l�����¾|&��[>s<�g�*�:*$�{Jl+�dr���!6p�7��b��Ԣ#m��p�?�))��f�uz"�R.ߖ�"��[Bb����k�/�]�}vS�w��`�Y���d�^��w�q-r�S@�����*be(W|�Y������<�`h��j�]u���Sbq��W����LMs���,���w�b��uºh�����/Ŧ$��x'��j�%��n���TL��8�B��IGOmi ��E�r�A��C��>4�:WkG�pa� !��1�1��O(�J�M��v(���tL��Hc�<�޽���Չf�1:�ia$��J4�'1����^�5�bʢ�,d�l�}�(� y��|i����VF f��%G�9٢[��@�<ƇqRУ+��\/����w���x��ꋧ��.v� `Z�x*��v������Y��"Z9%!j:S������!C�b����l3G�Őh*ѹ;�N0e� X{c���_l�~�c�#�+"{E��T1��/q���-�6��S6��w�������$j�v*:���+��S��!:ڰ�'$�K��@��'�]�H�P%�N��ؕ�? ����+6(���:���|����3!�y��T�ہ |����p"W��ܲ߀@���͕��<B4��=v�'>�J�]��r��H�Hv��ETdZ7�u����)`���	��[Z<l�R���%��4-�/cTu��_�%U���y�,o���_��*g�4�Ӛ�0G�XM7S���1ti�66�_&��#��)/��1��Q9\9��x���#�^X?|5B����X��M��?h������b�����4��C�����J��=�bIV��9Is"{֛��U��?�h2���z�h�|���GHʬs����X�T�p�#��&�e6���6�-
�t9�<��ˁ��%�O9~��!,p��e8S)J�a �<Pvr�I|���Ǭ�s̶�G�A�׾�sj��y?�B�����&����;$*�?Ѿ�â	4�z��e~�� Y��s���2�e�HB�T�3���K��/��o�ZR�,��>��� 8�� ��S���� ���Y#�#� b��R���$@���uH��8tϴ��!؇�3�������Σ"����J��v��ƶE2Z���t9Ф�2T�1�w��D��Ͻ%X����}]�pOD��d�'-+��ܧwjz�0Vl��~�[?�u��sȶ��n�y7�}�w��"�5Vt��x�����ԥ�e����=����"��*9�2�?)�??O��^'�{��#�	�
����O�8x;��zID���!�e���밴-H�jo�����6�0�K!�S��ԇyva?:`)�N�Ŭ�QTG�M��g-S����doI8ҧ-�G�F�jغ�͟��10�`���)�C7N���_�%/�ʕ�,�t�֜�FшD�
X���E��l�8��.͹�q#���:Gi
�/D��)�,ku�_%��RD�K'a�,,RZ&���K���7�A. r<���zG��x=���0Cdj=��8�5A~=��A�J*�.F(�S�s#0��)�AT���dexz�j1��PG�)�����T�-���ڹj|o��BfBmW %�E"	Z�g�����HU���2�8��7o$�����-�ͷ�i�K�j��	���6:~_≒*gix��g����Ʀ��'�|Ұ�<�~�zb��3� ��|�3�T�w�=Mi�Qo�ǩ��Y����I)����l�?zq*� �V�v���++z����b�������a�h��]�{r^`��+��J>������~Z�Vf�[�YP+u���pmJP�#m�ɳJ�W׈K|E �`�Қ�Ekp����(�/d{��~ "|l�V	i�����J�i~,�˚���v�	9��n�Q:lɏpR�t%��4c�$r�� �t��1=�053H��8g};of�t��4�Jco�e���5�A����� "��	s��Ұ�Z�6m���v��׿��	jjQf�ƼF[��Z�~��w�jJ�9(�m��7��ͺ7��t�m|�$ '���H��ju���J���1�t>�~j�eW����;l��.$�՚$g�A���-��ϵ�G��p���=��j���Ү�v}��J��&�b���p
ת�&���N^��f���.�Y`�M��1|Yܐ�_���qSG5J��.m`��¯*ͺ�_u�^��o��-}`�<t����Q���D�;K$aNc�3�,���$������U�fI^d߁:_�֪�f�YSl !_~Ů1� ����PkN7Y���2j�/0[S��/�^T�-�_��-
�v6O͋O"�d�}���훢?���'w�G�D7�����������n
SR{��](�^���ٽ��UʚU�?4�j�	bff�p�g�iQ�df����j��9=��Z߭]!�ӂ�����b��B ����;�Ც��X����6_���|�|����ӌ���@���3BC|b+"���RKo��Dw��l��!'a�W����>�п*�My��f�/�_Zs����Hy���� ӣK�@9P�P����@��_ס����W�ᰬL�]w,t����r���.⮜��҄�B�F�m(#�j��+���?ѡ���c���zT��n�Џ�tP���ڐl�O�v:����V��jIe�M��Fvk����Xʎ�*��|WDy��w,�nuA�c�[&�[��)�$���Lw��u������ԫ�p�9<$�҅I��yf��d�"/��ˁ�'8��P�O|<��q���S�s�9`��	e�������u�EW����Vw�������=�g�F9y�E�l
�-R�������3��M|��C��Bc���Z��s/���|!��^c<�`�G�i��������͠��p��u�����@��ʐGX�����������n�'��psV�d�:˯%@��� �B�t�.��Rg%υeAwUu�~���g����E�/ʨ9�ŭ��`o	i�	T �ޟ��~bYi�z��^�؆��ڮ����QG��(��37�u���vϿr�	��O���9� _D�M>������W!��-VVF�&�Ҟv?A�^�5�HH��4@#����4�m-�ha����[�DҮ�0Q+�w�.��K�@�x�����6���
��a&J�'6~�jU���+�w�r�"��Hl�W�_�#��?0]�ղ{�_e0��׋�o�L["8�#At`
"��x|�6JwUM�3�E��&w&�ko�u��y%ֆ[������݃.@ɾC����	
tu��I��n�T����HIV2���A�h,���{��D/C�
�8�d�1�	,:��j304�Mh���潀��ʄL�jj�4-����VpL��s-���,l���֔XKͯ��k�}���m<Z������y^�U���;á"��g$q~��N�%�����D_��cAa�n"�#hd����<i�-դ4{�I9��ηh��̑{���H��x��c>@�S�Ԋ��6� :$cT��A������b��� _��}�<�j�.1�B�kb�^����T@�9�N�������N��n:��Em=��:�T�R���.���a���@���ryȻ�=C��0.��R���0�q��yz����f曂U��g��\r�=T�����?W�YY�ٱ���UN�R�g��X0��}M�B��j�8���g�H��ēñ ��,a��c\k��Oqʫ܎ý!�_kT���ŭq9l���xw����*�3�U�^0��Gdo��K��aM�Q����eZ�ty��}�����C'��1�=��w	�+��;!w2��}_�pϲqP?�������thTe�}۠2fH��1�"��#���V-����$g?��T4�oX�
琑4��˲�!��4<�
�����	�!��M���ʧ�(g�W鷽�˓K?mu���;����Y�a�1���6��%-K�U��Vw�'��v��
�
|�վ���ۦ��_����B焻e�7_�^�EI��7�eS�k?����� �_ n�-����D7�|\L`�?տ�v��0P��c��m��}��Mٛ 8��o-�:��[�<���9s]�"֑��?�����+�/WO+H]�f^�,��z
�-5�d��xn`q�FT�70�2�3��Z������-i�S%�X-�M�_{�A��0qْ!�$:MqQA�W_YpcS�}|׊��	�>�6ގ�߅�����ŉ�d2\�����$�C.���g���f�%|{�]CN6�X�f!�c��:幘���	1<�Da��<��T��W~�8Ă��q8LztRˮ�����	[i�;u�x(��4�"���5��Ҙ}͸L��x�
)
e�wQ.4XGp�������:Ut�K彶3����A�:�Q�.�~�Ef$�OH����	����=���~�@h�|LK�۟�����CD�XqЧs̵�͗�!YP�T�p�7P�D �M�\�[�33��d��E-��<�&�pU�Y�DCJ$�(PW�B�e�4���,m�	��Q�/�s"~����v�6;L;��1�׿���c�~�^�ʃ���(ux*ٿ��@q��4���F��U�z83�**7F��(��G����� .��Ғ�|l��9��h������a7�pqR( S�D�@�[�������)��fG:'Lr���L�9�����<�=�����r�%�M�D^k]d-��~ݮE(rjD��c�=Yv���%�{�ǱO�P�r'$w�Q���ۮ-�P��ϕ
�=��^�6g$�},������F@�h�_H�sϣ���G�B��IW-�~�y�u� ]I��a�o�wX�r�������8�Y���^>��R�81��Od�!�(u�ʫ���"�6z��l���K�U�|
�]�؂�%�/�\�%-��>_��c�('k!Q����z�iIo|���I��H�e;��N.ߡ�ȩTY �SY1�f�pbi�����D4���;��.psb��=����̜�r���!7���ƾ��B��%^ʣS��4a�1�`�!qJ����BkP�ViF[ا���~��9��y���w~��U���Q� J��N�ԉ�~[�5ym���MK��{��|��Hew��V��6i!)���>�x�"5'�;q��&n�o�b�o�*�|���f�~�on�_�"x?�2va<�N|pa[�k~K��ˀ¯�,PĎ^�w���49n�}j��,<h����l�X�?T���N�^�ƥfa��qg_"�'��$��i�Q����7�e�#n�������� � �Ӛ>��6��)�'���0"��Gw�N�Mkq�C`�)f��ι�,�^��'�����i��S��e��;'G\�Y�h$�6=�;8��1�3��}C�"�,d��~�p��F����S��8��و�v���.���3�K��b_�S#:ȇ4�~�R��C�oLe�O���#ݯ���h�x~�Ah��4�Ǿ@f���&�`l�|z�|uK����̓0'�.���~>�^c�^�o�f�_+�|=HMG"_���c�g��{^���&送�6S�{O�#��;�0���d+�"�xq��Tz �!/��D.k�tS=�bN^�99�DA�u�QJc�������1�6
��j��^,L�d��X�@�L����B���脓��s�fWS�Eatee!����j�J��(,�p�Z.�P�M�a�|{���_�h��u�ǫ[ˣ��r�D���f�g,J��wqD�md�
���M��N��{"�~���,PR6��y���b-���Y�!�`[�D��WB������A�ۍLv˷�pL��בG��0�(��������>j�DGI�Xy#�W��G ��~@��)-)�	nk��<i޸��P��uO�˾�.f-hJ�AT�Lg;&u��˟(JF��{7�sy)����<Z��J>F:ҷU�y~KJ��Q�_�4'8�8�ٔ,ِG}���+�ܭ�>�\�J_���4�%�?����7S,n�m�)`�W?��C�����(?������H���&�Z&V�҆z&� c[)��:���`tE��b+sε(��#y&�z:���be�s/�:����5Y�	���u%nT�N��K5�Ts��H
Ǳ�C�����{rI�3fٔ����8��o�5ރ,|���
r@�;=��0�z &�u�4����%D[�_�'H��֛ n�*Ѣ).�( �S����&ӏk�>���W�;xm&
��,7�*}(��?C|6s'��3�����ɴ�$��tթ��ݙy�O

9]4�،�)�¯����g��8N��_����W%Jz}ZSi\���$ƬF���\�����^�����C�f��;�����Rl��eʫiɢ�q���)n4{+���&�P���ZF�qeo&��t��QM�!��)���i��K���6�C�P2���ǴH��+^���o3
���W��>�$�$��[c?���ڤi`Uy[�\�wS�y蹑N��~xJ��ǆyAaCEh�c�^1P�W��dG����������kW�ny��w�.�����S>�l��j(.�K��I����EQS�h���A�r�ki��T����:�3�4{�$��`����@�l��m�W��ʨ)a5�"��jc��`e�1E0�0�t,�[��i�ߴj�X�N�q?��FU�߻��],����rs4��� <�`hQq`����2���8�-j���[�AaI�f��	j��i��(<x����iR������~DLgjq)ޓ�e��G4�;ţ�/k���d��U�:�[C��t-G���p�P��q��������\�ؔ��x2�~��=
����kO�������\9����ў�9q�T���<�E� (Qd�q׋�?�=�(�?��U�@�5��8�����~ 5-;e�k�(<���δ�!*�Y+�ݩɃPH�S�Ll��e{�?w1e��i��N�9����mn{��L㍧�����Y+�-u�p��L���e�[�e�(�g�������t��?4Ls�c�q9He(�����9ԗa�X�+�GulUM���85��|�3�}s��ay&θ�s����ʄ,�c����HX^ԃ��V�����%�����2'V�}w��:�J�G�D$��ݠ�W*-�tn���O\R+�\�Md��9�.]����� ؈�0=�麱_t*,_@7��Dm ��C�U�S�%cc�P�a��]��X�l�9�]D[˰5�P�D)��w�~I�B�?Ti,,B��e��RN�%?�5c8*�F�lfS,���Θ?5
PQ(�_$��H��d,�u[��	"x�򚣰�;;#AZt,��p���bH�d)<E֏������Jӡm��h���i�c�0�槵�
�Q�z��QNP,�U�1�<I@69:ϔGds�nЯF�L,��Ou+������K(xG�R���
g�!$�FM�f���>_��w�xq��$`3/���5Z�=�l�9��؀{�Iy��s�نc��k:
�b�����v�.���$I�b���5�r0�G�� �)�[��D7κ)�-��Э.��Q�c�:%s-��؍�'c(���/�.3E�i���HZן��,#a��i}�~`���N�[K��V߽�)�Jn��5[����0EL�n�dja^����9�OB�	�e���h���!����N��V�����8�1���V���O��g:)ܭ����Q�Zǭ��E5��{⼅����[M�h���c��^��7��ȑ"c�7<��č�{31����|= �����+TFX����-� ��ahK*��[q���ǹ��2�Z�"U�)T��9Z��63��^h;�.Bݘ��S���OݜU䪶���pc��9uw�g�{��R�f�i���2�R�h���]u�
L�z`U
ߘ�Q�p�6h/!e	�yE�k.Z� �Ǆ�ۻ,�QT���U;W����xB�mw�����Dg���� +H����y��	4,}�OE�>b��;;u%���~�o�)&Uر��X����/D����I�z�},|�w8AƤt��mG�C!�����N�^�Y�'�H]���z��zaݴ��'"i$/� x?�k���08�$��h���/>`��(T��F�S�\5f/+���A0Z%xE!�_�L-��cL""dH(���ڠ�~�����^^��8�����qg�{gmF�����6Bnc��s��u�������-k3]v��4�b�9z�}ᘛ|�O�=7\�=�B�Ւ��q�}�k�}f\c�휵\� ��gI�����KF?�'}N��Y���8��`�^5�T�$2�7��+g�V��ڳ���N=e��0����X+�I�CNyv�t��������$A�!Yp&R��"��8�xPu(�9�)t9�B�Do3���JA��$�G���nz6~Y��6X3 ܸ��r��������l�>�"���"����>��3f��}���~�@A[��!=�S��]���.~�0$̗�u6�*���mWg V�K���e4�\C�0�KE���N���w.mo���+���FEB�p�2טR�&��"c5��(��+�j�Nu�T���� ~.����I}?kD������/��=u*�\�8%��|��s"%'���9I3!�P��Q"s���8n�q~Z�^�/p��Ni����x����^i����X}�2E�+��|(Pn�DV@�;K_��kקc�~��g���c������X$,����K�ң%IqYn��N�:U�{�5�i��Ӄ�-�3���f7np��$(���ur.�V�c|[f�(A�3Jzj�	}���_�e����,oi�fL�ڲft���{:z'����7ހ1E������FMo�D�0v�_]W�z�M!Ië�-�lCf��6x+Ss[�_���ğ%#]�N�����+����a7,���ޘ��Aڸ�3n)�5��3}���|�;�_ˢ�G���]A��<rA�>Qp��$y������rx��>�����D~�%��]�J��#;x�uy s�� K��84H������ve��"�>�J.X�LlΊ�n�_~���H5ʄ�
x��AL�2�9i-[g³I��q���g���/�20��ǵ�oP�:�nV�aJ�	� r��nG78E)�Zb�	.�M�oD82�Ac[dt��a�"��lQ]Iw�� ٓV��ӧ���qQ������/
�޺�q+QJ#���뚯l�u�D��e�R2��*�CH�.~�w�+0�<�����^B]&�Ք��,���زp}������<�,�U�:n�T�@��[n��)�u��	KT�>#�~jA��F���&P@�}#���
���vaՁ2Ï2�_i;�T���[�q�o��kd�e������=6��D�$%��tv�|������?y����n��*��bΗ�bW`�^��Sղ�-�\*oj�prj;�"Jf����x���g�X݂�I��SӠMc���_����e�4E��@u�T� �n�����BkW�nP���ɦe a�S$���z����܊�F_�c.���~9*)��a(�Ѣ�J�r��� �<5s�2N_K���N9�\��Mr���w-1�$'���f,I�KC�q�Mb
�ea��tbyI�)\��<	�B<�����	O[��N������"��^:��D��"b��~N"e{���=&b�T��n2��]�X���%����Tx^�����mAs��J+±ͬ���Ԍ��AQE�[<b�͡�?�[mkLX�D��b"ۊ_�9�gL���3r*�4�Jz�5����7rK{xeG���M��
��*�<�\��-K&�Ž�M��/�[z���� g�*X�O����aU��r�(R; c�P�~���
�Ğl�M��O���� ?뽽��d9[�c���Y�_��TW�a��e�~:�1r����lE�4:��\�`��a������U�����8�?��v� �@������Lc�����5,#�G��oF
b��fN���o������t'-M#��soSX�M�2�O����=�=Ր�@X���T)�F�0^k�F�¢�tc�w[v�`}�!���67��������n�����-�c��e1R~�Sz�d����;|mێ!{�xq�w��wRH�-#]�����ʃ�7�-��_J(����k�d'\���N��R�ig���!DR�GW��h_�(`:�|s��"1���D�:�W�1�~X��Qh�ŦJV���fW�L�dx���3��e�$�Y�q��c��S[�{�0���xƚyI��<4r��h	�U����tB�����)�W!S�Q��wj���B��޷_U5������P8	�M_Cw`A��pd\=m+6������YH?�k����4��;*�����E�ЛQf2��9P�8�%��k�b��{"ͫ��	<�2�yŅ��-�9��H�⁨z�st?�H$/�S��*&�����@i��t��L��K�Wm
OǇ�$��4�|��
�J��t���q�O%�;.4�#kx�_�?P�d�"���*
�6	�m��|q���d�\"j�':�#���`���;N-��9�$T�Ć,CI���'g�_����M@u��O�%�P��$
!�[��sZ�;�#�đ�թ��IuMO�P�\ƙ1�"^��p8sn�eO���]��X��m�g�^P���~�n{�[M��<E�Si�q&6?ZX�lt~��q��>�KxV.�&�L&�.l V3��	� IȱG��1�Վ����4�P�{R����m���a�l�t�܊W(���5��uX}�\��˲�y�/�PmU8���F�!l ��o{��p��[g���	�JBra1�g^�G�`��|�x��9w�E��d4#����u "�㗚���х���=%�쫓��dE,�{�0e%�
�0��r�c[k�{�~G`Ь&�^
r`i�=��|��x���)qiK������ř ;���Kd���q�#�tN�n�"������C8�����<�1�W~���b46 Qd�?z$��2#�s�`r��9W�r�ʇ�!?Z�'6H�@��QJ���r��fV�/:�������3��y"��ᨓ��-:��\"��Ȉ�0�B�n�Ae�(��feD�A(��Ah�k�,��:��+�Ϊ���K��uy.�&�c �O��%nZc��^�V-��������	)���-��R���b�^2��$�: Vj��*`�=,g�����ˏ�d��L��<@��Ȗ�}��TO�Ҧ�f�L�	a��oK0�Ђ�P�](̓��V���鴢)R�| ~�v<�KrE��O�{��aV�.?O�L�Ld���Ev�� ۊR`��.�j��	oUixMG8��q�U�Or{4�`ԣ^t���0j�\�`(���9��lن�&�T��4�Fp��B^���6�R�"�Iz8�u�� S%*6a8��w��8���@�n�ͤ�����/������}�hf�`C�J:�LԳ(�R�]�Q��6݇136I1�eBQ[{�=-~}i�n����Q���EAL��ٓ׽���(�D��݊��g�)TѬ ���5�GO�S�w�iN��dDHޥ�9�J����f���+n�|8T�t���~&�s��9fU��������W�s�̕0��:'R.\����,�֢�q�g� ��j���Z�杺8� ���p�MŚ���P��&�F�E�$�i$GI��ذ��ylL�<;�_��{Qf	{=��F|�pF�Ǘb�#�)>��x /AW[�`o�sg��&����W?�u��[�tv��zB�2Evy�jDe"��K(m��DT�����p	��}ؓ<)�QY���̒��@��:��xPǄ�Q�5�ֈ��V~6Z˰d�@� �v��Uv� 6�r��k��W�?I 
1���Q�/-ƻ��{Y��
J��gsC���5��%ō�7�R-k�k"F�E٤�X/�f���/tk_o�]\���*�'wuC�:�:�+�U���	yW�*	&�%frPe�6��]G�0�1c�!0h��lD-1��J�����"λ��s�U��q��_�|4y�9�fd���k?M:��F�f����ewin6��W78<�9$�7�q�H�qWU��*�{U'ϊ6sF-��Y�
�HH�6?^��>HŜ�p�gL���崘=�͡�k<6#����" 5��^O����
�W��:���x�=�O��X��P0-����0z#�^�YZ��П@���-?-�BaTᛖ<{��UI<�3��:��M�¤��8�9�|��M�	Tqq��\��u���D�۵Q��1x�QLˑ�X*�����O~dj�ˆ.�\+�]��
ݎ
��̩�/8D1co�f�6�^�EX�MU��к�"�����TA��i��mbA'�m���̈́6
�H��:�g��{'�#�����墿Z�hةGR�-qOrH��|�2���'M�0N169��)�M����7x�?f˚�y�KE
��7I[)w��fU΁-���Ͼ �We6��h
mtQ�����tE��)��UB_�5H9egL���o6���`{>ٖ�d�}�Ű{ў�84f�v��	��v\�GL��#�]�J�"��;0���y��yr�p|�Z*�?��2F��u���m>��V�z�������C��N�݃�es!�:��1�����J�^�o����4^���]<�tջ�K����J��$�yl����3���6��� ����u|~[�%P���Ye.��]����?5��e��E������p4�Q#k���<�ik�T=�g�J��Wn�]���˨�\٭�5��0S����{us,R�{�s�uhlU3x���H�cs���(k?q3��J��I���56a���VA��
�2��p���up�̬r�P� ��el�y�~Sf�.������uɜ��!ЧV���j	�
���O��#97��M�`��g�U� �V���|4N���`j��Q������fB�1����¹�䆝��ܗ��^;:���T�YTm�V�SHړ��:�Ky*��v�f� t�y��}�8��G���˶��k��	��5N���Q�z��%�S�;h�zM^l��'��6���~�oa�,P��U�S�gd׆��cf����?�P��Q�h�;[c������F�����B7���~�-Kx�8+��v�y�8�����H��ַ[�>��}��{���f�?!��x�I�l�������.cj���0�_�v�L�)9����U�/���-7�.iB>�ym˃�p��V��0O��~@��P���[nD��Ds�`���CQ�q�'w1���kp��A���q��b�Y���<2wx~h��|�A�3u=M�9~O�9�]�9�A0͟�h��`Q�I�i|0d�@���vY5�Z!�>�a�?��Lq�!�M�.�`_���S�~�j$��z������.�8�1��0�Q〴�X�V�^�z������{�6G 8�($i�!%�^��$ 遺�iH������o��Y@��<�P�a�G�6�Ǿ0���$s�8��RD4>sA=�gwy(�w�E��W'�,���he`��_3�~��Ђe��'l�~o!����[O�t���[��� Dl�%�jR��JA�/G[�>�v��|oJ7�]�$�Bk�
���RS�B����Zn��	�߷\����xp�c�jX�g���aKl>�%x S_IH�ng���P��	���8�g��5�u�z���&o�}NQ�p��������B�����(���r�dW1Űg�>�C ��vx�MX�p7�E�����HS+M1J�1�D��Ų�PJ��"fҥzŘ0W�ٿ������~y�Aa�?A���!a����k���k�!*��3@�Qyy����u*(�.\�{����5�f`$G��-��gY"V��MSqC�jӒI�h�c�497��%�~�w.@?f:�j �k�c����ʶ���R�H���ܮ�睧�o�'��k�ƴ�4䒉��Y�:	�+;(���n)��D5TGό��.X,(��{/e���l�З�;��n[�W΀��P-���� �9�,O�X ��)���� ]�~M��6�?�cP����([r�W�WD�Y���k�h��a�'���x�pָ��h�0�0U�P;ŏ&4pc"�x�̀�
�C7����o �C��\J'1��mگ�C�X�"Q��ĭ�� �!��P�D����֏<>��m#^q�&�t����������ڑ/��+m �FҴ���Z���L���:H�T	§��5��W�^i��F��b��=mU���x�ı�P���'w�#}�;j\Û��*,���;��_�ݘX���8��˕���*u���X=F߃ĵ;G�pH~2��o�x�,V\E��|���f����*���r�R3����2�`��}�S�q8,d�ۭn�"|������r�P����`�WsAAŇ��gP~\�O�J���كg��$�ԙ^����_��z�&�1K�n*�[�^&O���G��}��pɻ�H	ҹ�6E'��X��4����Am����uv��:3P4I��ߜ+��W�L��#��Oʢ���,���$����ܓ�P7ҨO"dM�x�FhCP���.<t	CHў'4��_��w�Reu���Sg��)�
1��>��c�>�V{2N��-v*�m����}�G)y&�S�o��5+��?];�J�v������K�Y��:*6�x:ac���誸]%���Bjx���1�e�VҞ6|+��"G녴�Q/�c�:(%�	��Ι�������fӗyx ��Y�F
{)iܛ����r{�O��9�E�iݩ��!�D�(��a�&�=:���w�,[�֎RҨ��z�-�j�L�iη��
s���$=9�t�{Bb��AD$5asa�>�h�{���#`����tI]wG�^}�Z^A���º���t�S�\�=���ϲ�U���P�*0����d~��Z�)�a0��H�i%�S�����G_�Btz�5f^J�[?8�Ҋ]X٣R���������$`��%��ᴴ�� ��+�ǣ���yՏz��丈�$.�տ-�w��E�b!�mf"��Qƞh�lG)oKb�tw��E�����J����t#��G �����z���R��\�/���4zW'<�RR��akL��^{BÃb�ΑӾ<��*�M���W��厢����O[LX]�̭Ԓ�<pP��Ӆ:'���&���hœ:�_��E%x��a�����+�z0�����[y�txDkkv�T���n\j#i��M���|���kW��n7̤0Dy���ɨ��.(9D� �,ܮ�� �2}�VG`u*��s)�Μ�h�߈��9�Rk�+^�GT��j�R���v$�a���%+x���n�-�

�g�#����K7��*m�``�6Y&��@R���6ulX
�D�-��~�+���]bP� ��egς���.��}S�Ʒ|J\*�u�Iz�t�1/�+��)4�������o�J�]��eE��ٸ��U�m�oD=8�S�
5�Y��,����R�X��n��!��Y/�3@r�`�6�
x�whY�%�l�����L��/g��@��
@�x�%�8Y��p��=3oԗ��mꫝ졁����Q�eE��pM/-v ���Ì캄&�1�\���w�H����bK0�!2��o��$�1b��`�ޯ�	n���Y��9��"l=!��SB�ĭ� 'S�׫>¬y�Dd���}���N�� ��?�i6фܫO����7gd��ᨽ~��Ѓ�0|W���U��L��Z50��biwM�+�e�7Maw#E�B��DC�����w���Q(Nh4�d��*�\�k��
Z��Ԛ�QJ���Z� �,�@aC�Q9lc�@*\���ꂘW^�ê�/�}>��Y[���H��<�s��kE�3a^��Gkqw�2�!B
dj�Q �i�x�r+�Mcj���m���a=x�\�&�>$�`(�:) E-��De��zYئ\��]��l/���$J����w��Թ�RYZ�dp��� u�����}��Q'��&	ڿ�-/��EV�����XRi!*�5�����"��Y��@�3���4��g�zU�t�Ǔ���a1جb� !�!9� ����)n��?	�>��k[�����i�����|�4�=����D���h�n	ǂ\�oL^�Ux�p�'���	�Ǫ�e��Ti���Zy�����-�?ೀ�����M3�&3�kC&qa��4;1*0P-2��%����ӌ�>�OhA���؆�Q\L�ٱ��3���'��.=�e!��`|$�+M�ql�(H`ۀ�}i*�3l����p�k1Ody,�{V�Y%��K���RP�(=�xj�QAo&I�K�Θ����s+�3:�6�ۏin�4�!k���[5����Pբ�jt��&��� �7ʋ���P�+�����:�M�����w��9��|�.m�I��ybI��]�i�7����0�[�����C#�)8�m�@_�����m�;�U�3�8��g<22\	�V�X�Nh�h}�"�{-LŭaR��v�Ӛ����1�R�bJܑ<����K��K=���t�J�)TQ-�$Kя�����zCF���j��{10R�H�_����2ݠ��+��WE����8�\���ƚ�&l�j����k���,��Ht��1�1#��8w>�yY܂�2����Ƚ��k����oa��<eu_�5I�:1��h<qR�K|�;Q���6f(�Wآ��e�]tt�^l@�Ae��oP��&���o���>]z�����a]�Siԁ���F�d�����^Q�I��ЯK��tz[	%��7U�S��D4ϬGx�F��VN�@v(�r�	�"t����N��wy�a
�f�KlY����ŝw���x>c�@g�J�&L�^։�d�4���<y�l>	T~����a5u��QJڬ^
�$�.�"ͺq��~2�?2�ϓ�o�bS���,�J�����;Έ�v�n\�F[�-�i�%4!g�q�̵���D܅��V"|Ǥ��Jஙǰ�j��<W��.5\9���"��O��V�<0���{�pjEc-Oƫ��S�39:G��a�j��b]0]	Wa�)�lk'�Jڼ���Ŏ�B�%�隖��/��9�k�h��ѝ�ܴ��Eȝ,U�+��vS�S�=�(��39#	dX5ӟ3WK ��z��i�q����܍".���NfW�.��.m��c3���h'�꼒r.h�M�|��<W�(+��N�/�=�"�@��>Ҷ]��dP�c��U%J�<,���;Pэ�������I6a��<���K(��G1+�3`l�k�"_u0E��_3�0�n^X�Y#������u���G46��[`��)����w8E��28�d���D�Uo�þ�Z�s��xHUR8'�����d$�ĭ�L�fq��= ����sN��hmYzӣ6����;����+�]ce��H��zL�,�I;���:��z��:�'�,��`K<�R�����0�Z#�9���Bٚv;�&UL��ϓ��2S��>s��V.�6�?xWv!fY��6��Zd����}_^���/��1��\H��Y�#���;T]?��WA�'���̩�e��7��FS�ͺV�*;�a���9Uj ���'( XP
�ڇ�C�"��N-������gRz)�=nt������lǹ�쥱ߙ���vX����AE��!��*_�K�f���cM'a������\��X��:�d��q�D��#�Ǌϛ7��U�`?�s�M/�0��fs�5۷��Dp��k�m�A��0�+�m �4YuJ��N*dW���fL����G�~#:ޡ\48vzߡ]0��q}��Dj4��l��M|���I�*�H�bW%���U���e��d�DC����^9��]�k2�
2��>�MF)]�^МOa�,��|�2O���ׅ$����@�n����|ݨ���ݦU�XT��F�.���ג�ϳ�X��Gu0<�:I�qML��[8.$à�9a���&h���_w	fžMw�eT�t�eRm�q�W���=���	9�xtW�?'TM��4�d!7�h �ud�+��7IK�yF��'4�%���4�\<P}�g��M����r6\J��A��`v{P�_�_@�I���̛T�6����ܑ�j� ^��AC)VkL@&�� {JX�ݦM3aŇ}�-��d+n�hC6E�V���S�RW�ގ���.GI� �I�w��B�6��#~�v0����)�#�1��n���a"�>�9�.��J�Ykr�*�rp�T�_����5�}#�[˫ى�e��o��(����������ݚ������l�ƎXN ���|�f���`H$l���%j!:���9G=յ�?�a0��٣���}�M60�z�:�\���wK���-�-�$K[�3���y�{�������?�Ǯ�(1b�x�d�s)��D��sJ�e��7N�p��r|�\Xǂ���"ίGa}O�g�����b�"J�蟉h<9�|�`p�n�����I_/c��yu��*A�����_��/�q��ӊ6�?�M��Mfռ�[��%N�@�9���m([���J������������(NR.^��I��E�H�MOy.����\;��jҿ �&����b�g������I�Er�µ&���s�$���q�������d�����2�ΰ��1u�@�L��َ8�繍P7`�K�?���& �����@�\�U��+�jrʹ3����Q�|���ϦD���d��hR �&��h�Ъn=fk��2h� ��t���%3{RiQ���y��������nt�s�f�h�3�E��ɸ,�Yc9Q��������v��<r�:�X����쟦��0*�Q�8��$*�x���˸����YA�D�ld
��֘�:��.��x�<{e��;j�f#/6�ӻuUC�t�Ժ��E�xp>�g<������׺�c���^�*C2 �,˔A�\��
�ΐz~bԬ���
'.�r�>.'eؾA�`	rو��M!����OO����f�bQ���tH���l#����{x �� Ll8�����T>�����@Kl�%�a�
'�B)������
�q�?�-��ޚ�B	\n�|�[vcUK����f��3�W5L��]�<�m�� م���^XWa��A�#��wX���KC�I�.&d]�``�{u>��O"�[!W���4�q�M�j�����!E�O�R����<�%�m�k�B�E���=�D�) ��\PTycT,��(غ�!٥�w��C+������o�^.O���tad��n�^X��S���JN�oۢ�u�qh�S�jIU�g���R�� ������a$%�=n`��[S�P��4*�7���DcA	����o��A���δx/ǹ�|+�����+��A!�I�:��~�j�W�k�S��HsMU�f��+%/aq`�e�����q9�!�����|Ja�}�ѕt@Z�+�ѼI\-
��RH�W�W���rҴ��~�j�N�q��'*RY�y��E)�"�*��U-�*��q����:o�w`���H���ӑ�%�.1f6T���G�'E���_�40�>�g�'WO��҇CL��x��3m.��0��!TQqY���X>�E,0���V�-0NX?T���|G��l�Z�c�>�����2�A&?�Q��	�����Y����38���>��idY�XP�գ�ҁS篊�u��7�n�PU@oQM�z ɤ㦰��Y˞��s|���"k���_� ׯ%[���rc��ol�Y�/mY����T\��O���50w��3�}(�ҥo�nj5�z�K��Č���["�C�u�D93ց>j���[�`�k�rgB�<�o�&"�����Yf�D�N��@��Fo����+N�V�����F�B\�
���U�j�d.�_gW�������_�i��5Sӈ\K��r�6�"c`M]�����\v�|d95eX��˔@
uNZO7�m_����h���=%���-+h��k��ʕĬ�����^��w5Ҟ����7Pk����U�k���G�wFG�`(Y_ҁƯF���u�"t+bh1h�Ǯ�і�D�Q�=�\��"M5�uSŬ��D�?���M��K�U�HP�"	?���3��H�"��*��#������=G%��!%r�G>F�	���1��/�.����z�N�l0�7͜ɵʵ��h�Gq�o`�Q�~��j:�u��{x���_���n�^�Jp����4M�O/R���i��(�d�x0eN<�U����i�%z,Ҭ0F��F�jM�e�O��l��i@�D*Z����r�;9 �\!��'�D��p��Eک�y�4l��t��Ds���ӛ�����'�tD��
N�A�F@f���P��׊�!��W޳rht ��������@X�ހ
q��P+-�+���w\K�8����ɫ
)��!T�=�D�ĕT"~��U2_�x4Zh"	�Q�,aQ�R�H���cg��>�gۋ�0�@0�ɇ�����Lp;1�0;iX�l��ՇA¥|R�]���Ɔv����J ;S�2��i))�063�l�e�>������uI��1΅( ���V��W� � T{��|��O"���_
����LAS7�#t�4�_�����wnLr��l9�,V�2�&�/�=R9]�����نTm1'�ki25��o�Y�^dQ�E9dI?�]��헀j�b[����>b5:�?�gO��[=��A%,"�������_o�
U���X����n�F�?��dt8�ʒ��a0b�kG�S�}��ۚ�o���A&2�_���K�*#W�Y�8��p]�c�?�Ҷ�g ���3�:}!�������be&D��9C �ca7uu����E���|4���Kx�Vb�-˔�&�%�4ǣXP���8U!!����'y��ϗ#f�Tr&.��/�R�T:��׼�ɡr�6�e�1�s����{J龓P����SѼ 0�0_�1��Zb<���#i�L��_�>,Xƭ�ζ0��LbxS�N孵���dH�&��/�<�f�(I�s}���5��
�lU��l ��θ�ϒ�੺!N�8�U���� �:���g�S6l�#��c��l�˸u���)�|� B�I�@aU�ہQ؉XLx�?ɋli�y�!:	�0]�vW^#Tq*�]ę�8�"�n�
.)�[�~�v_�N���-6h��[�r߃}���XҌfV������W�2__����}��v��+�[�.s��JY�^�/Ʊ :]دy-i%z��do�F�{gͱ�9���G24ib�*2h9�?-D���@o,ˋe��� �+��V�@Ζ�r~�����jRI�I��@<��,�"�0i�>�@]4�-��ͧ���0��h��&ԁ��[L*�u�
�9�wK��u�TG�=���@��"�`U��֒UvC��9�x���v��r�d����r5[P�&Լ�o�(7L������;���� m�;�ysYT���g��j<��a+2[+���1��0�9��ί�*�+�@�6Yr8�Z� �	�UW�V
�ԑ������0Li2�]��M|4�:�n&�-�O`c�-���D�x���ŗ�3�
Y��Z:�a�5�l���e�C,?�������4�/Qw�|��;��n��2�u��Cl���m*Z�1�i�c:gk���ywem%LY��SO� �w\��;]�ys�^׸�!�ip �K�9��Dp�r`Eb+�>�+_���f���_x1�b�{J���&�$��>-�E{"nZ���O����r(�J��ѯ�51�fҐ���9�Áq��*4C�( ?�� "����j���@���tg��G_s,�%0.m�3����$x���q��,���	
�? g�l�=�>R����r�0^X�4��@���`���l��^>;��/'�b�ɠ�I��6\�TC���%��.�uH0�J��#�9�K����j��y1d�Խ��O;��5s˖�:�b��zA��1�H�PGwA�c0L�k
���Dz�{�e�X���E�&/
7m2�2C[ )F���ꊉ<�z;���8\�A�tN	�o��1�����P��Mv�bmELj:UȤ�Y�u@�`!3x���u���r�ty�Ċ��������1?~�>�Bh��l�y�0�t�f�����jm�"��Ra� ��間���L��h���"]���Ff?�'��<�'=4��mZ���CΌ8��}B{(JF6��e�Ju8o�|1���('�f�0� �`T�7�Y��¸b�w`�J���E��	>��_�>�d�V���d�h�xMI��|D�~e;�E�AI�6�|�<`_����0� Q���$�UĀ1���ْd��{�km}myyZ�޵f��0Vc�B>�ձ�����?ҍ��s�� �2(�xi,��W�I�>���s��>��Ĵ;n0�އ�z�l�|���`צ��'��?�~�D�Z\��qdv�����A��<9uC�� jI\C/6[+`�_$�
�%c����͇V�:p3��H��4���G�,G�~>��Q�J渰SI�M��T#'��C���}{�2�M/.��:��v��9�
_��%�
%�s���5dU�B����e�KB.��Ey�ULjE�:�(%�q��V��=t-�n8Su�p�_�q�R�y�Z� ���m,��kԷ9��a�1�����S.i��{���U��O~u��F1j�2�@+��{z�[*O���z��Zع42�+�g(5���,`˾�h 7Ft�d���愽�Z���],�!����a<_�f��5��^=1��M�"�1��1�z�lJv�; )�%/<�T�_�;xC�+&b��|!��uIF~�P�t��&:Ѫ4��p:ߦ;zx���38�l#��\C�f^@�]nGg�X;i�A$�<<��ZKts1���a�����w���1Xu���]R@��������4Q{K��!tD/ܰBݴ�a�R�\s�\r�pr�٘��7�Y� ��*E��^͂`V�`�0��gq�����+����X%���f����=X���3��/�=���[[�Y��`2��z|��q�F�o?#ݝS��;��9��ͯ�Ş?�"N�+?;D�(\�=h�>��HZ�=�\��6�a�+��PXA��Қ࿕��Bs��U�j��2�E�L���-�(m�x_����{j+�Մ��rP�r؏-]��*�ˑh�1n�_$nH�]���fO9��*&V�K��D�Q�ս�L�� ��FB�<�?�aW�P����P��UA'��t$E�R��H����4�����'^�iV>9�ɯ;�X (��j�d����lZxX��oI�D�JO.�]��X5��(�@���`�������>+���Qo��Ip����
0߻� Z��	��9:f�b��&@:�,%��1mEyi�`8C��(3��Hv��p��d�� ���a�w!��Ã��w�'3 4��*a`�]mj/�Li�d{�|� 
�s�٬V-!K��
`�$:�j�5��8�\~-l�V���`��靱 ���5�X-�2+������PÛX<~�xU�ٽں�;=j(��UN��ŏ8��]��&s���mgi8l�GW=P0v|�E@�=�d�IīÄE�j!@Sh�(o���J�;�]�� ���
��X�����j���G�3����<�Z44�+D�k�O���S3�I$x�����%7z7�2`QX����;�o��5����+^����9�-$H��^�j}n�,�Ҹo�ޔ#�0����� 4�@N�Ҳ���CS*-}E���"h��`"���L�}g�\�<V)��g�7�褣�[�|q�y�{���o0�2�ﭣ
>��vz�٥/��\��*$���J���gѦ$�e�OGYV�N�(Io!�J��G�m=K���
�L`O��#�X�
IE1b�1!��0�`����V�P�)�޻� �+�ɦ�����N͞�p'�$��9D��@-�d2-�F���Zٕ��q���pG�!Uɜ`��K�UC�ɲ��]E�]��˜�?�q��!3��!aD��ςZĜ��u�������7�����bg�Ê�a{՗-��4�(i�$aOrX�L���Q�_���y��ж�����'���{ʫ~r~:o�.��z��b������0�Yvp(��gQP��"6y�$�}d^V�#(��m��7�a�pF3�(R@����Y���J�+J�7ȫ�֠����~���Ј��a��Xh��C�!}�f��[<�x�cÀ�@l=d��SS���t�������!.���)N�Dʣ���LH��!#/Mv��ՠ��k@�3&����p�""0��aS��FR�a��?} (dK�{����C<nG(��28��C��S��5�l�c���c^�ͩP�y�����>2dC#7��7� ���k7B{��&��o��f���ˋ	F}o���9�r �#�0��QR޴��cN� ��@>O-����gv��wn6��VC^��y*��G�2N��ӺP������d�Kf��Km����%pu�b�맖��o�lm���r�_�

m	�R(c(�T���ʝ0d3-$�U^�R�X?i&�;�Z=O7��w86L5 <���K=)b���х���6�碗)�i�ުs�g��1�/��*3܂�������0���DuK?W<����վ�#�W�ڷX�9aev����E����:���ʂ�~з�"���ůu�j�Z/D� ����3{�	K(n��NIn^�q��<�ECF�����9W${�]��)��ڔwb�Fյš���H���%�6�Ư�D���LU�U�D�\H�69g���d�|`���}�T����)9E�5,0�H�-����؁�'q�d��)�ٔ)Iĉ��V5RhD�F5F�_C��~�PY�L/�����`3x��i+����@��M���k�h\�k��O8u�q~�ZCH��r���6'8������`�n_��C���ݦ�3���+8%�����dh�͉��B�}1�1�	�> H���J0�C3���H�K\�e}��j��衝eNu+m7'縓8����(M������NƯn,6Q^Ek簞?�!'I����2�_�z�Z�!�w$#rAs�"�*@��~ZKW[��P��	P��!��A [���p �j�(i���o��z0Vb �.s�b�gf�w��LuFw���UeX������|`����c��,V>��ʝ�/�&�	��Of���v�T(W����G_l�Lx����a*n^��U*rtz��G����k5���h�?�B;�� lS x	jR#��R%���w�8�a�9惗4�SHp�c�}��׾J�Ϟ�W�K�O��ݧ��8���%qN�-?l�D�/�S�--�I;�1>����CM�v�p�B3Y6��)��(+�}��}z��mr>a{W���?�t�ދ7�m@&��<a�=��a>/�(��l;���ݦY�%�)�F�<�b5�h,S~��-@���ׄA�
*�X�������b��$3��w/�5�аU�?�<캼Yl\z��YQ�h�i�7���af+�������}���/�:Sdm:vms6THK����+���[��7�>��ʲ��ۼfb��:/8�ז�ҁ�F�H��@烂6��c�x�O ����d/][M���)�1�%��ZU�t/�	!V�|Ҙ˦	G�O���[I,.�i�/A���$z���^�r�E�-��U�}�������Y<eV7��-=O��΄������{�}�c�>������&Qp�m@�5��Ѯ7_�ɚ�p��^S���p��H�c�;p��[�M ����|�J=@������Q�b�l�l�~V�[J�M�����"n�-В�5&���C�ڽ#u'��׳�#�r�C�qx�8�P�p��	O#m��7d6�w��vM@1lG+����3ٜ��p�[�Gr8�
*3��38����l��D��kO��/�d/$���].΍�V� ����KG�ه� �#Yv~��#ΨK�+�)f� 峅!;��hjq1B�p	g&_:��R�o�N�:�:Lb#>�NX%C������ĥ��j����[�v9
�!�΄� K��g�/�������D=%�����h����7$�j��h��7%��;�7������'�qj�⧜2?5>��ǫ��۫%�y8{|n���ݩ���5��Ԅ[F!�Ź��'=I{`����c����{"����V?�B��Ť��?�D�t���P_�q�(��Q�ߨ5�2ȏ�-��y�5�@�rD�	S4�뾪�����E���ivQ������
Q�~�Q�lB8V���ʹV��~AuZ��l�R�������݋@0��~�Ȯ#�s���]W�bE�ϵ�Q�n}gv�L�X<���T�Uc�Z��q�2��fv�6!6D�˿!)*i�g_�LY麭��λ����+(�k�����M�\c<.�v҉����4E�siU?�2�m�M�1���AZ������c�B�k�)c\�O�,� BPA� ꌕ;��֚��J>�3�D��yE�Zpyؒ����`��X�Xf�/� Fu��{�r
����� �[+��λr%'5Ik�;���m&O����'=�e�4�g�sW��U��tijvz�(��µ�n���4-+����z��Ȋ����.	��'z�[t��q��Q�~� �$�ѠЂ����]VL��:7w�r�q�}cB�&�\��݌�%����魝 �u:?ŋ�/����4����>/������k�D����C��b��Waa/X�$ջ�h	�
`���G�ŀ�u�QǏ֥L�ma�҄�%�}\��Ѿ�Gۨh'=������jm7:u]U�XR����4�U"X�`WEc�R��,0",8~�osفp�	��\�	�h��Q��;�Vw�F�� ��򢓺�Db[d���I/N��xA��z��L��Y7�`�}�u��I���צ��1W�*�E�ە6�/kt.���p`S�WhÓ�k��z�ʓ��=c�IGS�����=�m3��W�1Z��e�_q־n�4��O�`S������b���5�$f��E4�M~l�.��pϠ{�y�����[U��բ�E�䀗D"C�m��%B���PJ=���,{VML�����Nӈ^I
��)�g�}�Q��7�+��*/c&�%�UP͵�e�K����X�k�. ?�쟒�s}�0�I@�1~ET!����g����W:��;)�S�	�~�c-`��M��$$�)�0O�qT՚�pҠv��vLe����'�;����fӚ�:�J�&�Q�tl8J3����y�q&����n�����feM���]��\s��;9MP9U-�^7��!~_<;!�f���9y�C� v�s�z��P�Vy%΁`���Is��EAr0��A�"��V9k��{�����h/<݄�_.�mZ�gg!�}#��p���$��,�m}:!�L�Û��T-�B���2)9qC�Z���3GR�FJ���B9N�Q^�W5.^�FD����J���Ȼ�;�(�RT�3yrp��Z}y�˩�%;� ��
��^	��ssus)5�RrA�\�sI�fj�ŷ�����U�I�m�~_k4pH�		z�@Ҧ.(H�b�6�=b���7�364��2+(�ָ���G5~�q�/-�\c1�4V}V�A�(����X�c9���^@G֣M���`kK$W�g��ئ�_�R��ﯣ�d""0��ⷎ��Q��;��0?���h�d'�3����"vg�+���n"�L�K�����MN�CS�NZ:	��7�%����pP�ӊl}1�5;��D��|~,4�ap�ԫ��VLp��M�Ac�D2�՗o4��⠧����e�+7��؊�_8F��jc'�7��+J�W�����3�
Ft�` "pMs�m �k��/-�CEmX4����:Q�>��/�N�TW�B}oI��S��(��BʠqxŇN�ؗ�����$��nhy.���'�z�
�0Q���[�q�uw�TgS� �/�qQ�q��K��K��XC2��r�o>�9�+��-���%~������b��^�C��m���$D����{�CZrJA�%��}ɼ玼��
��!b�իVSW��`�@��AT�%]���:[G�(���ަ���;�U	QV�T��!	�x��-9�3&:l ^�=�p�V<mJ��[��x�^��^a��5�XŸ �=�ꅨ�[C�O`h��$%a(ĉ�p-��P��*��w��쀔#�; ��%7�a��}�-�)Zo��-Z5x��<�m.�hM�p�/Y��%�ʡ=]?�:t�+�)�ϡ�Җ1]��v,�������!�Q^��+���[��cq�,�F���t�6~�кWX��)D��~������14�a쭕;�SC,T����R��"y��[����Yf�U����	�Z "0"�P�S���Q
n�@����<�a$MAa>�J_���,�y@��(�~r��nz����ѥE cswu���M�FHJ��k|��rSZ�fo��C[��"A�B%8Km��4S�(�,�����
�����3#���>�s��4�{��e.CB��	S�	x���"g@>����}X��r�s�Qiv	A�& �$Ѓ�*��eR�V��#�9h5��G�1��Y@o��_�kBR1�%*�ݧ(�F�i�W����>h��#$�<��ne��W�Ϣ+���+��>���ti���V�1�Y��$�1�K##���.��ҿ�#�5"W��s�W�{O� v������W�4��R�b��O=�@涀��.:  �,�V�L�_�r󒱨����� $I/?�/���m����G{��%�qD�1�=�J���$�����Ӟ� �0 ��eX�,�F������@u_�/��k�J�ty!Hw�L۠�:aTju�u�#���"A�'?4zΙK
��@�`�h0C˂B�*��n4�,%x�MN�F[�ei;&�N�ر� (S��8^�y�������w�ȑq�z�̤��}~z�q$s<��[�8�2{S
vJzER^�J���l� ���A�C6�h-�e.p�M��[��ήp$�&x#*x�B�#�5d��	���BF�s"E��UG�����{�Ō����Q#��%�!P���Y���/s��Hz[�
�ovl�F��{F�+p~�R0�J�d��鄹k��X@�B�q�`$���C�}m%�(�����q˫�P��xS�!�?�co��*y�������Q�w�x��IU�=<�?�(�ݾ�9;����LO��q��k7�i{2�����@_���@�&�ذ���"_f'%�� ��&{��8jୋ�4߻��n3�9�E%�}�{���ӄ/�m�����'=�����>���_"�B��U�o���G�\�O0�>�!\��9�]%�1��T�;�i���C�J�qS9�Tj�}/~�!�</���"��M��]��J�cڅ�ؑ�\���Z��VqMr���1�ŗ{Ȩ�\S��p�ڋB��(��N��'ia��{�X������6��Is�#��9`jkzۧdU��eV"�z��Ƅ
؜����k+������z�y��N��A���D�1\�Λ(֎`se��S��z �,�r�F�Ǡ�Y�c;�	/X�G� $d��N�X{���
bNg�)d'��!���V�؜�U8�rkk�W�>x�0��A��\n���G�H׉"6��Jf�>Ɛ�s��~Q���<������RNXԭ�'�m�d��R�������{���s�_b�T%��Ch�M���K�%K�TE�=�'J��Q��\f0��*�v��%b׭��_���v��Vphzsl�Co��T��� �4�JP�-�2�`/�G�up+�gd��_{I�%�� $�S/836(�����q-��O�%�ϱja������aa: �5��bKf����{e(bG�p�`����l$�!p�d=l�0�
2���a��A�^�����I���z�ٚ���k�q+��v�Z���H�y_"�'�#-f7.�w,��6q�n1SL/�xp��8�߫�z�䥃0fۊ�c��
.`��Υ���!빊�0�_���>ܶR�0�n���E�g�;�8��8���J��|*�aS�M*���ލz���H9�!����l�w;�χp��S���o�J1��vˀ��	#S[��p��+O�h����p- v��6�-��ϴ+��ͭk6z�F��1��E��B�3�b<=}"�`B��8��9�s�?��W��;H���>%x�Ϥ]u��\�8hm`��&�37�Ǩ�]�����Y^��8�1,$(:��uq����|ɍ���>��=�"zʓ?w�����w��R�yp��:��"Q2|�B;ͬzJ����G�¼)b��+���ܯ~1��,�C!8k���6�}�u��H��O+��UGA���%#��A���-̦�'s�e�[M<d��*�Jq���&jX���Mܩ;��p�])�B��E~/XÞ�h��l]xA�?���ð�Xd����"��LYM�9 �*<5�ЂX��'nN�}�9vtm�O8����빌*�}�I�K0a+A�LP\�}n��d�x��+ʓ�λSb`����7��c���Ǽ�'m�� �ȗJ�5�=�)�ޅ�u���i=iy��6@>�Qh�(H�ޟHhe3:�=h)^���؇<�9�CE�-,:� ��טƲ�&��	��%�/���N�M�F���_�J2��q�|�%]C��yW����
�Ho��Qծhf�B�`3�K�l�5�[⣟�!SL��u/�OUM|����r�a���aS���~T	�,1���a��~���q*�����"����V�ng��Rץ��}�K@o�)KЀl�HP�_W%Q��0�}r#f��}/�H|k���`;	ɼ��a���8a&2�o[�iC�Udc!�W2�XW�E�E�b�G|I-� j\Ul��0�z}(�4��K��@c����Np`,�`��;
!�1�#���G�]�	���s3�oӁƥ �5�R��&��~e�M���:�K;p΂�O�ڐ	��E�$�X��t��Bv=�	�X�
���x��cײ��R�Y2�1@�)��?�J���S�Y��� 6L�B
�1�?,0��p�cGv(ִ o���0�ᾟ�i
����3m��8���@�쫎AU`�Oq	Oa�u#�r*1t���b��[?�[�Z��E�} ��)^ը�/�V�xh��Y�^�����0�2[��^�Y9+�!��n�sTG�U��Rg��a�^���Zm�n�m%B�3�@�Wp9싑��4:E�/�G�R+R_uS����$&[9�vx6*`eu>�l�N�?��]����>�-��@d���E���/��Z�j��
;(��)L�c�I��n�!l���v��Uʂ*.���W�X����[ȥ&Z�則�$���t���ے1x��D]S}���$�q����gw�B�:�k�W�x�3t�cڋ%� �ܴ����
D��������0�;�<�3�I�I�Hj������o����Z�OM4�������K�C���s�;�iRTV��>��Yڳ�w��H-����(N)�ۚ��	9kv"�ڕ'�{Fsڒ�c_�R#�tz�u̜��+�@�9�q��i�UE�s"� ��M*��8�hse}ߤ�E�k�]E$7��櫆�a~�Vs[�[�`۴D5a͕ze68�@c�;bƻ���Cu��FWtN�N,L����̜�Q�T-�ic�Iz�gD�K�O�J5y�IO`���+9�OJ��݃���R��uKf�8B�~��� : �ޙ�4��m�M�X�M��	)��Z^H�-R�0�5��r{2�\&��6�H0]2DFR��@�bP�]�AԲ�� GU�~�%������s����k'����јq�� �v��WĖ3�81S�֔��Rғg�:�\S�cZw�D��E��^�v�F�|]�����F��y��������ēZt�	��"09��*��z�ܖFr��ֵ�Jų���O����UQ��u��}Ny��V�\CP<˴x2'x���j�GV
4�iss{�����{�=B����V�օ(^U]�&�-�g[$"�B/����R޲��0�5^R�\^&Q�[��'?r`�� b8xa�:�/�g&��%��:���K1��*�78��
���n,}���t�y��4D|lo��3�4$��p+����W��c�*�*֑Uv�>̇
������D�ͩ�؍o�J�ɥ�E�y잍���j����Sf�؉�J7��<aK
D��tM8̫���������l���X�Lj��l�Ή43b�p���ك��>�(r����r�:�ǈ� 13'��T��	}m���Q�mR���H<��I��|�w#�2Z>%�,�)�;�~)��]teKN�g��-ϙ�o�	q1�FCJ�pzU`zw�8�b8
�4�4XiOˢ��qv�`}Q���1i�l�U4��zZA��;.�M8'�@z��]��fA�F"R��H|t;s�s"w1Y�X���l�Rԟ�&��;���!�r����B�<����BlQ��#�'����*D�֟���'��:����+�,�,��G��,��'�A8�s��4ٞa��+�SG8��!�-�P/�W��9l��T����,~v�T�V�֋T"�d���ޕEK���_��t������-�S}��.�!�W��,�� F�$q�q=�ˡ�w��%}���
S���K�%rjxwZ!�i�@6�D�Q�0:�(�;�ZP���[>�-��i\�_F���D[��]eo�b���8
`�h�<5����4�����0�l(�do�x���&Oq��]���rcU�#�z�����CZ�����
Om5�h�#�*�Z��CP>wj��I�bM��i���(J~t_s�<ҧ��76����L ��Y�Ա�ջ�.c`Z��|,
#�=Q/u�0�����qd�'OO���� E�3�Y�\?���4
&�(��7 ǁ-�s��z]�ln�$�S}���k�$�x;q�v,l��?&�ם:bO�w&Q*s'����_����2o�9�U�V�e��9(�}2G�=S܄G���UM����+���,g!�ZF�""H`$N��Ƀj]~�]��������r��W��Pc�4α,�G;�ts)+u���������.���[��u%(�G����1��#�c�H.XC���:'���e8#9%��F
�]3"��654k������|ʽ���dtdx����L:j�a��WF�M	�.�Uyػzʛ {�=� v��RI����y�q�unY���tUIL�ۦ%�0C:*o-�g� �=��_�׸�6��.�ɯ�:ک>ÿ�?+] �4\�q����r�̜"�VYg+.T�����4��"��X�C5��QQ؈Q���A���7�'���۩/�Ca�.V!��%˸2;+�E/Z��u���JC확A��}=%�G��s�~F�H���>t����I�G	�Å��[�FY&�&�����D��3o��1׀S���- ��ѱu��R�&G�IZ��풓�ҷ (�Q's|u�cv��x���l;��2��ԝ;B#�1�N��߳���fa�/��Mt�"J)e!
e{m,�}F�|le0{SuZ=�G��06����O69�iS�I����W՘�·?��T#��I���7���:�ɍ�*vÏH��a$���6�G��,�@�1.�Ԏ�5=��fH��X�����u|f��܂bӹQ}���
�jI.O�����!��XuA|�C���$i�IS��J�(mWٶDM���o�}�[�:�66���U�[t�p0�e�GN��Py����602Eo�� �v���N.��J�r4������>��uE#�8�g.� ���n	���y��Z��?'��tm.�015�2�{�;�1�5$����U�>�i��C�a(�"�ϯ�4��ԟ/��C} 
��j��2�����lq,c�]?�GI�Ǆ�ҝ��������~>#��~� ;�=����IxN6�{�9U�\$�pf�F�|�hE�'aޔFK4���
���^6�O�x�+�� �.�bU§���CI�v������>]nz�#g��M�Лm z38����J���-�%��O
z��kd�!���y���B�陇�ғ�Ft�f�Pcn�%�mIN=KNiL���e)�������r����ܹ�0�2�M�"{��ڳf%��L-���)���ks3,�|A �z�|�9�Q�V,���w�tѩ�mR���O��%UAI��60�d�l�b!���ƳV��{��.q��`����+�tf���RI.�b�4e��1հxצ��&n'Ք�:����_���6��I���4c|K���e�{M��mċ�1��ى'����PU�R.܌����-�=P[����E��j�ҺNK�rc�:��ײl��i@�T��.b�!�K��z���b��I#�S��($�+��!���a{}�;Y��EV�W��$51ؽC��!���:.,�Y���X�h/Rl�E:��L���KcB�k�	�1�-��)�p��@B=���3$sS����k,L�pӺ{~�Qx���f�W_�y��{�ʰu�D��Lb�P}�:�B��eZ���V\���n�^��#��8�-�!�A�!~�k ��-ˎ� �W$I�Of��c�ŝ�K ������1��c��A?Q�,VCZ��@��a��)��g��b�	��A���E��vκ��tc�zcK�d>v�sZ���R|0��Wym^�2|��c6
+�H\p�+�U��vie�,J�����e#.|��F�hA;`B�^��Y�?S����M��05�Ƿ._�|�z��i�c�	�t0w��>W#"�l�0�]��id��t������97��<0�m6@>�a�V�k�"}Fʰ��%��rF-�G�M ]m�i6�4S�+���u6�3T�X�������{�k�_�ݚ��V��b쨐=��ߛ�6���cH�~��D׵�_�[��d?C[�jg	�Y�t?�pxib�zQN�n��:2m�f�z���D��6�O��j��mlh���>#�[ꑾ ���ٹ�����E��Tc��XK����xM��PQ�E���ԭ7Kwp=���XX'V	c������-��zI����Ϧ����~J��`���H����_L���|k�FV=v�K�|Bi���쑤}��X�m��8}(�y��T������/â��#������qúl�����z�4v-k?�ΟԠ��}Y�*mtHEx���e�1t��Mg��>-;Z��O���
�]�e4�T�`��v�#���Mv����AC�|������Y��"AG��a�;���!�80�h�qҵ����-K���2�����,B��!��8�j�e�����6��ڥ�\���7��֍�N��E��z��x� ��fY/>)���nft����^fl���� ����@N��İ�6�ȉ��
��EP�QN��lEvq�^�]�j��l��*�㑫c$��ə,�C��Bw�r�f�Au����W�����G��Mv���"�Z\� ^l����/<���.A�8p�;*f>�=�)�Q[�0�q+�J�!��=�C�͸ѿ���&�|��?��]'5�'O���hR��H�x�i���7>q�����X�R���t�7^6�Y��^��~̆�-qu<�����F$�T�k�9����pR B&�uϺ�Z7������p9�F	�D�&�ٙ�(����X������JXp1�(��p�cciS~f�f��v
�������C���R�A��Ξ/W����sZ&��#�}`�08ʃ�	�B�zO�� �ߴ����r��	l��-���p���
9��� IDZ8�fi�h��uqd��/�m�]d� s�f�U��vH�,�<����z�y	ԫ���! �aW[v�`��|/T�����r�,��P�Q��Q��r'n�eQ����Tޥ~:d��wp��%��jLB�\ �|����秊h��jj�3d�����]��,4xK����7�l��m���,6��U��{�C�g��&��)t�/���s���X��A�B����S�x��T�x�mE�F�S�G+��S�# ��u0G�#FO�� p�4�t���n��Z]�2�t��B���+��@���'#ri��R�,��+:f�
^t�r�i�o�q[W���6?�f���좞�N$�h�����;�G�����J��@�0�_Pl9�޷��;�^�	3vι1��-Fo$�Q�^��(�?r	<E�À����3��vI�Y}��e�����4��+�TS�i�~%��%�90�]v$l,�Ad�K�����ɬ�꜕�si��M����� Z���{�������|�m� .)"�C;�����'y�����^�x��b*��o������Jfd���`3�m�ȭ���o]�	[�+��{��H���+���,�`�yHy��َ�	��Y@����a��,$r5��=��7/A�iX\'���&��>�#����/J�8Ԏ��P.����l*�?��P����cHhj*ӗq�A$Z��Q$H`J-�<-9˙�F��JY����W_\����m@��t�WW���z��Ķ�-��|��Ϲ	�U�����{J�=�/��=a���[�y�(��c3�P�k9��rw�4�����j���q�I^[cW���X�����C8� ��#p�F&*'ej]x0����D�U�4%���7"��5 ~y�9)u� �.�"���[R�|��3wW����׽�m��Y4������⒉��e�*�d�=�,�Z�+H�~����`�.�ٞ.�R������Qd��L�Z��쒟mXyό#�9���\yb������P�{t�$�6�%�#(Q�����%�򿼻�As�L7��#J]�!H�������s�5S"<�&7���u�(���η���;�Ŏt��f�i�����Wᥖ�G�[ }&7�p���o�.Mb:��g�e��.c����L�~�R~�&e�y�gghl����]J�!|΂����V��M�* b�*�y�KA�h��ݴ��������:�|���t��Zk9�2+3���H9�VA����]��П���[�]�$��VN�&K��F+��x�<��q'�w�����Q;����i>� &��'}��"eI��sx����w�7�4�����Ucf'B��j��d%����H��{QĆ�C@��#�4%��"���,Pp��s�ǵ�0��� �������#9���+�~���d���J�e��I	����	�a�/�g;İx�ݿ^�5�ddv���	> @Mu� �v2�.�)���b�[>�����of�i��Vt��)����>�^�5ܷс�����͔��WCh���PH�O_�sfԝ���>m�q�ҥ�/l���FQ=����$��@n(���)()�bp��v�:؇_j+�Nf�-Z �N�OѦ�$���t��y@kG�$s�d
�w%4��q�-R���x�L�Q%�^b8߈^!��,nAb�^_�5iw�:�8Tj���.)C/�� 46*����m��C�Ń�V)�
��|"�a����	pg���$��_�K�_է��s�0X+.�����?Ӧ_�j\�����u.��]ѥ��V�*�'Sk��ϼ�{Fw8ח�޼{e��,"�-X'�N�����C�Zp��K�]��C%�o��|��봣�;��H�?���������l����E�L:�hu���|��� �u�`�U�v�y��T{k��k|��Sd�OG���I4��،H��Ӆ��A���Gz_݈M�S�?��37�>��4_J��%�C��v鸢a������A��ѸD��٪Z�Y*��?���_o�jt|\��X�.-�wʺ%A%�D�m��Ծ+R�y�-��)*�fg��,��ЎT�y��K�9��.id<ũ��S
,9}op��"��ڻ;�m�2������?�N|����L��(��n�L�(�Ai �]�O�f\��Ʌ�X���RX�`	n��j��W�B���%ѣx`�����*�����\4g���G[I���,n�)g�ђz�&S��Y�CA�������źyB�߂��awD���h��1�5X~�s]_�0��suXT�P��l���uP�;v�
g$l(gzh�iƇ��x#k儴^*\�'_�%��p�]�ZBr��^��K[`�_� K��
��\��4�]�cZs�w@@���E:�o�}!vc��|I\���q�#�'�,��� ���-9��>����������ލ�!ݸe�Y��+�d�n�ۈ�/\T��x�U��i�X	�<1���6HyK��J�h�υ�F�ˏMP�E��>Y�O���Q�9f0�p��b�=���9����`m�����D����j��A�,�o%�W�� b�
uf�Y3@SO�Lk��N5Bu٪2���u�q����[`��I0��4xE�+.�P�)���a�^����Q��GH���.)/�7߃���M�H���Cj� �rI^�i*�a�Уb3��� Zu�b?%��ns"��b�_�j�paHN�@�c˫�1��.��m@�\��YC�Nu�ԋ��XM2��	��X� R�܌Փ+���*|��J���H�԰�4D�3e�$dV����%Z+ۆ��<���ВxA��O�ɘ�p%��,�zv��4����wVGF��s:�m�Q^w��k�r�9w�v�%�X�wJ� `�kop�������4�E�m3B"im{��_{���ʧ0�Rur�p'J�M ��\[{��(���v@��;M( UWH3E3�(>x�:%&q}��6�z����D(��q�� �� ��+@�K���.%Dú��,���I^��c�2��Xϊ����r��s��#�GQ�UC	P�K�m�d�{�J+2L���?�6&�f�,����=?�����_V)���7&�%�=����ͷO�y���P�v�	�b�H�נ;�]6y�!)Q��m3��"�����m���^&u_Ա�K������K��Ҟ�6$���4]  �PZ8#�w0�-hH�?�0G��V �����&�Z�`�*�*9���,����Ā�R��E�^�X���VFE�`Y��e�A%����D�~K7��å���eY��Jq0l���Wa\	��Z$G@O�;�K�(����ٱ�d����Am�?�T>�����9�r�2��S@�#i7�O��wҜ+IR᳠�w�D��;u�Qi�@4t�	��id�𲻑���X&������th�e��?F���e�7ĵ��������i��)�����7��)C�h�s��l`��H��5ӌ�9 �~|�}"%�ɢ��
21�����JWܝ,Um �U.�`�����Yr��$�S�[�aU-V$���ii��iܤ!4�3T,�!��
f��w��i����=K���C���h�x�=��`*�8�#��}�� �dBF����)�(���fxP����\ʐ����#�V���{е͎ۘ�%^ث������YU����F
���UN���$g��=�5[f�> (u(�"dz7)���H5��߹w����&E6��oܫ73�ZA�c����H�l��vY0�"o��_�o&����T�pdyCY1]��J�ӯ  ��ڐ��E�
��&�������-��uvñ]���@���,чJ�T�MWj����[��.���m�+)P2c�dN�_V���&d�Z��0ܦ�����E��z&y��!�B��\K��/`�ۀ]�$@H�ȎНk �V���c�,BZx��U^�2��r�5�����-��W�p�'���tz3���;�,�lZ�b��A�.L��L'���4v�7e���Y��E-3����G@�3������������C�ȭR!����G��WB\�j���a��/ז|(r�-�0�:�I�H�IJ��`h9)�� ���ě��6�������3�ލi�t��]�w6���{G�o�g�*p��!��^� RF0r*|(i���I�t�N\[��G���h��:��Yw�%x�t���{% D���l�qj�2���g������4�x�L�ގ��r�~�Mo��j���t$�GC;��(3TO��_b�bqTb���;o��s��4����hFH�W���ZrE&��u�
��*���D���_��)U�p�����/#ܫ�$_�3��AFyQ{���W�6
����s�TRa"����M���_�f��K^>~4�-vV[��!{NZ�e����kWH]��O����g�������o"_K-�}�g*Q��?E��U���ɸAۄ̼S��#���T�]��%���;�t0W6_쇎�g�׋�J,�B���V��"�m�ԓ��y7��)iD�	M������ jM,�k�#;��+���]�E-��@�fm4à۫E[�� �8\��@37��/3(�K-�;�`Y^����r�Źѯ�@D^�o��e�R���_U�n���T�]#d� ӛ�Y�n6%�$3�,2<Գ*�lWLޗ=��b�OB�_uo�p�0�~�F\P��3�+�F�U`)#���2ߖ"�K�FsX�Q:	Gu�[�e�������ȝ?ٺ�L$H�7���{V��/�H���-Ͻ넦~Fq#�,j���z�����ǿ���d���U���bD��^y<9r7.J��ӦH�3ƿ�L��}V~X�G�Tso��3t��������� �Q�|��l䯚����ۨ��*�d$��V�����Xa��}�˛_��<+��b;2>��Y(�\+���7c;�,v{i���S#ʂ0Ml��J(S��9�~�޶���R�s�zu)*��^WC.	�����b�w����2Vhj4�u9WCK�r�gGЉ�qMJ̑B��䩮k�=q������on�Q�.�2���-��j��۝:,�h�<	z�y�l�og��׃F�;Q�8���G��AT%�CS=�kS����0��N�!���zpX��*�)"��)'W!cć4"�`�'��D�j,������:�->��U�����rWd���k�5)�X�x(��)�2��*)�l�To��)T_��(@�h���s�1)�C0&N�}P6�+�!I�H߆���A�$����2z�%˭Mc�`�T秵��Q���,4i唏�4
���d��v�Eˏ.���I�L���NJw��X��.�<̛8�2_%�%z�4�`���R�픜�N�R��b
>fΣ����W����h	�/�}��q�s�
��~,�n.� �P��,��K4��L�>�h����1+��5�%�5)���j��5���B���m�㥪i;6c6�o��Q�񉧠?�1%��W;S<�,�*���K����[~��zz��TA�'�#�������ջ�\?ݲڣ ��=��PpW��XE���3�LJ�=Nw�Y��-�'��]���R�zM��z?&�|�(5g�ƈXd�bUK�d�8�2ӕ��n���	Z���<��[n�vu�9���.i�5[X!'��H�e�;:"�י@|!�Ұ`�Q�#}r��a�����4�f۩��ٵ�/�9�1��x��#б�rw����D�w����
7m���s���3���9�-5�e������2i�T�v�dI�c��<�pWS�� ���}ã��{���N���0��j�x�:�=�l�{b|n��У
���{-��v�:cp+� �bw��n�"N�U�+N��f@�Hrde8��~��e��"-gar��+R���3����O��T$U�n<ЫIuʳ�:KͦJ��S�+�q�V�q&��L��.�׋��&PṬ��;�Y`�<���B���n"�2��F�/n��U�d@�Z5{�?��YP��߄x�eO�fty�}x3ت�O�b������d�6��#���UP[��a]�h7��.�)a0�T��nwԔI��ة���]s5!Ʃ=����]=v@�}��������4�8��׬�"v2�d��j��2g�D�x�o��9�Ta�HV��j��\�2��U@�!�{U%jP�w1.��VtG�G� aPxH�+jG�Avk�'�@�p��X�ED-�_l�QT�h�9����A�yAw2�����'�!lsa>_�;�.�Y�"��[�l����7�AT�o�eڽ�o��8�S���n�O��Fڟ���/ch?���ˮ��{�R(Vޫ�L �t���L)�Z�PQ�=�b��֖5?�"�ܳ�%N��J-�+��`�d��'����&`�Qj������^��� 17$��%Z��ݦ�����˻ 3ڊ�Ѯ5&<5�����Q��$o<Pg�Y�_��ͮ��yHT���@Qq��<�-x�����2Klj�S���`t�?�%��9aY��$�:]1%���[L즛��DeK�+���1��m��JZ,��Z(�
�� <�� -a�����<�v)�)μ��i��̓\����C(��Q�*���!��F��H����Ou*�=�?�*����5Bg)����7V��]���<s�"9�4��R �������o���B��%��̋G� 4:d���i�=�,�ćH=��t2��5�wL�����81��g��ʧ�v<&�YI���&��]�m�ڗN����mC�9&�~��,mg����%x��L��]�Y/�j����l��#7�q��d4�4i�M\M~�V�zĲ5�fA�?��P*�Iu�]�5��$��h���c�@k�̀�(�^H8�A�C%�����̫˴!�
[���5��΍;��+޻�_��&ea�a�� ��Ʒ��t��#P��!P�	셾J�bB �L0�%N&%�
b�Ƃ+��#kd���E�͝�� x.֋��*�Ϟ�'$R����rRք�!�ow���������Lss����a;����H�#8�X�0�r4�m�M�O4#A5���*u�z�n�G���/"�i�e,������,V�.���՝��k��:��[z@V_�����T��\N_��r{Ϭ��'.�T��MJ��IKɽ��n��d�����R�_>�w��h,~��,����V�R�STY�l�I�@U�������'�c���?<@t!�c���?��6(V�*��e��\�55(b���.7������q��7W����W�lVt"���=�$b	�g=���)�$���@g7���*�)Ü�y�ۄ%IN�z��"�f�6x��x�U�YN�& ��l�^j�T���:J#��7��,/�ێ5���?�k>�0��&!�7��#���Y�����qz�
6�'��[�����T�ob�u9���P	xO���I*o飸B@�K��aA�2. �`��5���_	 ���VBn��J�ɥ�ƿW��b��h���ߞe좂xQ��t{%_����%$���*���N�T�q��bTH�M�j�B�.7��.v����(�D�oB�e2���Y^�/����Ut�w�X�>,�Fw�v�����,����N=KR|aZ�g��@��s��[ۧ܉�̟��@:��_"�LvUsX0X�8��/cȐ}�D��ut2���e��>ꖄ�W�S�ϴgF���]�uCs�,�Q���3]���z����L��ěo�
��g��X�KC��-7?�p)�_Lq�����Aț<�Σh���ݛI���FOO;T@��ƣ���+B���G�N�d��8�,��S��Pm;۫�D�u�(_�9���J.�M�"ėꖑU4��?��J˥�1���!S���fa���VI�׵(ζz=pA(u'�����22��0��b}���fu�l�<s�?z�-m!�#RM��)(N��/9�m���\�Mkb���T,C+��!L^Q{��!��D
�sՖ��D�����9�W2�����\���Y)M)Zi��</?1�i9�s�>fb���lM���BK s;�O��p�'��`|��+���H������u0��;"�0m���;��)�E����C��B���DH @�����������:��&.VQ�#x��~�&ա.da����;��G�s��o�[����)/��(��3��iqNj�u�VZ��(H�-9��
�<�z��g����Qw,n�0���N��$(�������?W�{:��W�D��&1��i�Kj�vP�Ѽ�����D�<@Xdt����F��:,��_��>�p6Շ3��1��(B��c�q�є׮�q�a�|��9�ՋI!��q��ops�lk m��2�v�f_��D��̍Lp�3��OoͼrFbg�%�\�`ҔK��n�D[4�.va�\���!P�O��C�22T͢���/���.����C+�:,m~��6`h,�@~KWà>R�j7����9��O�
0�T��;s����{M�c�9z*��h��NE6�5�O���.��p�
zJ]]����5m���337�=��ᶀ�>`�	fG�v�2���&��椾޿�Qݶ���o�0��x���	 f)�z��X�?�T���^��W��\%�%��*�{����X^)�⳧�fpfRn�l��h��B7�p�C�Q>zi/�n���'@����ee���(f�ʦ��4ꌇ9�*���Z��x����f���������L��6�\��̏��e��5P�Qe�$�*x��f��pMh�Աg��\�t�Ί��x�nV�!����A���Z�ǒ�f=4� ����㌱��^A�Ժ��K�_��k�m�YO�k�`8Z�o�����YfL"�s�]��p��;΍���{c��.�� �����S8��jEp�>.�)�A�)Q�i�e�p�<
 ��_*Y�&v�O��Q&����9��yZ��b�cF)#Fƒ/���=/�n�(��|���#(v���'���ë�7'a^�[�*8�J���w�Ò[�&���L��R�eH����^b�X3H��s���i��-��)y�)�1�V�4p�����}�8��8���M�פ'�fI?��F�9�6����?,��!�6u��2�$�s80p*�3�y3\p�q���':VNۢ��}|eI5"�9QZ���#GX�E�~.��0���JȴxO�;�!�(�h���L��*<l 5�^:ȊS�[��k�X��A7~�$GS������ �6���2�wۨ�(�[[�dw�ڙ&�`c� ���'�wZ��'tj�E_]N��^@ �Ü!�u!=�o�0�ʯ����-��s��kf�fhO6����
��?%�)F�"�
_���N����	�^c�h=�	�s(CM �w0���ȸ��@�/��d�SPBd� ���EFC�&������W�K��������L:_V_�F��&ʼ��Vb�p3R5�R�p��ĉ͂�\H����}��	"�-��l�����!0R�{:���Ȓ٭�b��m����l!c̫�юa���">:�GH>��yћ��>��Ձ69{a@EG����ՄVĐZyp���o�u�z(.Nq)��`:P��5�ɒ��T�Gd�[ϩ��gs�s.�W��WJ�e���9� �L\0�0�9�O�3�\<�Ϛ�\t0 !s@p^a3�F�W=���
���v-&(؞�w�<R�ܗ��i��8Fs\��yZ�ef�>/T��%�(x��ewq�h.w�� U�b�l_C���ON���ֺ����y���h*9�*&ޢs��j�c7G�|�O�m�R�@�R?z��g�@سK_��r�D�"Dٵ|Qo���0~l�z��o�N�( F�A�� �|���@��"�~a�+ґ�yN��B�P��i*�z�M�*H�h8�^�5��pB�V��ᆂ`�u~�"�nyX�rK��8�6{ʁxA�C+�R�mx3!o'@�%����-�B[]JR�2��>��
�M������^���
�T�^���oE�@軌�X�NpYQI���\�r^��|���h�x�H���
ʬ�����3,�;xˣ�ȉ�׍�{ �1��Z's�9�y�"�d|��-p��I�q�6�=BK�<֯�\l��>�B�\�F[�P>a�P[�Fwp� <��.�-�VE���n�=�"�w��}8
@�(�?b=Nv#�
Si�ĸ�l5O�^��ԶC[��/n�K��k��43+�ꌘ�Hج��Q� ���A��l�������h�2v��d�PP{��Lps�{��עfV(���lz�%Σ2���7�QM��1%��k���(�Հ��<H��G�s#�.�زp����]m�o4�Kҝ���y>Ǽ����A��G�&��y2<Z���6D��~��Ug����t`t��@qk=�h=�{9�^��[�I�̬�]��.3�#�;�t�%5�~�RK�ɒ#��oq���9�8�i��o�U�6D�D���x8��O\�wB^�5� E8��p׳R�&k<2��o���SV33��;b�B:���i3�8��T��s�ڂ"�k�,q����0g��Z"��`Ax�v��(i�{每�P���{b��mb�Ψ;a�(���cЏ�o�MO��T�#��$���.*u5!��A?������S�)���Y�� ����Y��� �_��ƛ������W�YN�.��ɹ��X%9�����.�^.�C� 4�\H���`����]'쁲4������U0�@O����ֳ.�r�y!l�����^wF�X��6u6�K5:�4�{��#y����=e2���B�d�lz7�*��#�7�x }��J���4�_6�\��@�y�	T��
�&Ίֿ�(:]x�b�V' ���X�(��&��P�����"�DR�I�;|���WZ����i�T�#����XQ�_�� �l���Pt��.�撋�ZIގ��B����r���~H䠞�]�>�K@��i8�	v޿���uTv6r̕ �T��X`�,oXw]p�N�吗�6h�u������j�v�s�h��ߑn;���:󟻠��WA�w�R�X���6����ʱ�Xn����h$��l1:�+�B�`R�;��F���h�c)s0p�)�LY�	���:���\����R�6}���������oΊ�
��|{m�Pu�~f�������Qt���=J<h�U�����?�è;�m��@Q�����[��5nM�<J�B��'P�zΡ`^��ӝ�?��yZ�O���D�񲘐���D�۾[!���������J����d��s٧��@1���d����t��jB��Y��[=%E���LTXnk�":��c�C��;�w�e��J�׬����?�F��Pʡ��4�*�·�|c����<����?���e�TB�_6Z~�Wo-�Z��iBO"���	6�,���H��g3H����?�!�'�L��
�Ó~�1ypkkh��#Qk�����%���ђ���G�DПl���|Z�~-/��N�bɓ�N29��{�iKh��m=uԙ:���~C��l[K�أ��s�-s;��aLKCW׾lH�eh��WG!�v�k���'�^x4jH�Q������k�%₥*Tbg�&̊Y\Su~�v�  �
\���ygD%�!1N_���0|����z?������Y���P��~�.��٥7�[3�-ۺ�G\I^��ԛ�|\N�WL4�DGAYG�OAj�c�^Aɔ����A锝(<��ހ��K��q,��E�µ�.�H����[UN�@P����}����`k�Q�T
VV��6��W}V�z�jS�e�vf���I�Sxr��K}̍�2>������p�[Z�P�d�@P�s�jA��dJ��c,�,D��K.�x>��������E�oxK�O%\���ّJ����g�Q�+��q��
��=�p �����n~0�[�1���nC�P�mlq����]�����;1�������,@��>����z,�j��H���v�$�x@����N�G����8r��ܲ��)��@G���|���޻uE%%x�FC|6+몣6ٶ�O>&0��{�M����A��'��f�D鈰`gue��=�r�F���.�^"�l6�0���ɯkZ��d�;�z8w��礏�T'�㘣�E�f��jR���RD��v/V�Z~���B4\��I�Ю������pnH�����T211�lA]��C���7��d���i�%w&/��D�5��k*����ZM0eTh���H��|�8�vq�-���'n_���U�_(y�YI�_,?r�t�B��#d���.5!�M�V��=S��פ:I(1�L�X�-,˹9�V A5�O�'����E)d1�C�o$���>��c.�V�����I�����^�o����lL��1��a|�T���q�X�,Yj��msy�݉������T��c��u���b�����©l�O�SzZT�� ���5��F.H�P�o��)*#�c����O�X�4Hݓ7�B�b{�$�����K���-2DU2҃���R�_�g�Q��CJB*@]� ��j����yr<�C<G�g{�L���id����M��w������?B���Pr���#�N����Z��J��r�2����Ф.�`�b��g��>�j�`����|��f�����|AҩtG���,}*�!��.�]DM�jw���@h�޸'����9ƻ�X�D��[�Ki�|��;�A��=K�el`q�3G��Lom@Sv�?6��Ĝ�-P/"�$QX0�\p����
6)�i�򙯆��d� �/>�|`���.2�У��)>|1Q�n�%���l�T��=�$N�;����A�5I�1�Cq�ř�(�R�3Í0�2�Ry��4+$�Uk�)�,�k���+���<��Ƹ�T��V�Ԕ��{ڣ����YH��3SW��ᇂ8���\]�m���{�qq����e������m��I&�~��\g.)���!K	���w}rK$#�`��:|t�W�>^�}�F�_������HFkt	�s#�_����q��\WW�}��m=Ӑ|�n��~��;������T. ��!9ݺ��Ƣ/�ӯ�	�]�4c�T�͹�5��[�J!=D+Pj�ޅf}P)ƹ�'�٭����]�Pұ�V,�]��	+`�~��"���z�p�C�q�B��Q����!k:�G���O��n�^��I�Qm�i��F�3��W�;3�`��V~7�D_�$Ғ !��yJv��s����vd�P�����ִgrZ�T�CKE._�_z�݁�~�#���s�MI�|�9턏L�i)����gZ��
!�f }�����ݚё Y�Vy�`�LYi����У��=��t���\f�7�95,��
������x�� w/7%��0�o��b8���%�W��27y��n*u�=<��ߕ� ;���	3��g��]��}��5���\�h.9-P"I��r�l���f���^9	�I���G5��(K�?� ���Wy�gp�Ws0 ZQ|J��B9$?xw
t�y��鿃�J|�<�0��삝)t�#�g@!&�5�9a�oa��A�	?��Pئ��66�fd�Ů�{�h�rQ�-7f5��1<���+�.��u��>��'i4p�f�g'�WF�r����Q�8��5#r#��>L�b@x�:Fs)��
���0W�,A�1c��p������4K�y�R8U¥`��E�Q���+�Ľ�CV�N1l�� �j}Np�-��
ϊ�L��5>,h�潙vt���X*3J�P#s=���'L秄1��]Ƭ?A��5D�3��(��	���ݞ+�F̘�^+��*�S"Pݢ}�c��޻�_����͘�Q���pi�d1��	�{}�$J}KX�].WWMC#�Y"Z�XDR:���^"�ί�wzg·_r����SŜFtc�����Cc�ƙ��욋ǙG2�S6�d��~��������}��w��v�.Bd��4	Y�E_"Re��|��^Z���0�`��M�D�����[p��fEW1��_6Ӈۋ�n�G:%���75��<�� [!��/�c{���˗����d�
�f?3��M%w��9�co�yZs?�xEYRva A�vN���?�ǒrte��1^��Y!���1��Ryll�i7����(V2x��am�`tdˇ˱�
a�& ����4�G~y �=�G>��g��5HlQз	��F�%����/kQ݀?�"2�l��0D(�p�N��rXN�:;W�|�j*����	9 7�ʃ���d�����,_����$��C]�W����t�<�^��7 X�Qb4�ҥ�d����l�г�٧���WX`{�Z4V�b��������߷�"��`s���rZHF&��.���7Q�~�D�f��*qr|��</[>8���.�z�01ȬwzQ��ځ�cޛal����Ђ���ܩB!�ҙ[��HiCA�a�%ޗ��O�,�S��&�/�Ǚ-^z�y~�㧛,�7t�'8^�6Qk��G�ʎ�I�L�毿��u��ߦr������0��L�T?����=}�D�#
�����?K�/��V8�/�#�1?���Ģ���E�E=��(ݍ�+��8v�^�G��t`�pd�2L�Y>�a+��_xt?��ud�<��V"H>)݂m��~4��IZ�U�.���leU��u��L�_,��*��
[�TX9�]y2��í��V�l�����C�tf�F�50�?��5r��6�;�膖>�f~���9���i�� )�;iN�!��V���
z�t&V������ɘ���ۣ���=q�x^�g2�'��"T#���Ж��� �"�ۑ�萫���'M���H�dY�Λ���R>���9�=��]�e)x��d;�0<�x���1��F��1��&�.v��|���!0%6�+�@Q߶�b��k�^B�-H���.�d��3 ���=N�/��N��tM~��2P��� �����RqS����K���i�ߔEl�:1&��PT#�';�g��IG@q�Si��hCbi !�VRg�B�������֎3���d`5����Z�"m�P���L�>��7�x&V�<�X���ﯢ|�[F�At#���%'�S�;֓]�M\ҙ�VB
��.H��3pх��l����R����I�r�^�f�,4��to�����YL�@���ܼ����:�)�Esp�dm�+���[oCéq1���I��hKs��`��ܸ~3=Z�uq������~iP%�p#��MK��L��:�5:e��z�Û����M,���ڜ��f�c�K(��bE��W�[�I�v�k��>ߪ'쓹������n�L�dJ�P&�Y^8��#
߯=_5�N��h�D�B���)����-1�jk>����QI�������&p�{�$�����Z0�Nt
>K��g��M�5�3 ��]��C�gҢ�Aبڨɂ�Z�E����-�~Q��㵑�ýo	5�&Bdzp\�*!?ͫ��G��Zy&}J�����:��5̢
8M�c؁a����k|FG^��)�lꓕ����'��l�Z���g�fśma��/�j>�H���$O�L�+���(9�/mXQő�v�s����>r]��ÊbJ+�[E9�A������P�55a}i?��'�3�"�4��~�����
��R�$�@S=���b�mn��j�m��Ԅ����x�	y�4_^b�X���]���=���nc����[�L�Q�x��O.������*3"Q�C7�8d6�t�H���^C{���X�:"H㶜��jzfMW��tO+��'��'�.�L]��Q��m1HNb���u�QFSZB�YG��wU��������lB�����1o�[n^�:��ECB!�3��!Bw�,S��;��v���M����jhUb�է�&�a�<���a�dջKX�]�ӡ<��d������;p1�8����:��c��:�r7�|b5�������A�=���փ�"0�, ��'�?e@Y��M��%[u^3�����jŁ��z��p�:����[�tX
��ؤ�o�-�ݑ{	�s��|4f�y�����0��炕�����)A�.���|���vⱘ��w�r�=��Ւ@��~ :�\č�P�y�Y�jB�z��]�yYs�
�V��,�Q����N3�\���J�Cd����Ǯvȉ��Q��g�t���d��������`�����+���㿖�1;h���!Z:A�[]�]�� �g���s�Ab.��V����t����_�%�E�N�Ӹ� 
��0q�-�
h����)��>^�����1�$zd!$��P�)�$��+~����&���D��4Z�jB�B���$��
��1N	���~ Q)�[����d,�̾ȭ��,_q\s	I5�`�^hnM��L2�;�i?Ҹ1��CF�.�С���Y�- �jhUN)�u��75��,��q#����ܯ����P�.���m�q}a�
޵gUV��Y	 �*]����a�PO�AOG{�o'e�<�$LKB�%3	S�ɼ�c���Q����ݙ������C�GP� �=�Z�*ͳ�.	��0<=t��y���?uY�M��r��Ou4�x���8I�R-1�c���=��`k��vb�U�E�&ࢺ� @�]�y���*YHLG�x��`Ѱa\V�N��V�����w�5	ʍd]�B���8����&2G�) n�62EY)A6�p���Δ�)��_��;D[	rR��@�t_Q�:O������m<�ƆB���j\���t���<�7���B��F��;���q!����si�y�)[����z�)� �$��g��vK��V��*K�����SgU{p�H)���#og�p+�8i���LE6cfW�G���	+�d��.�Ϝ� �wˇ!�?�y7���͓�1�h�NY�d�{���ѵ����V[~u�L��ci�;�E��XQ��@�Lq��Y(~C�D�BB�El4�@E�L��o+����8Z��rfR�J��)��6��C����Ǩz��r�^�����C�{���</���N���&D����4S>)���.��[�y~��(�f'T�[;�W��whV�!�kgێS6��!� �������l3�M����k_���)-����J���h�KRց�[S���'�6Oᢩ�8���H�l~�Z�`��f��$�$F�̦R�x����Y<~87�-G�U�9졁�FZ�"e{}�	��"a3�����G�J�o��%z���%�]��T��Zd@m�����%���CWTř�����#�����4�1����*��Ls�+8��vv�qҙ�P���Pe��A:2E5Oe�<L��>���N�V�w+�9�+_�zKO<����$��V�9K	������]dz��ا� "�!H-�N��&�-u�3��H"H�{��UB5��B�7�U��c;�Q��c< �����d=!ߙ��{�g(���P�O�ND�$��=6a���`������\lP�V�����c��v�`1��ь�r/��f���%��\Z�U"A4^�~���Z��7��t��gL��$�ʨ},2
9N>����j3�+t�$���_;#���ׁ,�c�K�0+�8��>�)��4�����M�{��/0���_�����dm3W=�����1��W$W�t�>�e�/t�e�b*�5H���"�o���n��!��R'�3��զW��Wm,>P����*zٙ��ܯ�uk�@�w�Z�ߗ��u.k�C�1{�W�8k�j��o�k	�T�i�Y;Y[�,�����ȧ-�9H�	��)S�xp�/lJ��RR���te�DP�;�,�T�cV�r�7�*�7
� ��a�9e�f�*b�6���S�Lh�t0��+��	���oƂ�����}`�#�V=p�o2��ql��|�4 1��ҪV�����*w��G?֔�}g|v�~�l����H��pL>�^����f4��p3��C�9�؟��i��,q��� ��n�.l<H���A��d&f?���F0�ێ��. �<o�`ցR��!�!���h�շ;�+IB$���?
�,�>�J��"r��W�����䍬@�R�sYoč��	��Ӏ3���Q�s$����p���g0=;�z�M��l�����b�R�j�'ٶtC��F���͕$���Ԭ��N��(ڊ�W�5�ᨚ|�c�gr1��-�D�~�s�J� )Q˂z�)<̤�7�X�p���^�j��_���-���}VFn��?��?�*.G��9���#'f��	ָ0�~2��^i.�Y�Mœ%HH�?�;Tt�p1�e����8R��"���<��R8(��O4v���h��#��f ���_b����1��Q�
ϓP�(c9`�5b����&V��J�e�f��XY�A��!�-:X�P8�e"ƙ��G�Y�����g4:��q�X2Gpr3v��ސ�3 g2BN̟��c�cD	���ԉ�s6{�V�z�hB�����
V
ӆ;�=���a�)�/8.z��3��1HV��r�x6�0�ߴ��	_e<����k��uҗ���/p��ׇ����o�_�N reP�w�;�w9����Qn�+r�$�L��g�a5��6TH��]G����Fh�*�o�
���O]�Q:���'�r��
���0�U���Mi�n]	��	���Z�hͣ��%c�!�}#�Yr��v~us9�,�GΉؑ����܄s�0�n�Wq�ʳl�g���dg'g֖n���m�����{(gqЭ��nb����M*�p���K�mm�b���m/M�S40$��P�Z���}!?�����s����!\q��r�ᖩM�k~\z����f�����/	�8Q�����i���m����M�{d��}7|�$�utP�]乜�8�ڝv劻�nW�;�I X�`�<%����Z�U��J+d�.�h����0Ѵ	K���<�&4���l��6@�ߑ����KΚ*�"^�<G5[�C<�P��B�깙���	䟋�9c��:d���ղ�4�b�2��~�M	�g�U�����,��&L�0�aL���y����U�I8a��R�8���.���cZ��Qೀ��ۨ�Ky^� ����Ž��;��)o��¼�s��{��k��X���L����e�����<��P��=s;�������N7q�Ką�J��[ʽ9�6}�e�Kĸ�:^$���k�ϻ t����BBs�G4=L1a.A���@����Ǥ\P���IofڄXڻД��@4��}���h(7�t�pHG�]>�\|i�.��D�h�V<������Fy}�u"I�)n�L�=�ҪP�A'Q�׎��q�J�����*����w�k9a����)�51���e��.�2/�i� ��(�$��q`1�nv0��u���$[׈���E05���C���`͆8�0��\$��?� N�\���^��kᘝ|��C�d0j9UA�	�/P� ���p���3�*.�M������c[Y@c�c<}��V	$ ���ΎDC�������{�=��h�W1¹ v!��3�_�uA�4���-�t��l�zAjt|�rlHb����#�gіD�mng�3?�PDՀ$o[7����+��s��Q&#��dw��-}�:������B:�ك� ׯ��Pi�Wo�44vVk|�I��+v$3��|\3L�M��Q�c"�ߗ����}�+��E���Z��!�i뻮L�c�rc�"�5��^�X"~��9�M���E�N�T��b��Fʟo�R3!�x�/߲��-���Uvmk��a\J�~К�!/���Ͱ�yD�#�Y׷ӕ��e];h,R�sX+���tS$^S�A)y���5A�Y2$�W�� �	uR�[	΋�%]YWS���I�=%��8�5�B�5C]������/V�#ͭ�5/P�G��MAN��,�\�a����I�m�G3�9\s�]�Z�?���9c���U�¸�uCN:fk�(g'����'��ݢA$��۶����a����9���}'o��L��p�X��HW׺wu�8L�V�I�N2�y�\�%7T�v���ֿ7�ƙz�~�#�z�[��v A���AM��W�-��z�.!��{_�d���ݐ�M@)�����x�P�Pv����� S��2 b^�{�-��]���c6$�	Nec3���vTSr��@N�8��;i?M�(Q�vO^�8�ZR����$�H��dh��BS���T]Ů`6Q��R'�0��,^Z�i¨B�F�����ks�6��.؈n27Ы���3!�[q�j�����3a�	�V����3R����k�����b�0J����my߀Pe1Ti�������Gnd]�@Br#~W:��ͻ碅7"K'��r`�`�+��x՚]%���~����<[�ۇ��C��-��/�ۻ�9��
O�b}��*Z�)�o&R5��J��jg�HxI�p����#�d�Iy��lkl�T��������pE�;��P.��ؤ�Wd>���~�I]������7?��0!�Z�'q�1n=�����"���_7t;����Tz�3�%�� �+�
T��j���ϱ8�����f�ͳ��9�Z��n�����'Y����[QCN�����fߐ/��b�<�U9M� 3V9��5@�E���7�N�;8��S���6����tb�����Y����{&�&�V�� Q#n��%��*���}b�'�J�z��0�i~���G@��F���X�8_�mZ��w1���R�9���v8N���]N[1���Ȅm�����	 ���F����X�Xbf���U9筏�5�`�c���4���3:���ȗ�t�͒�-A.��"YFO�Mߨ�3�&��pfQ�:fo�^x�Q��g±���I��8P�%��|5�
�E>�:��#T�j��K�_X6ӵ�m�s���,)�7bV���9�=����D8�ق�k�]Ir|Qj"V���^�A��EfI���VU���E��55&����6�_�ɠ���G	�SG߶~�($QzI�n�>�Ro��i4��Z%܀�tX�=!?aǾ����R�'Ǖ[�>E�2|������|�@�	Y�,�Wϯ�׵.��7(�>Y�C/Fk����q�}�R��s���B�i�ɣBq�q�&�+��N�yZ�����8R̀��9I
ڂE��N������I���r���ar�FV��.漎�����h���+s5ڕs�2�WiX��1g��2����]]Q�.�0/9 
�xE��v4��zr^q4
��C�^�S��3b:���x�E�;(��J�C�UI��H�4����S�����+��.k#J�LAX�_�Ϩ7�O�F����)�����ʅl��%��
G�F�|yH=��?E�̊����{Xe��5�I�U��@�����\/=Ɨ!�3�I�Ĭ"��O\�R�rj*F�Nv˓�F"���� �_�*ܻ��'�L�9�y�������q�U�kN�8,�~�h�_7A����7;KJgo�w�L�O���"�D���
����uD��A��2{���y���6�ʠ �V��Q��=G�A���>����4@^	PӃ�fˠ�:�"���a�r(� !��o&��X�-�xQZ`.j�z�[�8�Y�q OJ\�
I3enN�rPoCeӞ��o�5��64��tv�e���C����t�OJ��أ u@e���5��#2�eX+�(S�b��΢�)�U[n���[\�t�v�̼���V�9����6�f1@2�/ 3���m��e?3:��(��.TH�R./v�"�G�/���g�p����I`�l�/�����s^�z�|�d��Z�͹�ha�8,s|�]r���I��.�d{��ʝ�>��!��3��t!�[�z�w�* �ei�e�ne��(|Z�-��2�u��^� eK�7�Fa��ܡ&����?��6!g���'f9����M�������̼h�AZ8d��H��+idїG��3���-x��@��V޵a��������-]�q>:2�>!�a/y�VL�̶m�Qe,�fAaҥwk�%���c�N�g��-���T�K�HR����}�&�=���T񻐤��y�UQ�p��v�t@p��sPr}���B�L���L����{T6�˶LG�����ts��N�N��cӵW�D����.lr�5Cs"���=���7nr��ƃo7����)s�7���xl���/��-z�1w�|����+'	��h����!Z�s�+/��TU�� {HZiKQ�u�ُ�s�I���c�#�QMb4U�*��Q���jm�_�^��H��>;ˈ>?|�6��U�{�X�h<�G�u�v�� 3�Ɯ�u�(��ٽg�չ.�f�6a��C��,l�M�l��'��H���x�7��s���j���Kq_�ɞ���?(A�BX�G�OE\K1,��EPN@j1�����~>J-}��B�]�e�П��A&R.��<]Ǉ"`�E�ٙ/�4�-m�ӠxЅ?�,4��[�`�����^�e�) r���tPMV�����|#�ٓ\��Ɠ���h(��"��B��LRC���CV���!��	p$;���R/@S�#��`�G�)��Cǽ� c ���w�c�������o�Ry����U,'��\\Ʀq"�~��CU=
N�)'��4�4Q�Wj���l3*,'��f��g���o�P&�gT��]ٿ!��iQUZy��x�Ȍ�@{�z9��J	H9�5���@���0{k��@wx؏'�NkxblPn�w��ʤ�y?����Қ=1��
��^�`��4����<QK*��};��̅��v���W�m9&�J*�B����V���T��{�_9��yD�}��w y�W��u��]��0q������w��sD{[<;p3�$�c�2�L���wy�
�����w��K���G��9���r6��+��^M�P�Tv�n���VsW�D�5�y���z���|�Os�.~d�5�\6��bp��ac�Hʧ~�f�RT�i݄��1e����YKѤ�RV���ԋ���^��=�P�h�f_�����W6(yAa>���~��x�ޑV��2�0��v�/!�Xd3�_��v5�/�
��.��~d+�"Eu�}3�ު�f��9��A+F����X�4�˯����|u��Mǆ�Ǽ����=P�Ǎ�z�lԟS�Yf�)�9І1.?�h64^���{��]�W7�_��dqX���+*�#����q����Z�tҗ)���N��[�KܗR�� ��Y(W}[������m�Z^k�:��]f���J�-��,}�y����o�G�r����QAD#�`��A��'���^e�"gNئAU�@�爀��sc�EP�-��0T���=�88�.��A����b�����Y�[�R�b�I����%��A�r�]ؤ�8@ά+��{�kc,�Ø��Ѥ�v���NQ��MԨ(��v�L�����=��J�Hݥ��N�hE��v\2�D��uue6�Q�mgϒ1D���
fv����[1����G����#�G�]�K��2�Y���`x�O�AH�}s�M����Ғ�rz`e���ٔN:��H�����>�7�(�c�����Eh^ۇ���C����:�7N�l��8-M6qd��éqL����.�P���НhեS�����\?�]���L�����l*Ab#;/��W��ݸ� OC_D=B�&l�aV�6�Ȱ*a��HN
o�4�k�7��m�ʼg<������9���]�����3���zq�H�ĉ8#=R��-:Y!�1_��O��M[�ğ`Yc._ڱ�����j��s�����lۥ:��<��8���M� wfY��%{�M�`~������1�{^���hQ��HV��a�"Ä2\��Lg��	OR�-�Q����C�{�~���y�>T��}|�iD�^*��'��c��􋕮�h�w�#�odi�w�K���M!f�jUǸ��1�\+��s���1��@{*��=��O8����]��(�X��0Ć��Rj�5���|�9�`��]ÑEr�U#!�vmۑ���0ώ8�9�iw&w�&2D@��^E�t_����Z���S��:s-7�]EW���R[q�jQ�ׁn�Gk��L�k�E�b�4g�=�Ay���;��T�T��0�]Yw�0o�LJ���u�������^.0W�ئ�kE���X��ՅU#�y1�Sv���HyKyf(N��1O��W�L#E�{2Aw{;�{�t ݜyU�����nS$!����Gp��י;�:X�?G���rG�K��qS���$����J��Y�M�B+h�,ǣuiC�9-��4a[�^&N�2O�,�sW�-|����-g	pb�$��$n������2ۛY�h
|��{�
vk��z��f���ʩ���_�صOq%�s������\��g���J��O�O�߭���{�>l�V>���i�s�j�^1̋�b���r�ֳ�'U�"������w�m��ߡJ|�9�^���Q��i;GCa�v,�����q�~^a�:[�v��]�-g�f�Q^�t�"wN� ����3.�f<��W��䖩��کwЇ=��Ԏ�K���K�S��J2{�4f���Y<�B�;+���c~��]2l��;�k�;8����O#I�6�@�x��GV$B�
q
'����Ybg�ݜ��ܴ����` a��+Q������[^�כ����ŷ9Q�"4n�$�H>G��=qw�{����0�y�|;��i��@��y1���2�t���Ɇ6�.�H>X�ɚ	B�`��n�Ki�U��/�W�����f��l( 6�+s�����*�g?��Ө�W]�s`�P0�N>W��>��0��_]\"q�� տ����N��o��2����*Z8�����]�����_ӏ~.X��H����i��hr9{��?�ܐ�����1~$>J�@�����Il� ��h荚�_�.���-?!P�L���5?�$8w�:�蹤l�$�����JF�҉R����Y��D����,�ݔ��:/է�'�*B]m���N�n�e/��J�G�b�Ş:5�'�9I�<�O�~��SW��U�^���@�d���rӭ8� ���\�<.Q�G"[���%	/��z�?89kLQ���-uu�t�^.� ��sͳ��~��mH�uX�pU�D������K�o���o2 ��	�@�m�R$Z��Q��>�ɱ�	9�i���@��+lOo})�K:+A��dJw8��!ilσ���&9o���$���˛k��,S\�D->���-�`�I�/Htތ�`&�oL��b��`V�Ӓ!$�I�ϖ�����8p
[S�9��Q�ĆϠw���4��\���[0�z���Te��DT�Y�ݠ�I��*m��� j�B�=/3�g$WL�7�9z������dz��ב�8��bn��z�V0�Ld�*��Ĭ�Z�?j�eŚ)��b[����+���;F��<�%`��N�����`?�\�;֧ºׅe]�[)8E�)$_ JAl��䆯��dU,zF��,�qǪCW��}cq�U��c�)�\O~<`h�ԇ�bS�y���9FΜ�W2�J���/��#;�Ba���̟���ko ���F�T�AZ�8�S�����u�N���!eE�wr�Y��|�j�BNu�}�����)���_����;��Z�So�T���k���^�'M�A�#�6����66���z�E��[��:
�mI~���Y��1ED�Q�{���sV:��ύ�5�zMJo$�'Qh��x�N�`#oN�S�*�$;�lH��ζ�W�dH�B�V�:�s �v-lᒝ؅�BQ��4������C���#W��$s>���ng$Q��(�J�N-\��,8��kb�F�_S+ĭ/yw�{5� ���|BCE�&�����DaC��T1��r@n60�Ɠ�9Z���������&�<��8�d!8X(�j��~m�pH�U�#��^	"�2Ŝ��/�Z�,{�.ݮ���B;y�����79�T�<�Um��n�G�}pA#:ƅ��aY���'Ew�A�N�>��Y�{*Z�V[�-n�t-�ڗ����hI
�M$�̂�k~��=���0%*s�Z���@=����ԑ���q6��LcSCW���V�}�g՗ZnVG�T�"6$=,ߛ��[Y��0 V+�w�Ԕ�i�L��]¹�ܼ��]'g����0��*�He�u�4I���H�D�9�Fr�ly�>��^��/� �{a���|(ۇ�X�o�i!Fҵ�ܒlKLۖ��)<J0.�Vh�/����LpWa�0����=`��C�sp`Fc�C��`��s8?T� ����Xd�}�o=�Ժ��mG�������������m�Z\��]t=�Ⱳb��I��f����fR!>5�iת����GI���%���wkٶz링E�Nf����^.�?���bd��CLJ�Mw3��Ο�yu�q�F��v�Փ!�9k�e�m&��{EK�$�m���ϋ�H:k�^���v�����%�U�����M��������rfV�G�����燷�@E�<ʡ2"��n���Iۨ�{C���>~U�.�)D�4�������`��yE�VX����"�}=V ��������W�()�{=�v}��	�ډe���F�#�����tuqF�Y/��90m���lw�
�Ab`�P�����A��\[�_>� e��Z�0�>����Dݐr�����5�#ў캼�Z�|~�Z��b���p��V�"���j� /�<��d�wlm05��1��ၱ&5p���&,l��r���f�C��������je�&ҁ������<B�&�[�wp�)w'@e���+p�2Pܪ�Jl��f�#Bb	M�N��+*1^&�x
l�� �L���$���:�H�S0�<�X\����Vȫ~��3�NrC��r�w�/����1eH⽖>�;�+���m�񿜄5���2^`3wV���n����A��??.^����]����~�/�E3��t����֊��5>xl��	��6)n���8k�?�ʝ������\|�쏳!<6S���\�4L���g�S)��{sq�����L�e����95J�˺G���k-�4v�QZ��.a<�@����86@��~nB���y�p��@^�HFfb>������x��"��4�%��_�>��q�U��|�(�}nS�穲��	�R>��O']�L���E{
�8�P�����a�w���7�B�������e�ԬD� ����6I�>��(�$�tf[��a�jq���Ȩme�ӆI+���[>��V ��j������.�<2��{*$����<~�Ć�M�\�w�i� $��Oxab�(�`�c/�P��9�i��?�%�������+^s
_6c�n���ݻ�!I]�	�ҷw���g?
��H��G/ȓ�-i�,���حJ����n�_�g�FW�|Ѐ2Z�*�E�/,Pero,�P�����t�:�Y�E<�=[�/���R=��[V�8��_��w�h(��G�q�r�9��=�Jwh��G�����l V�����?�T���[��e���%�y��Z�s�"v	�aNy�����Ÿ�[�$�r���E������T�Y�L�����߅���#�g��&!�r(��%rp�ә聯�
񐍗�"Ӆ�^5�v_'Y�@gI�)�X~F.&!ǬJ�G״�wh�΃�`�D�����r�Ţ$G�w�c��46���+���jU>	fB�XK��egf.�ί���&t��	�F{�T����P�y����k�H��S�*���6�������*�Y�݂�=D��:,�<������I�?���?�=nѯ{��Ϟ�Vy	�8�V1o�����P$�Ll���)�F]�O�go�G�!T'u��o�I���LO��B��7_}6-g������i�Y!T��mra�4��8H1����$4[�SW7�N�D���(���2�ڬ��a�d�f$��k!��v�d�*�ω���}=��(���~��L�S�Z'|�^c5z�]ZH~>"#�j����
�4H��#�%�
�OO�EQ���&�_P=�]9$E�_���b����G١��Kl��)5%�Ai		���G0�dv-a�aLaTQM�� ���~R㙗s@3��a�'�-�StϻI�PP��0���r��]Y1���͓�J}����3+FZ�:]MWO� �ҫ[��TX6;S���e-W��1UN�d�o�J2�O��9�����Z�w�!��|nF�t^X��޿,�����u�W�HZ�a]/S�B��hp�<�r��5|�Q������hZ�d���š�N�oQ��_J���zw��Q�t��3O��"��Bσ1�*�q��
����'���,^�NP6'=$�9�BA�r����ܩB��	�KXc�iE3��
�(�R��c J8~Ƞ��D)��B*gEʫ"��������l��½	�̼W`� ��SN��.1|��'찼n�Y�5/�!��2%��c��<����:h;�J�����l ��V��!��U��i�1��m}��?�|܌JM
�����ז\R�%.0��n&�n#�6�_�Х�A3���٫�=��6&%ql�9�oZ$��+.k\1QJ��q��z�;v�E.
gj'%ʿ�??���)yM�ucl�� )!']��wP9�(UEK��\�z����:#/�Hz��oF���W��B��%R�5Gi�@�Ë�-%��I��Ț)|�ƶv��w�'�}��t����:�gk�Rk���}�{�@t���d����|�t ��p�J	?�,�����9���Am�Փ��cvD��������1oQĸ;i�\�<��9n�a�n��TS��m;�=m�m���Z�B����(�wf��'����y 0�a�}�s�CG�� ԓ%�x>����d��̚�z�WZ(cqk�\Bk�o�&=K��<���G�U��'�t�Y�vm����^��(T|�a��_9.~W`Z2�ՃI	�P:]��~C��?'%]�*}�m ������P�3t�1��m��tP���M#P<�m����*zB@>��yU�M��/�k�.�%l;�TCoUho^TJ�$��ݛJ�y��=��_�ۤ��wi�|���<258�uWUQ��V�h�ڀK=�o�Z����v����KhC��v����傪&�яʛ��E�(�	�5'��M���9�׳�p����"f��c5Y�}����V�"ȟM�>�T�-@ N�@���5����bj��Y}�����@�nD�ce�0�@(\n@��F��/t�l4q���i�ll����2��b[M��Υ6�A����3u����GlRHV����yn�c�D����^��jO�w~��n��_��Հi�W��znEe�ji�{k�U��S#9d4z�pHEr4ˌLC�s[�\Z�>��0���" �&ڋR��x���&��S4��pha�j*Rthl�j�� i�b��&��ZRcUv��w��j5g�
T�R����5t;`�ȝ�m69vt��[9�z������'�c��dι38s�t������B�׉���yն���4<>�m؋��7���$�p,�K��Nb�d浄N�
�<ݝ4/d��gs˛��C �;E1�c9�(|T8NE��k ֳ���>�d���9E$Il��	�/�J=	��Pu���+��)�a8�r"�8!xhL?��c�m�܁ /���,:�h�U��l���w�F�痏�n�����C�z_V$Kk%����b�y�dM =H�b��.�U�xɤ��j�gzM&d����$�i<�{N�j�ʄ[#�!3�P�~*��/�@�af%�;y�q9�t�5�T�D��&���p�>�k�%���(9'r"0gB5y��c�f W��3�P��HR����'|;D����4���{A#F�V�R-��sq���Q,Q��heُ�qWtXι���^Kky�A8�{�3���*3v�xp�H�)w,+��h�Zt�r���P�c5DRV/��*	uڑ���}�w<�u�uYg@����E�tE	�C�(f���h�?��M��*�3(���K�X��Sj2cM�K����%z���	�QEg�3i]���~�kI;ލ}��)�_�Xu��ȅ��L���k�������3'9s�K.���K	X$0*��"��im�S�4�n02桉S�L���K�4�._�٬GY��D(�8��}TZWPd��o��g�AF�\���$�ð�O�*]sBF<t������R��#9��[�~�ri�Y��"������'��^R���^R�-�^��ZM5��~�J���U�D�xP�G��Zė���mL��2��jլ�X3��᎞��C�u]�3�<�*ۃ���t'?	��-Ҕ��I�p���s��i���{�A�5*I�����x�X�<ԡ��0�>��S�nlT�	��[T�V$���
�����}�/�wֈ]W� ||�fr#�y���p�Y�ʯ������5�
En{ſ�n`�ؼ�!�}MU��fצ�����U)(PFT(Y}U�~�dLo��=q�����NC:5~�5
U\�?�Z�����&��t��4r Xn*B��<yi��*J�����5g�+�j�J�Fֺ;�âu%���Kא��y�l�^�)�y��z��}V~�@1�X��	3c# mn梨�c2L��+$N��L�Aɟi4؈�����4�LH�5&���=��Ŷb���ǝ�5| h(s��r��!�nDU?����m�<?�M����Wx8��-��+�D�������p̊�zE	�pDQ'�.�v'Gd���\��YD��B��#Nx\�9�W���}����Z�c�@]��y���6�d�g�~Y�u��|c>Ҧa�B�:U��4��dj����=�M�$c��1d���l}*��u��R�ۯz��:�E��t'(�*6��Y �D����x�B��H���ƃ�A�;�8 \6+���9X���O�`����Naj��+V"�C�)	��{�+J���Jѳ�������A���2�G�Sy膀�o�ot�zbS����d]3x��l�:�{;�'f'/H�S���)� �͖�m�D��� �c��;VoVS�BK��騚�a/(2��Gx�Pu?W�w=��ep%��6�-�Fx��~�}ro߂�����~��܃�$dZs��V���r*��i~�G���e��d�&HRr�:z/\�X$�*5��b�5��PV�b���ˠ[������ft���ߩlG�$Ƹ_�*/��[���'��V�A��6�V�gC�/�Σ$��Y�7e��>�kbX0�d1'�(Te�}"���<�z"���%xhb؍�m�~���)@�/D������U^�I�A�ȡA�ܣ̌�/O����u�ۇR�]0���L����q�*V5�7�@��+��3Cxͧ���]���D=�V�� ��C��$ߵ��t鶟XQ���*�V��v^�8RF��5�n����u| )(j,yL�Wi�LN���I7��S�J��x��iƒљE���c�h0���^s�g�t"��2�>��3N�X�������Yk�T*]bx@R�x=����\���D}���d �x�T�u=MV�P�-g/��6iX�5��RG�UU��,rA�RUJ��F$D�5p��2����M�ײ��O�|���d�7�j-oa.��1����X�Wbh��v��h��E��K�z2�{8q����l�@%����v�����׭-�[�I��
��j��
t �j��8v/Bay��$8�.�/�a,�\vbTn���D�T�.�P��1<{uD�����LI�zK����^Klzp8�cO�b�������i��9��QJu}͹|R�͠�=W�׬��=�3)���&����Βu��H�l��g���XJ�$ �4T����R�.����L�!n|e	#X,!s��5�Q���U�� �)���h_���u��Y/��R�<N��s3��Á���㾐�-";�9 �z����L�ɤ����7�W�>G�@~m������y�n/:$�����J���v��ٞp�!��'�%2��ݿ�6��n�=�u��g�t����%!������;�<��Y�=��$\y�<��!�@�1�
��i��S�E+`č�ԓ!���u_�=���=9b8�;�'���ɀ��S����&�h������n7�~Ƒ݅��|��yCJkܵ.� 
�Q��}��0��s%S���(_t��Ԍ�}	����C9�Ц[+�DH��&~�par�(�1�'����c�(�����&��0��J�_��ɳ�Y(e��^X���I����:�Q�؛J��ȴ\S��I^[���T�wEn��Y���v
�DQS�5��pqf�S&W��I�*'��Eל��"�*]w-"��Q���ڌw�Y��Gnϡ�F���ٷ��{��t�L�SD�Q�/�!�[_'��T" �߶t�@Ӭ�]�u���D~Y����T����-}��.���T5$jo� y�B�����vyG�Ļ_R�t>7$.� .Xv�LZB>	����5�#:�mj�A�g���)��w��=f��4�M���_��6�b�)���:����Wpo���#��Fp����/-�=���
o��h�*N7��'���ļa�FqWQ�%��J"C�B2x�i�����6:aR����@3�SvJ����ݒ8T���+�a]����������ר��~�8k�%���z���i��q���{�/���E��w���eպ�+�.�Iܝ�LbJL)_	ӡ����2g�'�m�$3�є
%E܉?�-z�b��#�O"����&�`�svkXě^�?M�{��`+��%ߎ�����?���4=Û`u�d�#��{[?�e��x��S�y-Tȗ �*9:����Ā��'�H���3��&5�S�&ў�_�y��C1(�D嵈���d�N��L��������g�2*8���� �rK&[���.��"���h��|C�l����@$e�>`�sl�",7X�z���0#J��0#v�+�~ޯ���j��+��5����[���ݵ`h`��[�®4��+��d�;q�aw�̸jJ�պ(Uy���W���T$[��+j,�����&z4��I��^eT������T3�czݏ ��}Q��t�3EReޠ'�5�nl�,�� ��F�*ƗfV/|��S�8�b��G:�H3�ls���9al�M�׉}ݏ`�'���=�:B�C1�\~j�q)��+��;f��$�ដ(����>�{;���	1���+�Y���i*)}Z
R|��k�V2��ې�1��<Kb>�}"�|dej\��7h`ٲ�M��%�#Ү`����bn���� g�_��e��m�bo�wez�K>A��n=5��7/pWǗ
>�>�={X_b�P�.a����pُ|��k�Aj}s�.u��TS�a�2&���dy�)��I�B7�8e?7�N��9�w�pP��c�O)��e�.u>x�Q�Y���'����'vw,����-]�|U�?ѿ�c�� jef!$������h�`)����/�z��x�e��\�V�y�@1R�����3X���(|5=�P���S��K��g����=[�A�k/}a_b���Zz ��CRX��7�6+���$�"���{�*rT��P�ZI���≄��4��͜[��0|���qk�����.�Q;:����F�,J�!l}��qF:z��i�ho�S#��Q�Iߘ��=�nSg���6]�wO�Z!�5"��g0��b��}��c, ���GZ|��w��B÷�2�Ǭh�}F>��nI�,n�3$$X���և0�KP�f�|�ܸ!�6^�%+�(RQ������z�uO��tE&u*��s���bI��V����k��L��w���{GU���H��G 5��c��C�4:�����˱IX$ı��뎏Q�����46~c�Ѩ=|Y�9����!iΎ#�sxS�A�	�j���|��a�	�٪�c�C��!~R�@s!�9ߓ�fa�o�c���v�ƷNj5�B�IY,��"� ��!w�����&�tԼ�E�M�b3J3$z�����*���ldd�י ���`��\�]���Z�"�[&d�9Y!��^�1��'�}�Z�f�X�$Cm2�˪�bQI�45���_�6r��E��#ޣ�ޘT>KN�U�j�r�: HL�⇅}�V*U3|EJU�ޥ��X�������>�5�����p��<�@t/ݽ�+�u|��@����������6�D��I���ΊT��7G�]��X�?����UM���$:H��̝i���ۏx�F<,�&4��������/�c��}�	
�O!3̟�7�3���P0���4}D��Ϲ���v��h�=��;��{Ȇ�)Z'�;�OR$�>�!��|*m������Y���㈞�/�h�:�o4A���Mj��h⠡�|-�����g
>HY�t7������6"W'r��;C�K�E>�|#z�X߳cw�Flv�6z�ȏ��k��Ћ��ON����h��.ixX!*ӹV�,c|��]�YA"�Q��4��"O�q�|�hR	"SJ$DA���N�l��'	x%��J����dg�w5��E0����DV�1o��c^�ǰe��-v��362� �L�����!RW�U�@;)������h+���r>�
j=�q��V��cA0��z,�ڌ�x�����I�5/߃�Vo[Zɫ* 5 e$#��l���x��>5Z1|��	<��c*7���Oo�n^�rE�Or,��6$��ߵ*�j���?�i���6����M���℻��X�R8s�T[nL,��W�3��;ĴLc3U�(��K���S����"YGHTs����u�^��.�7WK�������́�|���H�*u<�G�l�5�z���#T���j�t*�O��t8y�{:���6���\+�|���2SE2������M"��t��/���\���,Ez���xu��(�W�Ql�|�.h�e!<.G�r��M�H�^���U" ��{�(\�z��[�g�(,�����=E�[����o,#��'�gH�؟��V@&�y0�#����L��֕�O����ܵ�m+W�M-��Hp��_-ҕfD��3�>����v��\CYЗV�$"7��N�+5�@Lh��k^k��n�+瘏���`1�c[�&@AGT��Ѷ6	���co��[�l��29�Y_c�򒗱��k���W���h	�Џ����{�*sDM�k6�fT�A����!�Cv����M#��dS�F���X-�pk3ɒ�:��V��2��<�����F��i�e)�H��p��&ju2F1^���Ħ)U8�Q��!��,���]j`�9}
�.ɏO�H�opn��ZFm���Üc�	�[���f�n�4Q��ҹn�|�^{�WvG�7�"6|��Do�o����-2��Y�}�<_A��B���f��y���4�����' �y.�w:%=|�p�����[���V[Q���B���S�܍!�R]���NT��3X.�QK] ��V�C;9���,�Ŵ� WNBr�4��1y\g���)�Y)�Aq� \oeRx�G�� D��pf�&�U$=E*c�A'P�(��|�B��_��i&�2]��Հ��t3R�i�j��2��SB|[Q�wωo��F*�JX���/3WQ��u2�*� >��h�Q��t�G�_YP�i��H�E�K��?p��@�\���-���U
3�J1��'jY���yՊ�a���n�0�����ѡ+��'cׄT��¡��H��Y�)��z��*�MLP�j�=:0�W��p�ѝ�lV�u6f=�>���{3��=H\б�Gm�>�{�	'�S���	��胄��t�W/�8�s�+��j�������H���^OY�8����!əR4%�9Ϡ+§�����-�9�zU?$!8����>γ�lT��oq������w"(h�{���R.���i���"�	M�G���D��0~���+���vP�@���e9�#�[*���$�u�>��hmE��[��F�d�q�fS�a�:��rՆ���-��p�E�A�{�ʏ��]�D�LP����V������n3Lz�A�|�4�?�6�X�����X(7ગ�"���A�0�I����_���lrt�X��q�M(�|Ϧ��1���L��3X���k ���M4���M��rW��$��w$C�UT��Bp�G7�Z����g+D� g�R��;^Y8�1ط�ZfHG^H��a��V!�>Y��8Y�k��p6P&Oe\�1r�dI@'/�������z[��2�*ea���00�r����;��3��uj[w!%��H7�W�'E���r��*�&��yo*��]�\�,<��*�6:�ƌ���D��Ey�_)J�&�no�m=GFn��%Ռj�NT���"�v�����XK�w/��F]��*$i¡����+��̶�Y�e�Ι����(u�1�`����@�S��������綑�
���.��+�"����.��p�t@<�;Ր��|{�Ln�r�H����BOq��P=q����D-JJ@9\sƎ���p�	�c a��E�끦#����>XD~�&�w��U�`�|@#�Ȇ�Jd����}_���m�%�lΤr
.,�&K9�̬��1���g�:�`�a�RS�z��pb�Y9����[_GŐد�W�d;���T���K���N�K;�cc��
lo[�5����O*���*+wC=��_k��ִ�;gY�w�㵙�z*�U�_4{7�0����Q�|S�
��bd�|u�Y�����9�ۘ��S��ڷ�<�{�;���q�@w��z �̜�;��Ј�TՒ���M����I6$�&��t� z�%u�5 ��s�L�#Oj 
_���5�̵�2#��IE͋�%h/W��>ܒ8��m���qŒ�_�[�Ʌ���A�	�AE5�~u��jKdG�7��F�=Nx�ؤb�.�;A5����cߎK����?$A�1�D� �:F�44łF��<^Y�}�FZt�+�Ö�E
�4��K�u.�����!Q�����|�t;�0��b
�
����CY(�izEq�y;��t�_0�؎�v.�Mr�8s��oz0��j���Єj	{��Q6͑�5�
�<jW����v,�a௖����z���}�-� |/�r��?���S���[�Ij���2]�7���@� �;J�ژ�1��r	[Q*L8.�'y��T�=�nk}'��5�\0B�r]��ߚ�����F�8i�2Ѧ����Wxl����zz�������U ��w�yf\L�Ծ$��;DC�(�!�=�e~j0-��%�n���1R2�%��XD�e&=m�&���"��t�Iű�T��	����c��V�̀��"��0�rnI�� �<�O���I4j��+%ە|�9�xj��Q��'EV�
�t��F�`�^�x�Y�'��z�[���l�^�G���H��"���o����Dꐏ���]�@���E���GI�po��[x�G ̈́����^Wc�t6 8�@������ϧ��zQ�_�36/���סs?�0�c�U��T�
��Vm[Sng��<8�|zD3����=f�kƹ���o�kY�<N$U�چ�:�l]��w�<��?O�����6gKh������ܿ,����Z�h_���@$T��c&������Jo�G�0c� "7v���U�
)���X~~aj���Gdh�:��v�3����|F���l�"��=K��~�1�Y�vJa˨H�ֈ>G��L}�U:�����^�B9u����}�&�b����;�V�0Gv?�Fx<��N���-l)H-^a�R��H��-ٶ��{��Z���.\�W�\��?���Y���=r�n�_Dֿ�C4�m���r���P���/C�Q�&����:�֦��+��{��~>�u�"�������(�(�CQ\���-�m�s�aI|��!�?;cR
dy��<� ~���]!��ѹ?���wN7H5	�t��D���u�n`|4\����7���*�H�g9+�#ߣC�Yx~H�z�񉱚��{�"?���`�^IL	���*�����.z�)���wj���!3W���D������t*y,�q�/|�μ%GQ���@�[x,qv_� ;����p���sH�훏��cw��+�����i~e��U$sv��1K��,��w]ӈGA�;��*bpSSq6NW-��X��?G�r�s#,H��/�40����fDz��i�K����l�)����	6�'��n-Au�s�����2�	��#z�T�׈VX��5u�~�ۥ�5���+B�ę�-��a�e�B~}ğt��!*{�>��5�d�V��u�����;FSQ~iI��+�JN�+`+�s(1߆�q�XZ���	s�yY��'b�QE���ϝ�x�� ����UM�SO�g���|.�T�0x`����<˿�^�e>��F �r�BJ����S��U��əm��Z.f�.x��.e�2��J�\��-W0<_W��LQ7S=�]�R��P�W���a��Pe������ɮ�A�<W���A�p���_O��l�
��$���/����e1�r�0�dc�є#j��F�$p��0�<�ݫ+)��w�-��,�������b��w�����	��߻x���Ƽ�rj��7�k�2��C�Z�a
�6)W]8�X`{[`�4�0o�9�������$�)(�Ey�[�D.�#��c�C����\%�q���ZU��G|#(������F�>ZvX��f�zn�$�U1:H����̧�՛�'>�줝I];��`׀$�U� �D�}�Wq��񢣢��}���>3�
�������AX0���;���cn����Ix�8u�>g��m��fb֭L��I��q+�'SȌ�F�b���]ӀL�ȕ~x����&����B�������_I/w2�'艃�.:�u��)?���k.u���o[�o�Z"�,�Hm��}u!����h�����a��7]���-B��G��Y/z�H5L���\��0+�Z�q�1�w�0nis�ŐZgr�/LqI@�daA����=*Z���p�������b&��u�ZR6֥Gw�2�D1�7�T3��h;4,��*q4������"���B�f������ó�!0�/|h����AE~���[�/�Dj�����L0%�zj&�W7��*_�$?3�(���ЇD.W��3oe��W�$ֶ��Q��bT�6�	�CW�Vy��'S���(�)�/F�q�l�;�>��:�-`����ݤ}���Ӹ�O�{j��|���rZ�����Br�6G���ɓ�C����´z����$j��-%S��0�6^�E�iJtO�NzZ�=���P{ �\s��!m �DR�޶TJ<��uh)��o�Qv\�tH�Eo���SM�
�J=Me��k,�S6E힃��꧶����z|'pJ=	��H�R.�"��\�Č��.1�ŋڎ���빾��+;c��� 4P�}��_�ỡ��84k�ӕ��y�x`��#Iw�
��ש�"<�X%�̶0�MؐC��R�oq��f1�3�X3�N�pP�xw��r?Hq�T,/t���Z��-��,��}���<)x�W�%?R��'vfo�J��a��\8��o��9i���)�ܠ�����厠엘9|D��3���?�-�>�N`�L�g��@�x��LG4����f���<�����O�:��ܷ��u��
�o��L`��yw0�Ā��a��*�VO�2'�b���K�.�'1H��7�V�'��
�$��\j�G�\��}��a(��?tfڐ��lJ�E�ˊ��Hr��X�J)��~L��*�6���*���A���2~�/�[s���dO����V�R�OrQ�>5���n�����p����{�mGm�����0Q7obJ���e��SJ/�c�s��X�ͣ��}5[���Hd��d�v+2M��4���F�������ĕ�9�ֳ9�E���)����=��1T�u�ſ�����S��#!�»̊$v�]�5���n�rP�\
ZPԪv'`�����2�\�a��J�ˋ盌F c㈌9��v ���Y�p�&�����T��0��d�;�V��9�co}��a�����;���'Q*z ��<l���H��2H鱮"�v���g\ص~	#�mӠ"p% =���O�,-	s��H�+���#r�������Fv�0�.wN
�*���IM�f&�]�$}� ����K�+�}���;Ւ��ۑ��D�1��X�%nR�
��F:�4k&�V&o�2�I\�BL!c�Κ Ƽ"�$L�.|:G$r�q���hz!0u�XCqXQ���ކ�*o���;�ޥ�I#��!���=�O%���Z�Ɖ#��_�:��ݶ�C��7BA��X���{�T�|H;�D����O�[��y3:ɤ3yrͷ�m�Y����^WRRx⚑3�*��S������ j\A����6�r4��-�?vp���7&���6I�D��X�F��]���ɇv�m[K�����e����oG��(IN�8�`���\.c��ѷ�3{`�B��&�59�s�O1���Ŝ�B���O �	�
��k��k8�HhmUr���s��w
��������>B�|���G�m���f��W3%d����m�8���ؒ��9'�a� ������We�������ᝪ��R���c�);E��Y��i���d���V��P��
,J�P��H��R�b��������/C��W;F��|"ZH�OMJ%{�h���	��I\r�;!t�⫙ŗ����)�j��(Z��u:-����MQK|.��ݾ��MT����y�8��~����+;oǤ�� B�e�p��>�;��K>�C*��	�д��e}H�\�p
�̈E�*�6�	���$旵��Ο!`�9����홭�_z��L���9�'�#��L�-�%�.���˶]�1�/�:gxE�W�'��+V�1m亝6y��}IB:��]�Ɖ.2N���#����k�a�?�j�,�N����Mkp�����nDy�Q��A��֒o���$��g�PƼiƁz3K���Ƚ��P!�A1`6�0W��kaj�z�8�Oy|����m��3-�Ʈ�v~����(���g�ߐ=r��i���b��ev,mT�8Y,�Y?���#���H��(k��2�(
t�AQ���́M����o�eI���l��#�ܗ6�82�f�|���*=:"2��_��A�8ࠄ��l#����AF�uw��M�#~[Yg�������z��ã����?��x�Ϳ��W��W)��K`-�H�(=&����� �x>�ŵ�Y�]�:����]c��~;_e3� ��Ng�m\a�9J�?����/���)}��k��j���}�X�.Wԏ�=�0��m1�˛ ���q{s�NWJֻ��S��0N�ɉ��08�jk)�3��¨jů��x�а
x� k|���ˣ�-��u�ר(�����sc�s�~��ٽ����Ix���\��M����
���<��/�?��jE�0i-w+Sk�QK�e0W��)���t�bp��4�V� ��UG̷���(��W�
VV����l�1�.�o"��1��c�'�\g��{|[`����׽�+�<43����@�Q�wu�����]h+�A	>f��of^�.�e��G�J�N�Ʉ��PP�/m������l%�E��o�o���*_OϪ��T��B�|�x��,uj�h|����� i�i��w`�4��iDOQ"?��|̗%'`������ �3�z�f�S�֨�@x	řY_�
�2	�q�2���#4&�e�C>Yp����R��~�|��t1GY:�,1C�����֜�?!J){��*�Sh���#at�ғX�2s	�����G��Sy[�]404d������,t�S�7���������0��gI��D 5W�by~0pt�a�T�D���'���D��ob�-���A�*�
��,� ��t�n��C�������zP�9����S,�f��%�MQrT��.&B���ʵ�cK���^%�ΆZ�i��(R��W���^r[�CD�UX[^5�� �;n��)�F�r$d)��OG9<v�8��!`��]�,r�H��?����r�R9k�O��*���@�������7��>�_��e��ù�e�D����(ܒ~ú]�᠏aK�  ������A�v�j��vz�}<⅋��KP߼�k{T�Hw���:>L0�20�Ý6�&�gs�	�Q�"��	Jg\������~��ң�Mxk��CIx۸��g��*XA��I��i�c������V�o�,�ju�o���U���<' $���Uv�p��`3�����L0Z;�'�����э��&�#�av�z;�����YO�h���I�{����
�FzT�t���(��m��T�ܾ�94�J@a�ñ�H�wS�#�$�j��{�O���7X��d}�|qsU���e�C�C6~�e]���Q��x$Q�8��.�����q�[տ��!�zS�#����[J��u_}�|�ٔ�����Ǒ��}3�u��K,O��h�͆5�ٌ�ھ���/�4ҵ}�M����#~�=���At��}x}��VZ��;ll���l�������3�'ZfFA�o�("Fm���q�t���OG�KD2��pS���0U~�{�w�9=��7�"�&�g�lh ϲI�K.��*�T��*��9�g�Ր���JT��<gk�:a��a���N'Z��H;�mF�\d����S�ڞ����׭ۈ���lpO�N۱�>�1�=o̭�:�����ɝ_P�ڮ)�a�a�/��]�Fm�C�iC�f�YH�+-=�^9����(! U�Fs��+qC�k���Pu�/2�����M4�M�5.�V�SΌ 7����o�B�#���#,ꞙ��*\��L�F�i-��� ��� &�9��R+6�%6z�%�%Ez{b&EW�����й�Ra|Bab�!�2���sk�;���Zm���Ĳ�|H�{5�%�ei��ۨts��.R�t9�%D��g�Q�X�{�Yd���0T����fF>��+�x|�V�,{�Rl�v$8�  ��Y�*��T S"��Q��tO*�J������t����E�fY�DFGl�`��_��\�y���k�Rq��}K|r^8�c��U�m8��W �s����SOw$^ ��l*��vV4W1 ��J��Rm^D�ה�TM�H�'�ǔH�Q��DE�ڤ(��wHԭ�i��4�p��tȱ���e�7���I������\�s�n�&�©+����
Sύq��;�ߗ�6��xh`B��8�e�}e]�r߅wɆ[�]���q��8�#m���ـ�PvH�cEc��&��o�b�ڴ$f����;�5�h.�!АT���I���DN!���%�N�4�C�V3��F��k�K���g�{\ _}:�<H�/���2�����C&_?/G���j�N�'��f���p�Q݋�<$�/e��X�A�!<畖H|�X���z�1ܐJ��x ^�zL6�)�D l�Y�=<L�1��"@ӹ�7��0�;c� i.p�ld�޻�SԴ��EDn4!�P�±������L��Ϛt�_sյ�� ������\�{Y܁�u��8'Z$��MK;c�� j����A��iZ Q��lQ���T �3kg�#c��+]>4Nx4�v|�Um�m�-���o�Y5.d�D�b��w臤q��,7jO��J�(1�9ıHa9��� �!���l��Ӑ����0%o��"[�� ���Ww'nshx ~�;�z�&2��-MCaq�����'q�=�&Y�䆶D�����.� �b=&u��|����ZFw�o��İ͉Ĥ�����ğ��n�o4䗈��!�/����+9L��3�l~P��нB�G�w�c1籚|�d�}к�E�3�D�~d�ȷ#�����xzD&���~�5��;~(�¼�C$�C:8�uB��֜��l�T<~��	��^�u-����-װ��e0����1�㙞s��Y���vP|(� Aa����=~`�k�3ꋼ/#�cT��S�)gN�����vj�ba&zsLӯ�0���tU��Ո�K����ö+�O�e�.�A�F����VB�HTE�p~Ƭ��un����<������X(�ג���%��P���9�����u0����&x�\�+�O�#d"�A@��^~����s��<<4~�a��96R�������D���$}[\I���D
*��A��������`�7������~���O�1C+)�o�����z�4��fR��+ ���b�n6^����_P$S4>ջ�������İ�	�>mJeZ����7�3r���Ñ��>~b��d!�f�҉��4����$�I�"��@L����*k�S1	����P��J�����Vt.8K��	��CJYTW&�PVPF� �0�0 �����x�ʓ4%�3�4{�c#��<�NmԼ��B�����;�i1�=r `�%��e�	(K�#F�wZ��굗�!�x������oi;�w_Va���蹈��v�ݶO��xP2cu��^a��L^Y����tLH<00c��B�k���r$\o/���V3��B����5g�X�V�4�j	3'm(X����Ņllw\qg�>��V����F�+}��*�)R����	S+�*eT���f�)�)m��\(P+����}� ۑ���d�g
���iD�}�sC��
�㐻$Z�LC7�	�fy(���F.Wr�?>,1�:3��Y&7��dJ|93*I�t�q��͉��[Ѽq���{�plB��U�W�<�5�����t��o/UA���Q�[�J��D�|9m#l�����a�����H&a\d("�]v��P<it�9��=Hla13<k�~E�+)"�M�ّ� D]��L?��\��?}�B�q-�X��Y�Ʊ�ρ#�rX�D����D���~�T�бDL�`�z�&R� "�)Jh�<���\��&q�S�|�/~��
{��,[ߕ���WH��يr�� �<Q0��K#���y�q��DgLgG���ɏ��d1l�����snw=�>��%������F����au�3u?�����a@p9�f+��zS�HϪ{c���؆���ke����  o��*8�5̵Dwo��2N�Q�Zx��q�e��Y�����w��@t����qĩ3S�U~6�����DyF���eo��|�O���px%�j�sϖ�htJ���qUX;	�H���f�.{���(vf��I- 7SP�Y6����ݰ�=oS�����p�Ң�#낁�\�q�e������Sit(3*s����z�]��겳@�L���?�y冘����c�����z����e�X�\3��OeX-�Q��rx��X���b�ľwy+v���I�{)��8bI(S`S�� nl
!��Vǘ6b�u�f��m�#��q|fn@��.q�d�)Sd(�j`	�sLI�-	���#�TiD�b�*v���<���zs�W���)�4xዝ���[0�[6l5z���TG�����F��J��5��΢��s������1k�
�<�2V��ʛ��e�1x�K�Ƕ�2G��N(��BѓS�����m���h�ߛ�h1�}��!Z`	 ���Q��욆L6�S��e�o��Jsu0�O��ۇ�KSek Ā�P11.�=4{o��ӞԖۥ/L�/��.��@jN>�&X��0Sow#f�w�_��8�.��ϮP�za�f�	y`w�w�2�Hڦy=���gk�Q�uG���;��P�=a����f����ϙ>� ��ԲZ���:��������g��u)�����a���/a`#�(��U}ĥ�~W�B�$N؂O�SJh�=����/�R#�hd�t"�&��#|�D���:I�12f+��J�[3v�r'	���:�U�����N�R��*9�����*p��,�o��#vA��Y��9�l��S�a��aa�G�� �R��{�l8[�7�"%�3Y;�����Θ���L�	{	�6��$G�$Z'�����135`��cS����K2ws�E�'�W��]DFiru��J�F����((��dB�K��)��D:n��F2Ę����� u��N�^I;<�%�<�Ŵ"�}���ܘז� S#��8�5lKB`yhgEch���Wˡ,|�T������O3��[�J*�1���7�2�:���Mm6c8��P����m��XO')'�S?T_�B���'��R8��s�Rk���W=l��{�W^�\Һ��'�b�%�,�,��(�3�TQ^N3��(��0�H���<ɺ�f�g��k�&��z��T�5�	]��ϗIA��N�K��B1�D��"�Q�����:���y�{�=�fL�@a�w�N�@"UOxVc^�+��ӭ���>h���� i�WPm&${��7�̓}k�rCV^#�X�C��#�Z��C���W�(G�w�iT�!?��;�'�����C���|��)8=��ۆ�+p���xYl�s�gA�.���\��br�0I�܊A�3�`�?YY�X����>�iӐ���Ó	W�n��X�C�o	�3|�����;wAīB�l��mtj@XւZ�m� B�I�$W��c6
���4?^d\���V�"��֧J
��?Z������Lq.��>�M�^���d2�'��QDS�1�\���F��N#�����Ov�%<4�D��b'� ��[7�<1����%F�Wk:�7��j���_g�ԃ�x�D� ��b=�2�4sE�s�z�Q����;�./�'Q~���U<��=0`��!8wA��r����x��R4�����7y���g;(���!^�m�6}����$�N�g�_��	1~���*����k2Ԅ���ֻ��o��<�Jaq��B ��G��%?<�6�6��68�1���heF���i����V�C߶H��]�+$�1�i�'���4X�8�㔶E��l�	���=�����J]Agn���ϽE��K
~ٺm?O�[�����x�yʭ?��F��Q}�k/��A%W|i�{٪ɴu�����ce�]?1\��!�L�NZ��('�\��$�YeӸ-_��/�ul-�����I���	B$/�[�mD��vJ�|	U�U��ϸ��(A5�M�6%xFfyO�C��a
n����j1��y�۩�	��؂�0$m��q?6	�������j�m��wD�"�3'"V�]m���<�ߝ��@U*��E��vg�����>������V��8PAӳ4�:t��[![L�JP��L��yWw D��G����Cr	�s2Yo�
N4!�`�^�&�Ge
��	���>*F�|^}����r<y�l˯�AJ� =��"�U��8�:c��~W�+f\᷀Pįb>�:M65y�]_����4Py�U�!�T ޴Z�ՍޱW�~�8��?�x����G>�8��ΨU�ʫx<�R��wd?����hB�*���?I��V!�2wR�A��%�Q��Y揯��s������KcvD\߷�knq0��]���u���r�7n�܌�A7���@fik���wX�\İ\)��y25q_3�=N�J�� �X�t�$�d����UW�����2�&S<&����?�$n�}�x$$>[	�L8Gw�a`Tl�!^�E��ӶN)��
�5D�7��}'�Pv�� 855o<���Uҗ�G� ��8�,�}�O�%j�uxv�6$N�=��y�������j~ev�r��U[���!���1L�UܸV����|R�y�G��(k�����a���g��K�J�7�F�sI��$J~��u���Li%�\I��1m^�|v ���~��ļQ6z�V�s�sj�n=@��Q�p�g�|��X�~,���-��iV�t)9��QU�Q��ȷk�_�F��;�����n�(����ۃ^z13�!fve�5�t�|����z�k��T��L��vc�P�/���Q%e�#p8�:P��	��޴�p� o����6�G��l]�^��hw(�&Y:�M~��U��4�����Rk�ιm��J8\�р��	�eM��W�����q��ʟdK�ɠF�D:�V�'L�꿱w�����/vᤦ
��~/����4f���ĩs�r��dsh�F�J(�&���pE:=�*�xǼ�:�Wx�-?�w�Z9A��ŖS���*�\9V�,fk�
�V�H6����;��~��h�jɔ�{v��,m�X)�����o�;nt� �Z���X	F)��H{�QK.�cG05Jl<EJ$�bԩ7�/&+qY��Xi��,�oPej��*�m�����![B�L���y��~��P#W�L|�����1���+�-c(ι�~M�Wa�Z\��W�T��=u�g8|Q��跌���CW���7�J���p�@z
M�h'��-��Y�[���심�V��yy(��lT%\��[�tW���E�/�x&Ȗ8h�U�H�(����H���f���)J܄ ��$T��#�jj���0��V�8����dm��c���-Љ�)5jѼ��GM��7�|��`	�3T�3���Q*�'c�^��yw0���h�ū�������@����?W!�{�D�9����y�;��Y��Cǳݘ:�]<���åiޞ5�wp^>��p�xEK��&3�Զ.4!�H��"h2�'ܨ@p��l����jc�"�n|ń��`]v\�����-o����8K�����})}�������[�� �`ţI8}�੣N�8�{@ +e$��� &\D'���:�XȺ?0�~�O�g&��-B�sy^zlo܌,��l�Z�cP������X��5�!2�':	��*:q?���ںJ�p��i0=���"���3��$�kR�3~��'O���Qc�*OE-s7��_G
:�^j!���r$���U)	P�4��S�Q�=��i%�������eи~_���3�e�t&q��u�J�}gt���-�!��Z���K	x���Y�D:ܱ�G�&�2f�I�j��N�r��@�s+��-݆��es�Qs�A;���O���Ȳ3��qQ�����9?=6\���j�m�Hծ7�s�&Z6�]Os��1d�
���%z
M���A�"��9V��ƭɻO{�P�`r����T(K�z+��"�/p�qCĕZ'g'�|*a�w8���l{������r�	�`(�������i��C�l�t�����|� �V��@U�@؍�&����t�3?��YW��ICh֙�qp��Ѡ�dYe�χvj���
-�EQ�h8��B\�.����^�&E�����u�;kx�#�������~{�B�nCK�A/��Z�B˸N@���e%���?^��:k����#��tY�n��_�"���k�O��=0�t�!�+��]#�[��[쬒UsuQ%�0'Q/{�ܯh�B��c=�:�� ���b�����o@��*ba��i��H�cQ�;�9C^��e�e�:H�}�Y���Fu.i?��԰�%��(�;�h���V7ٵA�
tq�A���e�'#}ax�E����WO�X�k�q ��v"�lP����S��(B�X���w�O�n�&�4�4�W�˔���B�鼢]����t���>�)������,�)�2.3�^�%{{]J�ǃ���	{��oZ)�n���1x�t03�#];��A����������صد�=���0��{)�/�Dŗg_2{0^%�Y��J�K�A��j.���.���+4٢\�c�<P��^9k�T6M=���S�}����ŉ��?߹B���"��7��#��X�{P�l[CE?����[���OMZ;V�Nx��eĠleb~��sl.dA�auR���
i�o$���"�b������`ü��z����igk0�b8(��z7$}�n$�G�gnX�/�f�^�\��]�o	Ӵ�R�'u�حuY���b��F��N\@�l6h.O�@�#n`7NT�hVk`�Q��X �2 ��d�&�ca�K�Yw� vM?�s8uu�+õ�0��Nt����r��3����G.�!�{1�Çg��
��qo���m�k�wd�#1ڽ������w`x<�'���išk��0,�Í/�gF��x�%	�g�Jg���f��U�\_ �4�4�vjt�k2�	��HL���@�+�N��_�*�ʌ�>���a�5��*�2�hN �F��t�jq�3t~|>c�&bY[�1f�T(�U5��\fNQ=|���\5�c$�=���㑳��4$�R�9����To䦨��q���>��9�6�6��"�x�Cќ�� ��NASh&��qA�7�����vW�\)h@O����8���1�7��w��!U�V�M?n0r"�>�ȺgN��V�Q�X����~ kQH��,��8u�=Rӳ%����C��TDtZW�:,?ж��7ƠJOa=Q+F�y�hX՟���HG8�WS�[%6�~���:��9pw��h:��-�U�/&�ΐ}wӴ��?9f��,ɴ��Q�p}u��o��x���e�-(g��c��,7 0��������SZꡲ����|D�*A�� ���ϦC��c�y���RanI�U�ǥͥ�$n�G��uލ�m�H!E�^WD�._s�Ο��'�Q?��j8+�.-�w	#"&��x�Ʀ�W�0p����2)�o�6�e��;�Y����R�",�Z� �Yv��b����gdo�rk�n�g�hT���	>5��[p
��~ߢa�~v��r�o�`R�[u{E��:%��m+�0��tq��I}�앐;��.�zc%���p�M���(�g�g<I\�XM������bxS�b��"�eP����E=|���}s��ˠ���:1��g�$����[���� �;'�_-��"�tb�����g�4�f�"_��*�dtY2
���5-W)��xz�*o"W�yW��*�f�nz����|`eV����#5��5�G�0�=ZA^� ��fv�2}U̪��4<ۀ�cӡ�w�7x�ˌ�-S��e�zs���B;���x�m��v;r���t;�I��N�LX��=�����+��v�;�`�quNT&�#�6���V�W�f�x�Np���#Ee���9��?=\;v�,�X�[�-\�a�%�����2$تA�jf	��߳��8�H5�G{}�����p[E���aD.�����NboU+3��)��|̿Pdm�x�ސ�єϕ�+K�W��΍^������k:���u�̊�V�@�{��榓O���������ഒ.P^��U(����2��I?gۢx�]��  	2_�#����2M��)���纱��Q׀⏂��
J	qc�X�{��g��gZg,!�=a�waHL�Ƙ@�_��%���b�d��'Zֆ�-[BU^�i��6E�%�`�
���5k����')\>��/���=����n��	�5�:4����C��&�!.CI��˺�Gv�T.S�~��F�Ƴ��U��u���SU��-/"���v?��P����f"��C �(�ƃ%�H�?� �Fļ��o���|J���$�ej���㔪�V4T|qJ�fV���������MD'#��g�ӿ��%ַ.M�H�8H�ʭh�87	�A5��(P���ȇ��!��I<0�J�?/	���aBBJX�- ���Bn��J���n[�oP��L$����O+�k<۔j労��ݼ�Ɍ�j�ZY�i��	��^P�}j)'q��k�!1+�7,O��9�B҅,p�6��_	/{��f�O��V�0�=Gt$�;�6��� �cq����T�'��#`��*NQ�A�+l\�&[ �1�m��=��Ir)u�\����6�"+7�c��<B�x^�_�p���x-�3N�X8UFO5G�N(_?�M�ޑ/lfJjTT��\ȯt���zTi�f�={ ����ǉ��X;-��n�a��.��*Q�1��`�F��G�T��݀��8��8���f�_���� P.�H��O���tk!F�7�	����U�����:ǯ�:�7v[��$i������{$�����_!�i�1�iPཤ�Jemێ�P�V�Ehv��խ2|�������8���N�w�1|�?��t�a9D1ˡ]�L�lE�ǽ|��Qt���L��G;g��0c�f�=��]�HG'$F�S	�q ����q�ٶ�ǨbW��w~{���1���� i�j��%��y��E�W$�q�ܪ�?���h﮿+,��k�����2��D��z d!t�-�V�D@X����^w����oa�-m��`$*�7�����	`B+Pѡ�d J�m4�>�U�f��u���.�{9��=`�پ!{hZ�n�R,=��y!�nأ�5۹Ε`PQF���(�4��X�O��W�4xZ��C*�0r��r�;!��>�n-��cά�2�wֆ�	
چ��\p���q�^ӹ)(�4i�����-ʋ�s��Ħ�?Ggr����!�U?Pq���rY͍���A����ɔ�4��RS�'�S˰�UR|�R�u~P�%�u��Z*<K����l��o4�Qg:�n�-�2�$�t�A����1��&�����ނ�1]����-A9�*���J�sL8h=vZjy��7�g�]��)��4u(��є��A��q���(���?*s�^�z�S�Ɉ�c"tT.��yo^�$"��xn�EI�Ҷ�2=��wT��{�r�d�f�G'�D���� $Y�%%D�zJjZ۰7�X�<���+�����vw�A�z�ؚ��8H�ЭT�ȷ�*� ����,�Wb��M�(��� ���a�����ir4b=K���n�H_���LE3�#-�ncQ�g���W
����/��Ѐa����$�-�,E4w5&N~C	F�Ӱ�1�+�.r���v�~�v��"L*v��ހ���`�W1:ؙ�ؘ�.��w�'f���ةk ����3+����$�n��^S�� -����u��"lZ�'/���y5�S��m T��#�`�BG�Vm#�5�jse�������3

Ә��/n���S$9)��yS@:�e�����㼳q}gʉ�D����u�F�Prg��U�����Ӫ������(�
���I�)L-<-�d�$��f_N�g���R�&n��x�k3���)�Y�#}>�*x9��m�~�\8�ƻ�d�����V"�#���S��b,��7}���b��d|
�s��m�X3u����zkz�=���<C4�C8��H��]^�>�$[Ŋz6d翧�j/[�F!���p)�>$��;���__,[/���"�X63R��A0���1c|)#��H8Q�.Gw�g��%��\�d�p�+F�<��� nX���E�.Z�N���% ��u5����X@a
R�,aU��`��X�:�ۺ��,6��%U�+1�v���d<˺�ѯf�d�B��o��ʜ]X���o�� �S�<��Ј�M���b!Z�P�k=$.�$d�)8��X���K���(7��[�UY�
6�kT���jise!
������=4�4�<����1Mז�;� 5�E!�)!Mx/�{���p̓yz�ۭd^�/��5���M1$��=��\��oi�>�|S~���}�M���A���S��sԣЌ�,����F��(�ˣ�V�6�ʱ�w�	���o)�Z��,��v����<��������DbI8�V���ɨ�"Cվ�Om|a�h��l�b�0[6��;�Q^<W#�5�=�*֯���aH�bz�'�
�3�7 [�Y�������7^a��IS೟8��v5	�&�]��T�����w�[�,��p ZIp��� �c�\5�~,��G$���I����
7!)S�a���bU�j cz�:ˉ��67��j̧פ�ֹ��h8�y�za������#��
�j/���ԣ.4�r=.>�>!p����{Cy�g��B�۳\Xc�e�#^"{��ϳ���c���6���ʡ���ߠ,e5ƌ����t9�bWFrǛ���g�ԃ�I(`/��������9#�� ��V	W Hl���CR��p{�9�V�
�A�9u�7�U��{l,VY��'\Ԟt<!�r���tFDY����i�$o,
�.z�Swy+��je�Mfi�����k��m��u��ۀq[��Lh������'��A�73%��<�i��9�A�M%��d4:H�X�Q`n�.�=���z|uR�V�.*���v�쭛jwТ�C񥆳�N~��.^f��Aj�n_/C��o�	+�K'pz �����2�5Î��y�M�P���TͽVb<3�K�r �6k��W?��c\��?��g�?��Ю��O��k�8���M����ÌJ�z���HQ�yo�	�;J��cJ{<����vd�T |���BLe�7��$ԣ�p�m��Sf��B�g5UI=
���������5D
gf�s�'o޲�1锻�*T��	��T���(��EmWR�h��;XP����!�d��ly�����]My(�j�~�ݳ���k�T�7�^h��)�p�m�3�ͪ�WE!qY��П���M�M�CIfP�����K&1r�u��Q��t}�
Y�z��D��v A�8��A������D䖻-��˟2Ԅ+�ֿ1A��>�m��̤��R?�%&oS��K����Q23�7sБ��ϊf���3<����p�V��
:����T՘o����9��@3D���?�����O;e>��ƾv~���R�["���ə7w�f/<�uB�L��#��z��������6|>���u��U���7~!�����p3�HXl�/h}��t��z?1��η��8K�J;c��V�p���)� �����Z,�?rb2M۶�:�n 5)G_O����%B�W���F��%�>���Ɍ�D�9���
�Pl�.���0�B���3G�A�u�I!`��P���ڿ��\luؒ�+ٵZ�c
�j�����,>�!1-�Ʒdn�j���߉A�����^5��|Z��L�-��.����(υ��cHm�03y��[������Ӽ5��5ݛ�g�%ktZ=�m��2��[�t(�% �^���us�(%�N�<���>P�f�S��Γ�Û)�����La��Ke�z��hx���+�6K����&�5ӽ�VJ)hS���w2UH)���F�a��W�/�p�
M�Y�[����J�M^<�}�<)/��5sۙ�`�m�I����β��# �����n��kI�/L<���� �	���;.�@�"�c���i��0��:�j[~����)�f��
��-����/وgT\�����(���»j�nS��v�������]��%�����E=
Z'l!���C}!�4� :��qaG�}#is�y�_�&�����>;�X��k��Y14�N�Eg��t5�領�T
�o�z�`~п�Z��Y���5��*jE_r=i~�|�f��y���7�q������ vߩ����NJ�=�S���E��J{�^DjzHQ�N�d\��A�d�'�N]3�(SH���0�]^_�O��+�8���^��L�Ф���TE���M����2ft�uV:���`�&�� ���"�7� ���>mi�l<hQ7� �P=fe��BP���鼳�Qbѡ���*��.	e��=�j X����`r@K�KQe/�Q��/�X"M[ƴ�;>��������Q�6�?ɚ��=�ɘ�����w�zK�4�^�ΪU�@f�\҅�~��M�v
��6Y�u�v�r'��5��W,����[Tu��2_c.?m��'��~��/��C��-7�~�A��V1R��w�SE���{��5�$G���fP�ܜ�t��A/��sqOG�tY�%�ke;*���u�
��<`m;M/����o��<7�� ���@ĥjĴ;������jV�W��a��(P:Z^�x��.��s3�~��I��ĕ(��e��p�`j:��mR���/,��U=�����e����Q��-l�Nj��X�cAZ9�ߟt�N������Mw�f�\ϖ�3������rt����>�~���Hc?7�9Yκǥ��a�Pj�Z��]������`vƕ;�;#+g�^���=YB��B�]��w��Wu+��Q��틣4!�Z��� M
���B᾿���%����_�Š�d��P$d��`�(�������|9ׂ��|ڢ�D�W�?��*4�j}qէ��.�T�D�KDÚ]'�?�|�*>=����7`�êj�|�!6
5� :ΓA=Wvw�L �n+�� Ď+�>׷�]���֩v6������%�`�����ߊ���R�:�����ޝ�>v"jp6��CA��}�|;.�g&�u��v]0a.`�� U��%Q�qm]y��ޠ��X�Ny�Ɔh.�{g��$������������Og�^(v�������~�k��Lˀ�ߖ֊&�{�aHx����6��f�>M���
\�_�5i�C��Kr����yy5GoeV��,5/N�"�q�'�"{9]�Fj�n�'[��k��a�O�viD|�^�`LOc��P=EsE�1�*�t�Xu�ޣ�t {���pN�v�6-�=��˃SU����-���%��\H�7ƕ-����..rQ=
��?'g�9�To�е�R	�F�>�!�Rp��.�+�4K�p�� �'�V��Y2��1��U�
� >]<��[�t�$�LEO��4Y������a��d�e|+b���t���6��8�KCz��uL�����s�˻߬-�˕�az�8�7�o����RϚ�;��������qb�6< �@4Q�7��#^#Z����S F���+?V�b�a?�	kP���,�ήWS��X_�uP�'|�*��Q�2�C͌��6^��-��0G�i3>���B��ʷs��{y
e�q4�(�u���
-y��XB1Gw�mi����pr��3�Y�2��/�,ϕ}/���Ɔ|�l��5"|��/	��Q2bN����Q�_�,I�yj�i�א�.R?���"��C�b,��\�1�uWZ�\✆1�'��ЫE���|�(� Q���@�v��#XJ_G������5����?�#l����˦ݺ�~�^��hYAe@eER*u��؇��&Q�,m���v˩�nmI�b��@��F�T�)={2*d={�4�#��i�O��凪܈��,X�r�ћQ&��LdFQ��o������~$7>px��A�t���ē��'����m�N�4�{�M�l`Egr	�AÅ�P�
���©q�������9���1�Ю+7�}sd�j�֡aQ�����^zo�;O��x��6����@Q�� ����5�`}����E��/-Y��>kKA7�PY9	\����1��m���7J�ko͈)(������E�|�Z�����b�t!��ܪWb.��T�O �U̍����|�@�S�;�b>�O�0�������(�'n��#qBo,
����p����ƪ�}8)̂6O�hE|!5I�M9އj�'Jqآ��O_x�)��p�����7`�C�?��^
��zGރ�2���f�?ls."<�8K{��n$c�o�m���*���\6�^o�G�ɲN��=+ǎV�BV6Y��ϩ�d8��x�r��d�QK��6s��� �4���v�8LܿNBO�� 1�޸�m�u���4)F�فU������'_.1�%xK��V�2���Z���?�O<�:T.GSN��g�?sW�������K��8)w�� 
���k�S1�@<J=��.9�+��c�Qg��v��2hѹ�Qsj:�ms�6ы��1�Tc�Ex�'�f�wp�G�o"ɞ���g��J�f	��m��4o���s�B5>̍���ȓ��`�'�4y����t�ZӧLr���_%}���h��n��,TL�1Z���7�Tɇ�n
6���c���c��Ns2�ёo�0����'�� ��_M�<�u��k�qN��;ֵ9�W����ADu�@/��L�`�ͤ��Iϭ�}��,����n���LN�1�>�=t�OF,F�iKѡo�*q�5��KӤ��	'���15���*��n�d$��V:G��n]P�Y�����I�m^2b�5��	���R��
����5l���w|+q0�����ƙ�X��'Lo�Q�b���>���_=���*k`i��Y.Ity�40�Ald#�^��V�C�g�GF�2E��'zF���P��0�P�����g��@�4=r\���/�S�$�~�{V(�oK��$`yp2�����-Y评@6�9��f�p Y�6w���@��b�k53��߰�2���,�[hN���	ԁ��1B�)�Ÿ7�"���t���C�Q#{�d�yd�0�����?cZIМo�j�F�P#7z&�_��q����[��3?Sn����H�-��q�ߙ���\v>�A
�/7)$���Q��>`]�ˀ�o.?mŮ���}>���3Ф兕
�&�)p��A���*�E�����6yyv\O�n�vx�r\	0Z���5�������D#��>U}��0�A�T,�O�e��[�����e\���������O`�l�1�$��	�uE^^����PШp��uVf��M =,�B4ʓ_%֛SC��=�inr��PWׁZ����k߲8J�����.�5���kT}�J[�b=��n���3?7�N>m#� (�vّԫL���`��屚��S�[�xP�w��V�����o�) QrVP��	T�	C��r������=E�2�L�7��;;gH����z6����_۲@8;���W�C��r�����r}��%J���^���*J������*&�>^~5�Lٸ����4	=D���{J"7!F|��>��K3B�����+�)'�n�m�{�Ɍ5WwK|4i�%��'������)D�����0����Qhm}۽Z��<��1�4�Y �)~Ϗ�dqH��M9�N�RA�n�O_&�m��Oy!�x���(��v��_7{���cY�e�&\���xj���B�k9�&���0BQ0�x�����Ƚ��^.���$
��s�7u�2C��Hک�A�+��1��e�(VF
�9��>z�}�́n�ܰ��O���?�Iх�h����	���@Z̿����x��/Z�\�U�Q��q����}z�S���Ƅ˧��Kc�$Gu4Q��t��ͺ�x���٤�2�ˬ2�� �hz6�{�H0��k����������8�?�Ք
�7%�qӔ�`_���!1�g�s�WB��pf��q�E�Yǹ ���ڃ��[�jp��=5�C�FH�b�����2ށ7�΂UH8��=���y�����؁j��<W�q<���@oZvN@O`@,Y�4ohc��!>{�墢y��|Y�T oe0�#L�C�:��7z3B9�~�z`�x�mk��Nk�z�������\�=��z��#Xj[�VK����̈`G��+��}�Y�����t����8�j��T�V��n���&��3gĹ�SB2WAτ�Vl�^@h�9}�!}�πa������ipt�b�F���몄�O�P�y	2�
7x���)N�}�]Vρ�����9o$+q�������Bft�o�s�r�4�yV�[!ݐ��6I$�FTb5�|~�?�����?mĨ�h@k�$��k�L�9��t�񿕓f ��L�3K$OߘqT��Lu*w�4��w�LdoOdT����Y,sm�3�g܊�.B$�-�_v� T5�H[
���G.l�6�S��4|I�I�G�S���~B���\ĽW0o���b����<����-w��\�1,C���t�f��pWA�cHP��GC�:W�8P��c�#�`0!��=GM˙(��5HC��Cm�^�_�l/jx�eő�G� �"��1�9 6��ú�#��Qo���+���,r����P�x��n��SËF�f#p���v�kL��meOQ1E��8�6�[����:UA˸=(-V.s^�|���-;��ʏ��b��<���?0���c>�^����||���/����o\�_Q��Y���ux>d��UQF%pj_�]HքX� Lg�b����Z�����f�B��m�B������)b|ג��7Wg
,��Z�yv�q�;Jm�H�/@�H+O��Kg�V��TLD{�@�FF�$I�'h��G:�]>��)����'|�S�1�#���(�G%<ч����਼ޏ�=8�GG���V,��{�=c���m�����8Ḟ�Ú3ù�������<@$ځ䠹�^��a �9X�z�:�^�0Aa RS�����T�˔����L�R���d�7ߩʨ�G�������s6�b�Vdu�ޞ7M��k�hK�}s���J�I��xP35�+H��C�@Lo�����t��M�4&���޲i��a�>/�U<�xXR���I���� _�FWtd[\���pl���`���[�_�C������R��g�=�3�v¤����Q|= V�j�Ň����":�ǈ0�,A�)o��=O��AA�D���UX�	i���)�5�B�FA 4A�b���N�V\��YB��,sp+�
���ถ�-�F���Iͣ]N���l��H�=�ւ�`��f�*@]Y[�C�6*yk}�SJ��;��?�s�T�u'|j:����Q�Q�]j��@���kW���
���c��7O�u6�p��٩-�H��(P+����ν��ް��F�'���y�F�p�E�h�^�ԕ{y2O3���1 �/��.���ޘ�~���*�@$A��Y���ȗZ���.�~�-���M`D��`�H�f;�3����r��NȾ�f���D)���]����Ͳ�q�b�ƶp��z|����)��_��l1f�
$�37��v��]��m,��rZy��G��u�	���d�k�!�6���N��'t��B��-z����3}������Z������x�c���L�;�mÞ@[�%l�eᜫ�g�!����f&7}}�`lzetU�ր�ώ05O�u��fh�4�|�7�Z�?�Ѫ5�G�V�-p���ϜcZ�1��3M�O�DY�v@�9^��7=r^��E���;�6W�=\=�#��������bD�U��\�%��W��\Q@��`F;�*f��T�[��\m~L`�f2a�$�Wq}e�UEߒ�C�;3� :;��9�m�k�Z����������m�y˞�(r�&�_�y~������&j��-�O�IY��F�0��)�W�vۂ?��CR��`���K=�?^{��6_�ur;j����>S>9~�$(>�C��fkF���I�݇��6�F�>�� Ɨk������mh�Ł�5����݅��:�,>�����=Ŏגu?�K��\�#�s�B5�����{���#>C�=�a��T��z�� �ģ�3�8y�.D\�BV��E��OJ�"�6���-�C�>��ه��|m���j���|�%z����z\-;T�(��Ԡe�|��E{=Ɂi3�����7]Sշ޻�a�X��2Z+��^q?I�[���_5<l��wi�6n���7��͗�G��+��/X���ꍧ,�l�=��4�T��{�;�#x�=E���w8@�Q�NH��=�m��EH�Ӯ����OĒ��/a��g��1��;\��Y�PSn��LK0�ۂ?k�?�'��Iz��!�U�g����`$����˒�gz@;�I�Fk���ؘ{�+��R�jg*��c�1f.�,�Y�[`����K���,D�ҝ�q�!S�w埇J����9��+��cK�=$�+��N�D�q�8��C��ON�4*Rv�P`K�(�KC��a�?�h��G��*�Z��u�u��A�}�=WӓS��$�B[�������%r�@M(v�<A��w4,;3��W�-&�JTk�����5\p��$vAL���B<J,�wAW<c��_�_M(���!��8��"@�X�>��Jn�\���[�e=N�T����W��a����h�/�	=~bG���. G�#�?Zd��zG�j�D�&E��Ӭ� �^�����fi��Sz��	���)��񕩀�ۑF�����y{z� �8Qe�q�r���\�p<���Y��H�a�	X�
�y�����~��=-"�BrLX�|%������&���+�*X=�c�s�ޕ����+A�[��9�R������Z"}��5S�2�v��b"��~�+���-�,I�m���E�hc��R�?% ��n��_X�r���`hb����)Ĺ廞pE���[73|��"�l\�Ƃ��6�h
��y!�*AG#r�1�G�I`s?+q�VMlG��b�E]�Pd,o�=����E��U�2�:;(=���������o����%i0�ϡO�[C��p��8��!�z$����(���K�-��U�����L�(W5m�(�?�gM���Z؆Tu! h�����&�gI��	>9^Ǝ�1f�<��~$��A#B����9�L�4A���w9����N���w2��Ay�Jְdcg�ü����61�%�+��U@(�TP�RP��,��*��DI�����\�`#�F���� �g����z(Ε���A�~�9o̘�(��*uh�=�<��HͿ�>x�X�9�1URԚ0PI���z�f�ÃK��������d��7;zu+�K�d�7öJ���b<yf�Hf��]P4�G����?������em�3���f���}q�y	�2��_�vI��gO��aY�QWpR�Ya־��FhY���R�~�\�eg�`e��5�sa��B8���r�B8z�qN:(/�.�x�UT��tq�¼j/�eZ�z��r�GWQ���g�@:fRL��;��)B��5�[�K5A%-v������ �۪AC��o}��/���s$zЫ�ŷ�L_��EvG�pZ��,R@�ƪ =\F"�����W~�C1�l�|��xt{L-	(���ؖ4ӏK2�qU�z
 �7��b���ׇ?�s{��$���&�{��F��� -\���bB5�#�s�����[K[����{�[�ɭ����L�'H�޵�}q4.�WJCmIF7�<�4�"�K��u<����E�g�c]v��d�H>b���=#{F�8��Ծ�-}*�dJ)Ա.o4t�ԭ��D�U�sq+F'��L��^ߚ{�.�f�Ic�wB�9q
�l."A�9���-�g�AX���؂�C�9��R�|�3���ҵ¥;^ᮛjA��]�m��o"-����T����j����f����#Q"@:�C��],�	������ߐ-g�񝻫QCD�2U�w~�N^�w���y)��F��8B�B�����5��i}H�k_I>ۓD�@\��z���¶�ף�g�Jz�+O8���#���~][
�xY~��~���9靌�����:&�S��8Zߤ��ʂk����� �oL�#Q��V��298*]���1����u`ցO, �˚�̱�ur���>�~����̪6��8�;���!�{���%�� 7�v7 �� P�gz���-�Nӧ�k��vSV��J�.�siȏ����R��ACn�Gˏ�Y�y�Y
~�3����k?I��<�N?�E	M���#�$W�dxd�����Q��͊@�t���K����'6n�Y�ϩw�)���D���ni_��	n�vy=���8 �ȣ����l�#�ʏ�\Wв)5FП������O�e|R r
�B��'n�1�0�1V'���/�4Ɣԯ*���������l+ 8V��*�C��]H9S����R��Bb[�7�w��r��9������"�l��-�h�.�� K"s�Mr�)�� ڝ��Ş+�­�b<C�涰��M۷�_�9Wy�}��^���$�lJnRH�_�t{^ ��ϭ�˒�S����(^^�~"{��g����9�!���U/�x�.a�KX)bw����Tb��x��9�ĳv[<�UfK�\�q`]xob8EF4�X�����I�{?F|��'��\r���2D��ʮ��2�u�'��}��`�b�V�Ϙq�<���ո�u&H���/��=����9��!&�pGP�� ��r����) !1�PC�.LK)�<�v�W$b&ٟ�)c������z��ܘ�ԋ��B���Nw����-Ο��S%�L��n�2}F�B7u���ӱզ�҉�6��S��d��D�8�� �rwd��"�&�����A����l�fTȬ̫8���uR���!����;����W|�󃮿��fy s��#��C�}�ނ|��mV�3\�:�b��1\;@]�:�n��K��&-q�m�Dr�$�=���@;o�K�f�J}+�d��Lu|�k(W�<���ݡQ�aLQMp
��v���B�wX���L�IG�K!���e5O[S,
Y$Ea��y5:���< vHA��y)�^�Ʊe�Q�z�z�J� ����L��ׇF��ϊ���_�4����g�d-��p���~�@���X�3��l��E0�އ�1#���*�px�6q2��	�u}�u�0v��?�V�9^{�ǑB�-�U2['��p�Ϯ2Ĩ�@����_tުK�� R�}��FTvEJnQ�}�3�E���M�En�*�$��x��s>w�/�"�k��xǭ=7.�ߢ�]��z$q�����L�R,��;�u2���{�m!o�s���1H5fX�Ȕ*c�%���%��}&�u�􅌷5Wg\��7@�G4B�a.�Up����������e[l[|93 K�Q�;	��J�}���PQI�����H�^�c��f_�cj#���=�*@�N��=3��
@�l��R`���/箈�+j{ob�o&N��o�V"�>�~
�"�7=����MìE��Ш�y����D��]�!'&-��j�jT�-�	�S��������1	��m�~�����<�ɤ9��:$�7@�3�:h/����B&	�i!&͉4��z'B$�"��[��؅��,�?���n!�����ۈj�g��d�4h�p���[l�s:K�@d@�/�Mv�&��R*ޚ�K�]�u�p��n��#C3p���F��8{���s&c�{L�q��R���cu�� YH)J�����Ŀ��f��G4�3?��Y<��|�P�B��tגi��%MLI�|�-��k�y���?����I����%���Rv]�|��d��y^~��I��D�X�y���l���h!'��X���;�mDј����"]�*�8'p�l��M�%�>���-��f\]�)��1��=� >	�4qq�D\.&�����$���NdKF-7	-x�8���Tl���W��Vsа���3�maGf@zi���h�Jk�Z_��� htq�6���3S���9�g�Y���\��̿`,�?��mo�rǗ(��6�#�w�ġ��iF6�9:��iF�D����5M�f�/a�bJ���mU�2���5�q2�L����h�X�y���:�l5(>�����?�4��F�e��E�S?�cg��ܷ,�Tϑ��|�/ܐ����Ow�����%"�]ϙ��8#O�Bފ/�H�]�q��\k~����2׈qP����e�f���ͥ�>@i8����{|�w��u�����Oo� ׏���xE�����?�զ�r~k���`��?`���̀�ы��f[�M�ڔ/��7D���&0��GI��_J�^U�:��Nc�[ț�]v�k�#��e������)CA�F�������0���_��T�	�)�7D05��U��c��@Ù5�� !�[o!�����3XC�'1�<�;z�9���eIV�c�)����l�f�	��X]�-j,�3@�~�����H��Z�H0�z[}�(��%��-����1��c�Zv�ɮ6���1�m|��z�Xa�X�/1��}���3��D ��`gk����Ԉ�Ϲ!�-�cP����4��x���"� 6.�n=��3d/������F��@ڇ?n�?_�yq�~i�he�1�}$�<�D'�z�n�K�z屣vRڻ��w�ll��So��X���y2V�2�
�е�>�0��Z"�L[�j緹P�:�6G��}M��2��#�8�����"���&����ڔk���ƙ�W�>|+�8�X#�c�wO0��2�%:G`P8��g��,f���aU~)ާ�gC�y*���A�M��`�<��yV�ky���1*�Ka�G����O���϶l8��.'\-�(b9.�7/�&��7\�%�:y��8��S�Ný�-���d�K��X����O�ʞ�SR�V�KD"�N�f-r�)����s�C�Uf[)�����v�2�K,| h\Y�z�i4�mt��
�y!�������GX^�>05�cO�\�A�*�	�r�"�"�o^7�M)�)3����&�L;3omT�k���[���<���<�F!��kөGeTAT;C��78�l�V���6�J�%�:�c�6�Ki˙�sy��x,״S�}���ڽP����,�w��A�f�=�J�(��Va=������+�ۀ=�����>Ӽ��hv�_h'"i$]�^��}�i�i����}������d��/}G�����,\�e�v�)�}|��/��p�V�/��)�i~W&�H�G�w=1���8�L���Zr]_f�_�ۇdNgu +������X�9"��<������#������,��R����zr{k����f�~�޹0��y�N�49����\������x�p��<.�S�fvՅ�ׂ�qh#T8�B�oN�ɾ���S��gb�ힿ`�&�< F��W����[+�N��]3Ò�`�WG� �^s���!k�?�'��,=8{3�(����5�ͅ"Z%1�����
&���W7:Xn�Y�͖i=��B��������ȿ�]R�޿g?E�hE�)'���H,�q~��Sp�V.Y�%� �],�ͽ��p��6��۸���E�jrx`��f`���.��_Y*�v_�yX�`�XyA}?��ڌ'�7!]�9zM�P┹zRl�v�c���"�T�0� 0zz��c�c�h)����kDYJ`/N������\٩ׁͺ�H'r��m�^"��S$����#F9�`��h�Y�x��B`��y�I��E�i�w���|n�U�-ۆ�$������\�Ӯ�4�۲8�+��?�`
v�����<����g������dQ���[t;m�$��h�4�:/���L�ηj0��ᣩ�G���&[y��$���C86� �`��0�J�~���{E �d��9?�Y�:�4p_C���.��n��4���-�]�F�u�K�)�T�%Eȑ�*���E�BO���_AO�Jg5򁰌�Llut��Lò�R�s;K�RvwwI�!{���+�\NWF
2���o8�Y�xVgA�-|J�sӉDEK��Jd���ę$| ���$X/�B]#����=��x\�l=ƭm���o n��(��M�}*��fh ��&\�*��9z�Z��Y�L�0տ�{�v��;�����OlBf%���K��`0N�@''��'Bu�-�5�&%�ƛL�v�1W�D�w3����rJ���#��P���ǫ�H�η3���)���p�˦^���<)��I��H�S�r� ��:�Kl��\�lL�i�|폚]t��M:p?چb�o���'�C
~�ؕ/O�������}�D��9������l�&CJ�%ę�/�}�E��y<�A@E�9�}#"�a)�����Y��~��(�}%-�֥�o>�sOj�0�����I����m��.�I�y'�,_J�U�F�~����؈���o�
,��SG.�alKp��	���.�C�J�
ѐI}"��<���I��[=�NlK���mH��nL�!%Mg��n\�m�*��]���10��bٺ�>�g�e�I?���x��rh���tF�y���$�іB���'6}Ʃ@�/Ob��3D�b��, ��%��SE�r	�(��)���r~�pG@��h��@\^nqcp��p��!]�/��#[�y��bD>h�q��_��EihP��/��y+��M�G���������l�wJF�i�I��[S����X��J�i�UTI�k�e�i�ǟ�Dw���E��+���4�f�:I��$6<W��f��;������PI��C��y6'v��a~\(	����ov��J顴a�|����Xa0��͍8+�Qv��i�#�Id�ЀaC)�~�Y���	f���6k�*U�Gm1�O�.�#���%1�"��>�{������RO�s�6�	6���X: N�!A)������瘏5{�i,�ź��E���MS�� ƻ�Z��o��Z��|�XF���!!�2vx���Hqup�X�*�	A.q�C��d۟�-c���k`������̦
��������{���'�+�Rm��ʕ��e����J�ہ�)Q9kp!(Q�����R+�<'�T`ΚE/Z��jp��3q�t+1n���a)�a%��,󠏬��R����f=�*���G�s��3�����|��0�W�jQ��p'ʄ��g���T���[ʗ݃����1��QX����9u���qI�<�8Qh	��=�>����G̻��t�!����ȑŀƧ�9��F�b�\��ɠ�*���l�-~8���~�/��~O��q�&G,;�C�[�%�xU����ם}p8���&]���Ii��ņ��� s�]4�����TS��Ρ6��!)`�$�EA�t8���;��վҩ�N�e�"��M�~6�aAś7�'{sJ	Y O'fL����Nw5.g�=�����Av]��^�ǻk;�]޷�_��n^Znp��!��d~ߣ�iU�4��&�`����'<%���������Jv!�.+#�� U!�n�G  Ѕk�u�T��>ߐ�F�&��N4܇����T��ԫ�A��CeѰ�|T;o"��RF�p'�'�ߑ����e�'�_$I��$lb�-Ǹ����O����ėT����v�A>3�A�x��Ή�uDY֑Z#��� �ந)��G;�����>�xj}�0�NXfVSVP+#>��2�Ά�:�J��=z�+��aZ�H.��1@p$SKln�q�5��(p��(�ppEF~��7@`B]4֢�;ʎM��e6j�8�.)����ap��^!��P1I�K��b�(������?ps���x����
YU��Yu�`#n���H�<���E&��:+-H����L>P�(��9��0����gi�;f�(�A%�b��w
zq��_g�ɧ�: b�=���4{��[��讬���<F�h;��f��S/{��!�z,��b	=Ovg^���0d	E�bVE�2�I���Ap���ON뎴��p���$�<76��%1��`eyg-�d��B��:ź!/�&<^˳Gih+zw��Q~���.�-'���J��YP�}�Υ~�yl;��oz0ӻ���4x¡;�u��o|��5�4����\͎�0�T��Q��̏����E.%(�q��-0|�cR<��b�����NʸM�R�2z�<~���r�GK�)hl�+�@[t���=����Ƈ���uG�I������i�t���������b���7�+7��ʤͨ�3C�l�@�^Ԯ��u���� ��B�!?/�29�@VKX�3��G�ȡЮ��O��]��Ou4��D��6U��Ir�ņ�$(N\x8�zg��9[�@ݟ[�l�~�"I����t(���e|�-���I3(l������`|� �;�>�N{ȱ�D�(sq�<�� 5�5���'!�cV� X�����8���zL�L`��2!���Itk3��s�CFz�d���0��j
��Ž��"*{����)�%�q)~�ƀO��g��o��#�UT�yHA�B$�e��{v�A�P	�}y��n��a�$�h>���6��aIK�Pc?�Pr��ǘ~!�0���/��f��
�+
�ڽ
��֚��l�-^G0� �|+����X`�q͵j ����d��	��Bĕ�8{P������n7g�&�t�^�_�T��a)t�0b��]�N��q��kς���^�%��x0������s��6��ّ�XS���X��&��x�v��3��ŀyӕ��%�L�M�#O��
R��w�G��@�<Z�҄�u��w������N��T�5�e������0��5e'%��)���F��Ux
M�R� ���_ _�U�E��!���s�sX9�����;�p�^n�/��&�mf�T8'���
�/�p\y��%9-M>Fǹ����o��vLh�"0��������@�|���WC���{�:;��+�kbu<K���Oi18W�F@�o)��i��^ '�*�m��p �8w���Yă=V~��Gt�*a��EJSJ��s���2�
n�p�4�I!AV D=O�H��� �+����A�[� �T����`�Sh:12rc�	߹��	hQ�����,�=H =�'��q�Ռ�tȤ9���5~�!�>c�����EO�m�gv�zb?���q-���)�Q��FT�w84WQZ�\�{�:��zr�x�yP�b��|���sٴd�� ��Id�T1�Eq����u�Y��P� �:�2/$��)����s�׬t(�T��G�y�t�s;��4�OF�zl�.���!*{�l�r�v�c���y 7�w�u��� �4
ۅ̀�ƨ2��
���$�Y���>ϣ}�~+�@���*��$����\�oUR�̔(��W���e��^w��^O$�YgVU<�=�G��s��'?�}n��WXag�����w�P�'w��䥢��k�e�t��b"���`�f䣎�Z�{M,��D��Q��ǵ�cX@��ˮO�������7�������S���׈��N^f	�#<��uB�e��Jq��QʃJ?����~OmE��a�I:�$`�������b��<���F�?sR~�s���]��3m}�=*��D�U���v�d@h#nHpx7F��8��T}M�Uµ(�FGhJ2�L��s�����5�)���-ʊV?u�D�K������=]�Qe3��%����]Xv�fn��������I�U8�4aV͚E^ÃS�,�ء�ftX'--�h���9Dc�(����[2�tvoAN,�?Ni/	>��j6�Ն�y��'������l��8��Y��k3O������w+�h�*��wt �0��LKK�]�,,<�ʅ�������8[�����BIVc
����b��x,/��'LF��#��Ő� �����>~���=���o䄝��gW�UW.��(�UQٝ��>�s��l����C���54�����<�W}��\�`T�'�m�4���=|#Z��&�f'�]Ƈ�aq'..r}���*�	;���·z��E�09��ˡ�FUn�<@��e�c���LWߜ��45d���w��ހ�"��I�n��;�c���p�8�0�xO�L�5fLhqq����9��i�h�i0��3�ׁa�`��҄�ϋq��|�J�Wg�]%`���+��0����Yۖ���:ȇ��;��	#�S�z�n��Ϩ���->J�x�8�����<i��o4��/�u߷*�7�eLu\�~�?���ݶ��(���>���M��(Ð�3)z���5A"�g)��}Fԕ��qb`|P���v?h�;�Ӆ���j���?Z�9�5�~0��9�'�p��q�YC��:7M��:�ڭ]S)����o���P9tE?��ۺcpO��0�)	��7���n��.b˨�B����g�{���~��o�wP�`�3w�6wa�<�-V@���j6VȂ�ˉ�{�`0T�Ï�ra�|�#������3%%��Əy�ys$�Y��)��;��ůu���r	Ѓ}}Us+�cԄɓά��#\��5:跈~JL��c=�QT�<����*]���*$m% 0�?�D��9���Jd}�¯�d�n��8</+��gެKS�5�g����{�tm �po/�*;Y��O��ڶς��X�~��2s�b��J�ɪQ�8���0�GcM�.�{�z;\3VQ���l�I���0}ڷ��f&�z��6W��C��c�ۅ���3��qsؘ��X�Ю�RHZIu_T�1��zd2g�%C\��.�󭨭�5�����E\��>}�W�����A��J{4 �5z]�Y����:��� 7.G��@����u^��ZZW/�1qIF$��e�&�TM9	¢K��0� ���8�����:�	��;�o�O��`>��m�#cVm �\|2�;n�*.�{{GIP��Qd�kK�H��q�9lYG�>�X��X&#o�����M^)�E���?
KA�3���>��fѓ��{u���5W5��TK�G�s��TuLmc>aT�{*uLz$�r��Qv
�˂��8��I1��u�D���V�i�0rR:��/��z���(��p� I�49��8V8V/7GTn <���z�i�N=f��7����R{�\�e �#a����膯U�j>���G���(�0���l�3^����`c��}��된^�qd�&�9�F���h>q΂��q�9���JK���t"T�Mұ�g���c�b>YÙI���h���HY�WQv-��E�־�&.Oy�lܦC ��V���Ϗy��C��7���:����[w�g�� ,�'�����T�,�!J�ց�K���^v�b�|�<����� >сt���Z6��M^�;�H�����wB\x�����?���&[��Go�+����熜�8�G<S,�����j����
7��ʊN�����AQNK<]����糸낑8ъH��p���I�9��~��M�셵ൃ9\՝:*6v�k�������]���v�I�c���V̒鉩#d�ćo����?x�;�����h}���$�7�a)}J��\�����Φ�=�Yʼ������_>1�憝��� {$&t~��K��`��B�Ŕ/�1�Y���O�Q��svq�1���A��ӻMo�vcw�ިv�=
��Q�� ��Oɯ�bm���-][0�(1��`v�����} �$�e\�yZ��v@���o��A� ��+p�IL������f�����6�uh��p�/�[\]��f���!�7��;G(߽^�f�z�Pߡ�fB�,�����1?�W��s�_b$��o�5�&O×��ٞy�B!zu���gp?l���՗�E�4i�6�ې��ߘ�t]nY�b��k�Am� R�`$�B���>e."���� eA86D|75h�)s[�[`�e�����lG�x)">��� ���i�� [��A?(L��pZu*0���pr/'v��������>K�J��ve�bn|2�9�ɍ�V
���IY�8�����ʐ�ۼgP�
�=w�^y��>e�9.L��|�^dcw��{_K����=����_�G�E��#ޡw}���}��e��������L̾�f��3B�+h���A����ٿ����Zo��B:����W��x!�&}4���R�-����Z�9+�����n�n��8ȁ�Q]Q�'��@�x��H?{?�~�������L�C"}h���7F�OS�h\I��85��A�zġ?F�AW�B+��B��1~W���������}�Qo�D�E6���xG�뙛ǩV�����ddn`!�p8�E~V��!�b��0��/.��QY}�q�����,/�f����Y#5�q)PF9�v�+��{dk#ì�$��$ߍU{�)I��ь��4٥o�O�+A�"����4���V�Yip}�R��q�`Q�1���!�וR��$��8rFW�b'xui�/���r���4�쬀{)�IR5����
?��.��j�Yi8y�a^���:!�Q���H��E��⠾��5������)��r/��oL�H�g�%�	����x3|�)q���@�(��h�O�_�nc���+��l�m�U��fa�2m8M�,}0l`�P��X�r�)@ĸ��6���炤��Ub�W����"`6���U��� �/o#U�\u0�_��tg2z/���*�b�;�����Ĺ�D���m��G�.���I�s�f�	�؎d:"BkFS���ag�UVd0G{d�YO�$d��vӆM.��L�G�J��<�RJ$is4f|����ː��{��d���E�Ö�"����<ja�|7����P�O���~�{벬zz��e��������
%���T�@��̔$�Әpc{g�4Y>�!ibw�g�
7�h2�%�"ڀ�?�lnҋ~����br����DW�Ӥ���}r�={�
 �Y��j��M"�� �x&���y]`�� P��[̷��z��':LO� ��{g�����$kڢ�Ig�l������ƣ�M'���h;h��B�ykg�r���7i��Q#��w0A�'�����t�p*{��6Z5t�拤�.@�J�Q�Cխ%Ử���ªO�{'+�(��R5���_�o[	��8��69�E�m���R<zժ�@��s���K&O�C��11�����bt�fEh���]�,]�%�p�	�j�_��ݞ/`�*SO���#�(W�,���30�dݵ ���	|KF} L�?4�9"Tt~?���qG}��ج���p��d��0��r����^>�"����?7�vOʗ�1�Fw��j��F�L)�"{��ҍ��O��3��kQ7�w� �.;Ő�C	�Pj^5�M�x���W������MCm����%a_�[��F)�g�o��J(�8�,m�7���@�V{(�qPh�.v�l��r�C}5Pq!|��`��n]����l�1�p��8���y�-2�J��hՅ	�&�z%hH:Ĝ���=ސ�@i��M���ɡex�ȱ�|����计\�>I���@��6'6�'b�/Z�ℐs�e�e*���&�#f`l��U��D`��hL��3<֏��w�_�D���/�A�f2�RL�nݡr�cj�m���Ғ���C��ʎl��b�Kc0>e"�hzf`�2{Q�������ބs��D���P��+R��b���,�E�;uXT����,k���+�h|��,m)�%)����%=-�HҢ��z�sFDKh�X:�u�9O�o=�i��K��BX�bs�;�e� ��*�)�ܨj��B������L֓e�,�]�a�Xz`��w�8~��sW/y�Q�)���M�r�`lh%>�
`Sm�:RU�k�}p����	�6Ɔ*��o�s2����}�"q�vr,Q��9��q�E��/=��\���_�@���=wRJ�q��bl����	NP@#��OT�w�E�YԸ���A��f'�+~�B��!<����-ѫf_�N�`�I$��(�i�n%n헉;U�/�߾�y�e!�4{3Y��;��߰S�g[/�3�S�'��kl�FO��{|��
�e��PΕs�Ԧ�Q_}%�m;�E�N�?�f��_D���/�����mt�I�MV��[>��Ƴ�>"*�"0�sF@cF���{m��w�(Z�X�n��IJ_bL��g]���֨��NM=h`�� ��l�s�����9]�=�gE
�ʡZ
���Jm�p�ߣn��a��5�q��%?�%���d��VGFT���g��ZUx9����Zc��f�{Х���9q�7���;�m���i"=ͨ(��f�S��@�$��*���t�'������L���d�6Z�o���&�U�F(+�Q-b`��m<p�����ӢG��}h��w��h%�f'�ȑ�΢Z4P��DT}�ٳd�6�
kЈ��A���1\~7F�>����NwrU#��Ƙ_m�p�Bm���_�LT���ϛ�8gů�`H�q7Ӈ���0�Vngߍ����֗����_�ҟR��q�s��d0ж]�o��j [@��I?H`�vCnV�|bt�a,!dp]AJ��o�Np���r��,Sq�b�e.��0�.X��;��d-��|��7�t���-��xt�5��Id�yp�u�X���/qe�&�k��sHx�t՗T�&��N>i�kX)�(`�cb�0�y+�:��s�V�N�S���?��9����+m�u����سo�5��Q!�i�ZM9^&��&;럵���c�m��Qa��]��Mt�2���U�L�aN�(7�A6	�>L
$m�ſ+����H����0]ڷ�ֵ7�B��:d�4WV
�S6�u�o�� Y�h5��X�	m�M�V��ב���,���*
2H��Y��2��_B2tDe�QN��H�5�b!gMQ������]��x�M��fj�W?	%����XLw��g�q��>��N'� {�rժw��ꌉ��_6��7	�����tDȯ¢��d��!)@[?���|Z��.�H��%h�4�<zt�ʕ������GmJ�T�� �>�B��Kw�������!Xm���0r���;ϥ���=PR�8�,U��j�.`�CgN�)�j0�z��]����E����&�ٸ&�7#���ƽ]�LO�P��G8O
��xw��*�Ze�G����z�<�
X��j��Y"�]!���ؙ���ο����*;��(�cm��P9O��"^��·�L!���兽�t�7E	��N��I���Jp��zh�LIt<Deԅ�Y"Z�v�F�{uX�R����u5�5�8��`a�9��뾎���}��3��+���� ��F����?��4\�����;6C̐��L���󊰏Զ$���:ok�8���!�!�<��j� �,�����G�\�����e���<�@	�s��B?p3.��r�2�P�I���y&<(0gR��#��W� ��6SQ6ˬU��5�Vf}��Y���7 ��$QR��V�ʀ4[�)�"�N��v����Rph2H���QI�ֳփ6�8P�dq����U,2�+�Ὅ_�gMCL��"Kj8�Lsrs�{�5+�o��U��=_@��$��
M�0�)A&R�.�h5�������X��F��G�s��ٰ䲪y׬,�� �������w!�BHΈSႍ%���� �WN�P�466��G�Br�M�7g�X�������D>?�y�������Z*^�;�r�׮�Ф�9�V������a�ѵu����J+����22��~X����3f��~���c|�s/zH��;O���&΅ʆ!�q��+�k���X�{En�ON08-g���Nw���Y)Tk_W� �ʁ��T��Rl��̟�,�O�쬶�@�ΕƖzi�İР���P�>.�C�ch�ڽI�"
p�d��Fϋ�όj�T]��2
��W�J6��b�y����~<Ok���_�(�=ϓ�_GTM��T�O��-�o{��7 �w���I����k�����o�.��8*SΩl�L10��۶�d�<����yZs��gEX��p�qn���j�[�b��\�׋��,���ؿ�'/6d�|q�Q�[�n�d�\G�[�}���h����4 ��L��{�X�x5�Hi�}(��Y���������3�f�~�(�@��\���z@E�Ն���lъ�]�zia''���#�`���LM[���bA�zˉ��{K�@{��5��o�4�1�H�%���(��d7u�.�I�m���J!���_R9��G+��`����� ^CWXX���+�A_�!G�|;�c|-n[��\�˫� \|E^�����]�� ��OST�e�vka�x���Q�g�9Z�-α���7"�*��r�b=Q�b܄i�h�{�Ǥ���|�Rݗ�t�z��B�ؚ1N�'�*�:���&�xl#J�@�.#M��+��`Ğ:7;�+���9+dS\Rja<������v��ne��}ZJ�u/�a�~��%�����-.$/F�!P4��;�T����mJD����q����~�~MP�X�a����H�U��:�j�G��`G�R�Ö�bK^oj:	6{����v@p����c�ykIjϝ!h6k����3[뼸U����!G�/:?>�YR��;�lr�imn�h9�m(�/?���-���8Š�ͥ�w.������7�x��T��|[�+���=���vYm+n�Ji_P�ZbTf�R����QH?�͢4.�ؽ��8�#�W!g'/cc��k�oq#�E�q$J/Ӕ�0~�[�FHB�.���%:Ζ٩K�:m�Qg����~�l2��])�a��s�> )aD����[_�15d��ze��u=���V��rSf��m��;:yȇPJ��#�P���8�:8$��!}�D��S��',����XPغ����Q��������ض9�KX(b_`A�j��I(mAwL7����/�$������+H�yzt�0͵IҦ>ؓ�ҋ���@҇�uh�4�t*��Nn�d"&\����O��N	w{����Ld�Y⡒�Q���H�{�5�B������nG��R?$u,�l7��$�;�0E��g���U)��6��L�Ý��?���J�ŀ�lŃ0���:V�-�~�d���P�<��^���r���S�����K�9���bh��Ai3NC=l�!�UD�6���ff�����?�c������'X����hfc���.�o��;M�3�v�:W���؀0�v�n�itS X;�	���	�<��L	�  
�N��YJ.S"���#mj�nKIݣ;X/V�})�׷��	�i��SEm�Ҿ��Y�JΙ�L�!}x����o�S��G�9P�ʒ�a��B>I�(�W�g>/*H�X�g�}v�d��g�QDb�\��9]p�ڛ؛��FZ\f%�Ѧ5Jy0M�Lh���[��h�L��H@�e^Pƍ4E��|�ǫ\5��8�}˛4��at���0��I��������`ZѷG�9�x	�[��+j�\�%��e:G�-@4_�k%MBc��$�嘕�7�Q�w���
��A.�K[#��Po\M!ڧ�����ȳ����^ዠ�)�3+��y3��Cˀx}*4�6Po��^Bo�e �����m��!�i�ea�'�>���
)���S�M���wrϩ5�VG�TO^�̷�ĩ�g��Uv��"8��_���w=*�!2��^���gz��O�^�{�jn���9T�(�Y�"꽳�.�nY��h�\HL�ZcT�H-ٖfx�z�/9Kv[��G~:��zT���b{�`��!�x����@`L�p^瘊lYqs!w�d5�Z
� gz*SL�v?�f�-���S��wV��Y�@ �Sԋ��.Ri,%��҇��r��
��;���Zox40ԪO���,"�lR��U��n�[�A��*9m0�"`)YRm�h�Ч�1X�'(�)���8o�/�-�t��Oeކ������(^�f�V&P8&���k�/!�4�4�Z�z�I�e�}q����i'���#��VD#l��lI �cj�!��wvզ0{ǖ���{<swH�A\�q_�a�r�첍�����0��ՅW�W+�����B��WI�'J��[�Ϥ�:1�Φ��&��j>�v)�D�[6�P����H2,S׬$ж�`�F^�Z �4'���GB�_��Xӭ���qm>w�*r`!�͖*XG-qN��/5�Ϲ�>9i���u��D�9�$ՋM��VlwU�h �vWi��$�"�����4�"Xd&�&��6(A�V�)�[E#�����a�T=�D0���
�([䱏أ�En�����
ݴ앂l=k��4���lk���d��5�c��)���nr��d)�i�ɉ�yr�v9ɉ�Y�7�~�%�,�:q;,L(b_?e�kSHw���w�9/G����<�&ܠ�I�� 4e��34tB
Ggc�N�f=p�����[bO\�#�D���O�!ڢ�f�S�aȐ0-��K;��r6�|��]6S�MMX�|��]�>"�Q�
����j|���(��0�[,'���Fb]xu����\Mװy��Q���0�E�8�}���=�n���W'H��Tx�E9�D������aj]�
.[�2�\֮�[�����q���샖�pJ9q M*k�^����A�YBs�V��F��U�a&[u��?�a���"y���]�(WQ�<X���R�%M�>7rX���S��<�Þ�R���0>�Ϻ��(os1�[�2�H�˽B��<�=I3T+P�zщ�[�vI@�[A1#�t��TPKw-�Ѷӷ;��Dv�u;V�̊֘��iS���F.sx3I�d��s/H0�=�_aX�!��o����}�+Ax���v0�:� _$j�Մ�V����Ly��������C��d_�V��0;e3�s�f�X9TC�P҂Ve��R�������D@�f]�'�<���vG�a>�3�j��������P���0�^�!rڐ�f�(�N���^���s���q>XF��H�fZ(/�{�^�ƖD�1>�W�&T���FL� ���������E�-g�ȁ����B@Q��2_�Hdh}��gc�l�M�}���$��
��^�@p���Y��؏���s#s.鑥�$������>0C'��++�i�ߒIW.g.�\�'gM!��v]
�����]��,�;�^N-� �k��{RX�?\���l*X��ʰ"����h_��j�ئ�Kꃔ{A{��I�]`^�#`,H���/���������,�}A���
������@O��nF~��Ty��{e��i>I��}�'=���ʰ��EpJ�H#��Z
��P~>��Q�!IܫG��i�r�⅝�S���}5�hEqw2�d�p���NO{u\��K�o�5��P3�L'�8Gku[�$d��MN"y8]ge�va㫉2|i`LE�z�D�A<ґJD�ĸ<(B;����W �ك�0������ۢ)1p�Q��I`�:Z�v@�x(�+���?�K;��@�,��*C�r��{�NƘt?e��'�8J�#+�?� 	��J8���.s�&��hܕ�}N�|�b�,��P���	��W��Tw�`��S�{ㄹ�UO.��%�*x�rj���6�� ��^^�E��`UF�yrkjM�3Bŉ���v����:�M&���BH�SR�u�l�p��i��<�\�!=KT�(��6�c̖N�{�V��mSI��bXd��i��k��Q^����|?2)qq���eG�W����m(�����s7�"t�+){)8Ҋ]V��~�2n��'��*����aX�qnK��I`���ܙ߬��A�����"��T��?�|��:�.@U�|7Z.�/�'娍�[W]@8+��K�U�	���Pv3�)�h���z�*,�KU�;w�~���u�F+8Kg��� 9plbU�� o��i�ҝqnYeN/��GHX67��~>��SA/[*>��K��wz���g��J<�N���?w�KC�����M�R�"^Um��<T&�G�#�4/�������7/�9�d�G⾓#`V Bv��&�vi7����-N�ņ��pK�E@�3��b�܀��,bN���BfS��e�S[(:Op�ngֳYR������]�Xaʫ����WM�������[��/y�O������5����<]|�hi�U�s˾-���hxH>�3v��u^�߅���{���i�R��4Xke&5B��jV����-��;5�r�F<�6�r}��{� ����o����΋3���A��1���X�~���}abjå�h�	�f��
�����a�M�Gx���/ՍH�����
a�Eo�MA	nf���)J֭k�ʴ�]v�:�/�H�L�p�ȑ,�@�"0�C`.4�Q�䥱��Rv����56,)rg�{���q=r�;����p�-�-�J%��	�N^��&<'FP�c�����W�*,6���>�xB&^i,��Z��K�F�)�L�bU靨5S�Ϣf�;9f_�.�<��p�Ȣx�:���bމ:~#ADي���Z�,G��y�Hd:)j�2c�,[HÑ��b��ΎA�J�l A�{��"H�M�-�P+_n:�6���~�~�b��-��~���x�ї{�v������m��R._�ܷ0�6��بD&�Q)x�����%5Ur#��&;�4.'�ZU@����;�&,�,U��:[�t�8a����D�Ǩ� \�}��k.��e�둗3�4���>�	�s�FqB�&E�\�[�nŇ
��v�����kۺ�[��P����G� ��u�%q%)�T�}\'�!�ݶNN���F�F���0R�I�qƽ��x^Z]Y�v�ag�W�,�6���_����I?aY�\$�;>�grܯ1���c.5M��Z�Yqr��T6�H� 
ļGt���>��޷6��K����?�:�xrZ����k���#�% �Y���zsֻ�Z�&������Ѡ8i>)�L�`K���\�	��y ���' �͠9��u���ṳu��P��VrYS<��,�J��mŴK)G�6'QtΠ��s!� �WN��.��^Ԙ��I>	q�Vt���e�R���h/��dܪNO�#�S��g��N�&!�zׇ�a`0u��x���$_�Z�q�o$�Ыqt5��s���%�EU�����f������ '���V\S������M�1��	΀9k��q�#⁜���ʼ��lĤ}�R!y��|� �@� ƀ?��wu�v��X�e�7�çrK%��
>�V`~Gׂ�ĀH�74�6�ЈW����Gߨ�?C2�d1�4vX��3=އ��ɨ�R�����Dd���"5[�[�L*���t�xq���݂bC��B%m}�&8;-��o�b�n�<lӅG�,���Ss��'A��R��'�@�j�:i�y���xr�$ߜ�1D���x�d�m5+��4@)p.I�s[ݝ�]�	�Id@����'��np;�
IKn�#jѨ�#J�*�
��xG0ǯ�*h�����9����ƒ���>%�h�`���N#�p�j�l���^ɗ�[z��PQUD��r�fՓqHڈ{8m'�y5��A\7��J��v��ma�Fy�̈�����Ah���M`����#Ф�+�!�� =R^��
��ʜY/�|���d�<����Εىef�%�<J�ap��B��F5A\oh��.W]��� ��\�#�_c0�?CO��Z?}������F����X�D�����a'ۣ�U��o��%)�*���|���=��\�(2��I���-J1��;,gqPv�/��ObbMa9X�����@QD���,B��i̼ �O?T�68�(�FY��x�jӘ&��Kb=�k�uV��si��>��O&��q�<�2��~��T�`!�OfJ���%��+Dy��(��������b05TQt�D�O)NW��c_�e><T��\uvA�/t{Xz'��SI���I٤(��n>��l�+�]:�栁7��ރ�KuM�4�����ö��x5�r;C袠�����y�DL��h^N�|޽���T
 ��M[̄ɫl��$%��/OZ.���+��[�3��C	q�XW,\ɷ���)JT�̿��Wiw�j8��q���D���5��p����j�〰[ Q�Q��ʋb�T�Ax�H�i��]��=�G�1����=���`&�G{�!Zv�Jd��2ĺ)�`%�qő�U�p	��9�7y�(��T�2�FR]��#�y���}_����H� �|{��\�qe�~��J�z�S�ŷޘ�{ݎ��l`4#�wcs�B��Ce^�ϝ-,��Ҕ1g�3k�w��k;|�	��g�h2yR���4�i�ZHZA+�򊀷��^�^�!M��qh6����������<�C�(��b{K`4�{ ��+3�����e�#Un{��R4��V� �Q��Y��:�W��%@�g�x��Gؗ50N(��.���i8/���~A���r�o�}�=k��Y6´�Jd����s��n������2J��=��!��ba����WE�ÿ�e���MZN]��g_�ޯP��NӴ�����1.��ҭ��|�4���7_�Sز���&�5��ރ���	Zدr���æio�Ct����l�֙�F�� � �?���|�Z��0?f_aG��MPz�5c(<V�y_sI��DD_�+��~_�Up�&M��[��-�?�u+�N��/Dm�Gdkn���=Ǹ�������\/����W�fuE��9���<O�7�=���!Z9r�'��y��#���%OHM��V�1!_�P�w�Ϧ�t����tڸ	�n������.C��S\q\*���RWN�#������|Jy(<jV&�u����\d7�T!-}�P��s��j�4���H�;�'z��=��\�}9�t�[{5[�cU�`��A"73��D�͒s��E������Uiɢ�<?����n^��"N
yP�4���廪#�~a�]�w��S��7���+��ߦ��\+����ϡ�7���@�H'��Ou'L�F�M�/o��<E���t$H<��^�_��
�\lL�5��%"藸�\�	��h ���A�EY�qsv�>�_Kf�l��^�t��@�  V@��f'a"5�o��a^��v^��Ũ�j~�y=7��>��/�<_I��M�0��������5�����T)� =�,~ܫ2'��΃�O8�[������i��4)<�0����l�����Z��Ҝ���vI1�i�E+�_�2'���`����A�Vi};2қ	 No682�N�I��n����`��~�����jM�v���g�aŻ��7E(<�f�=櫑��<eVM�f���ԃϹ��z�����)�'�HLI���<���X�a '�y^ N�SG�6<��~�A����������%Ƙ �q@��G�r���v�!��9� /�S=��	F묖�zQ}F����(�Hpg�,���y}�/7<)�j	G�Q�?.;�:�nn�N>S
I��K�U#1�JTyo�-`Q��⾅�˯���[y�H��Ĉ^P�t?��e!�4��e���(g�V7sJ�hX�s6+Ă^{H��8��B�����oU�߬���fG��wZh�̜q��<>�V���g҆���\�l�n��>�:Y�cL$>џ��)������똉�x�ʩ�����Eτʈ:p�'�b��~��v1���M0$��MbD2��Ė���ܸ��:;+"�t�����;?�`~�b��Y-�š���� ���2�vl����k,&�wM�W:��j�'߲�f��{��2�d���z\��A�����B�Os�G�VG���o0{g!S�h��W�'ϩ��4(e'y�� "\�ƕ1�
l�������<*�K�)���5 k3���P��40���&�\�����$D�Q�֠� mW���?i�Sd���LO@� P�r�Ɣ�u'��5�W�7)Ш��D�(��X-,����#2�	��4�{�15&�'d����Pֿ�"�3�u���F��1�iQۿrtg}A�}��nO�3~����Ϡ����j	L
?��ы����Li��ң�^�m��S ��_�8���.�i�٬qq\��l��cm�^L!������P�了�H�ҥX��v�K�5!v���tG@7U:����h.7���LN=�25R��=l}��x����K�����w1VR�$!�cVYP��g��\i�6�t�<L��l48$'��]L���cO�]W�Ƿ������tA��Ys�`o��r�5�V��5I�rw7g��>,��կw�M���٤�9�i�?{��-������g�<��o�����fSo7�Ѕ�,�'�t
�è�]�{1�iѵwс<����|���Ml�^�}s6�r���*�Ӳ�z��?'�Ò��y�� �"Ԋ�+��R?RQS��8���:Ԥ�S�\�/����m�ӎN���t�Dla3��5Pw\Ԑ���(�Jf#��Hщᰠ�Hӄ�!�=�����>��_��]U�D� �$�c����ۨ�^k� Ǩ��"����lq?� yZ�y�i�G�y�����c��� �)�w��uܢo�}����;<E;qb��ϊI3k���/ta��c`�P�E�0Q5\4�����<i��\�=}3��D�t�U��-��Nq��F��5�~���8.�MNX�J��<945Ϲ��k���3/����
�dj�]�i�7�O޴���۽�Q�$�ms��ے�r�O�5��G��0�!f3��2F�x�I͵�~�r$3�C[6���^�a�Kn%���L�i\e��8Nt��U��%�$P@C#Ȱ�����ܽ�l��`8A3�S�I���"+c��rF��~ֵfQ�DU �D���e
�X"b?�SD���BE�w	Q�q�h�<�dq����H���'�������AsRBnK�GF�f�B�f������?9(W�]���z��ư�	��|ӹ*�X�x�+�L5�6Vk�('�eq�.(��b	�p�+>}�=$x /����^��#1>���/�B9�~h�y�\f	��U5�&ď(��@,?�]���ڼ��Dֻ+����t��^	2�3���rd�@T������K�f�_M*+_~�4e$q��˜q�]q��b��{LT�_�X�jP��4:�&�)cWQ��y~�ޫܨ��C���fO5M���f;2(��;�*�.�	I���o<f�ѿu����	�-ǖ�֯ĕ�؏�쿩�e.8�������d��Z�Z�Cs�\����駯�dT���@K Re��H��?�ȩ^'�|ܠ�c�XIu~��q#�(ݕ�	V���Dx��F����
���
��Lȓ���P=���׋sW�j�c���;��<�B���>�.���
� ?�U`�����Ӏ���M�JS5�g���f𗿍�0UK�Fr'�x���J�/֟Ğ�"p��A������������ �F#sTp���)���A˨�ygG�o�U�lz�WλlI�kN2j�R�&2�������V0!�,F+���DndG��k�.��+0՗$�2���"��B@(�/k^�`�9��,��:����l�eg���Gd���D��K�HA�Ҹ����Ǡ�-�lR�y�Jkʿ95�-h*��?	e����L9���	qښ�L���:ely"��dߠW#S��������2��>��^�Z.!l�"3m#]D�mo�"P�s�C�h*�s��jF�+.��#Ɖ���j���~�ă��Z>┟$ʎ�P;(������|_ā�͡P#~�O���h-����ʑ�nM�J��[@ҥ����eR�-�>b��R(�	R5��$6��p
~
�)�q)1�c<f���}�O�u���QnQYe�*c�c)J�
.������[���������ś��Gfk]�6��o�C���)���5�Y��f'u�u�g�vS�Q��"c��S�
K�p99ҳZ[��q=��S
�񹱔t��ca��5����n��='y@������U��|���7�)��W���\g��_����pb�L�f����!Q��RڭA%�䨱���}��'��m[2r-��$[�u?͌�z�����|�U�N����-2�v��H�CZ��I�����B�,x��_a��+�����W��0����W�9��6��b<��^@iJ���KWtǙ�)��G�~��j[�T_�n��oUz'S�<NCj䬢�k
CA�!��t��
|X��\���e#�&h�v�J�4|pL�
���	��Q�nd���q$u�p����4��30Zv�<
Վo��RS�Y�nQO�F6�B��s����/��_�;���r[H�1��P�3�aJky��ټ��& �+�J�|X��Y� ?� 	dXJ�0o�-㊂Ь�sb�FZ��h�~��]�b��N��/���_�Hܥ�xܱ�8���i�	yQ�����$��rU��.�`���s�2a><�k^���&������������9o��ҷ��e�<3s9!�C*�-�AQ/��֢z����r�d_jͅ��B�D�������瓁u��Z6o�-�z���~ 1]f:�=8"���G���'I��ȴ�kG��B�W.��a� <�0�ƻ<������b33��%"�y�]�1`�/W�m~1}8�HlƄ��ɼB�VtP�[�|3q���s��f#��x8��G,F��Gv�^����D��6Sm��slBҘs�FH��C�B�$�l_^��$	�s6lECL��l3�.�a+䐛�S)b�jK>�}]��H�����)I�z����P����Ӡ�������[�v�Z�}x�m����.EZO��H�#a �ƀ�?K����PD�z
Hz��5��R�����C�X������O�g%��wq�����(:$'C��:;��ff-�\_4�;w�#x�Ѽo�R�9���[�4 Ÿ#��^5�i�H�c\���j���X' �K��)X) _�)u�s��$�c1HC�g2ubY�P�Q۸��K�v��X&-Ma���qbR�Z�/�ʔR��NɰY�c蓧�i�lM�<�D��b��Pp��pWn���	��y>�����J����l�l����Dd������R6����>�~W�Ո�Y�t0$]��>�v���i���Y��JB��6�2�Q��6�*#�����U�I<�t�>��>c��d^iZN�\�j�����sѨ�X� �pg������eRĿ�׆��v�j���c$ea�ቕ��p4�Q'�v�������=D�%N�B����3����yVq����k(!����CQ*�Ʈ�����5cZ���3�U�`"�J\Ob�Ki�ɔS%1m�x���32��A�1�#�+8ز=#$�9wu!�F��@��1��$E\ii���,Qx9M8�~��!������o�J�O��}$��8Y�O[�(�A5�"�z���ab�v�&Y{��yH�H��������o�E=���0Q���ϔ��MY@M��d� �o��;e�@05�7*��h=Ă��N�����GY�7��5u�����SV���"��Q��d��6zsCE������EI�3[y��C�e�Y����u��X.���%0Ӛ#�)���o���2L���->wN�2�>tTD�8
�4o|��~������@\��o��(�i��"�"��#t�1�u)6��m�9�Z,ֆ)qȹ�; ��g9f��Q�HK�+��»�!Y�G�W�Ct��FW^�oAj��Stm$�ƽU]��^�O�@�~0�f��3W%���g�����r}��F��;�(!惥�j?���iO
мl/~���T�܅��<-����|)3�A�/oD�n��Z̿s�%6�aN�������(	VhkL)lyv��Fu*���
'�8U����q�B�Mj�ڰ?RQ����F�F�$�lf(Q��'	k�3%9��5W��/��3�M���К+Z.yZ��?xە�G�t�sձt1��/d��"A�C]E��;!����]3d��ցD�:��9��!��L��W���|Ȍ�����h�)+u�̽����~�媹�YK���[v��a�]�D���L#+���05D)��(hS�Kg�ꑮ: ��8�K*�MH�
|��7��@C��cY�	�{��Z�l�� ��#�H�Qp�sd?~V
��BƎ�,�����Y�	�`�N�*����8����&��0���s֢�)A,<�����m���[(#,�wB&�&qR(3�Ō#�%�K@���K���P��M�+V;�]�SY����[��������0���P�_��S�\Æ���uJ�.���V P�E�Y��oϗ�e��U�vJE���7�:R	�	�����A��úm���pxP{�@z'p�"��:�����֤�Ӳ�^����N����[�qF�r��OڣB�q�����n�٦z2!o/�Uf
�]�$���������4�P���x��i��>ݧ�o>��	�=�@6���Y_v��7|���O��@�{n�8__1do$\*����+�+��<5$��g\�\�Ge1���Lh�B]M��~���
g+>��<߲n��f��Y+�
4d+Bؚ�.J���������H�U&ԁ	�C�/���f��*gK�ԃ���YW���^��I
������-:F�3}B��k�u�v�T�#x�+�a3SG�؈���4��P_���=���uT�ۜ���h0\�\/Z~؆oyTRv3�c[~~4����7(��K������?�>������S��Ri=��P(��;�E�?��vj&N�a�Z�d�K��^N.�:M�nu>�$�|1��nAG��� Z� >���E�C�?fL$a9Q�_v,����L�5?m:��r���e���3R�ߚ�ZK�G�影�~o�S{E���%��Sp�����O�S�i�o��0_ϊ�tu�W�������@��������_�:&���.�$���
��A{�d��u����:V�, �I�r曚b0[�ۙ�	�l���
�K`t�Π�[��3a���`��r����C�����Qc�..k1���e�rU�� ϗO��=����S�0���ԳN�nOk%�N������d%�%G�+Z�R����i���h��6������dyi�=I�&k�lo&���"$��?}���Na��F\ڑU����4��۰�>�Ӟ��2�����2ݯ�#����/�6��~m�^tpDD�-A�a;��\K���Ƚ��6��'�iY�
����E ֘+��퐐���0�t��X{xY�}���qHL��i\�� ����f=��`�}᧝2�\t� 9Ue����X���֪��#[��Xo�wҍf\�%�0�v��� N�En D�.�v<$%0�����j�p�-����F����W�_�Qyen��F�[� &PuR�6t�����;kw���(����L�UQ/��9pU���\��b.p}�t�S�Jb[c#J�^��y��և��4~AD]��=(��k@7��o���������ٺ��ᨄ���%}���cuUQ�,��4���D��-�+�<b�R1��Bo��c�Z�ޙ�&����#K�����e��*�
��Ts{.��T;�����6b����{Hq�)�=Pl��dY�� �Ԩ�oM���������'}���-l�o�V"��*����v���<	p���շ��D�=�]�����P�;.;���,�O��'U��2��|��}7�s=�z��B�q�9{~�v�3#�$��m�30� �
h���/c���@{=8�{��4b�S�V�%��P=4.կ�mٕ!�����u�*�*�a���e�
n�^"�S\W=�ԥ����
Fat��=`&�갑z.�gG[�'^�i'�QsA} %���8���riF{��s#�+��"O�A]���n�;���S����Cˀyo�3��`w d�UF�j�_�'�̏}�,��_u!A�+��4g�j�哻��<:��n��]�@e0���z6JЇ[`��2��0��w��Ed� �f�s�N�1�]�S��͚M(%�sg�!�63�T�G��Dƣ�l��@�]��վyA<����e�
%�}��Ȑbԥ����m8�B"��={�;��cn��0�Y��Xw]����HzA���L���C�Vä��n�PDt�ˆ� �����3d%\�{;105�xF�zu~��𰇉7������>�ĖR���e��v'���V���d��l)?g��K���]�y��E�|��4�D`�l��]nf`�=fw0�p�y)a��j=>=$)��d͇$�o��`;�=3���๿4z��1泰ʋf�ڔ��Us�d�_��.�Yz�J�����5�_�����ر�~��5,���o\��{ѭN��0�����G5R}�����ʎ�`X�ɢ��8��Wt��Oq���\6~�J�O~@b�&���A2�kYDoa��?b�a۳��>4�ʯګ��j��Q����6�����gT�h�,68�*
�U�۶��	}�(h�~�+X���;�-�c��`�����O�Y|�8��!���m��P�(6��R�����)���0*;�M��QH����D�Kxh������$�|�D*8�AuQ��c�O��Re�x*�9��Ƣ�_����6���Ͷk�F8�c���@[���2�WEڹ'K@=qC�d�I��Me��=B�}q��*��v#��v���-�1R-{{�kS�k�"؉�6"����E����S~��SD�8LѺ����=#�h�i��|q�ѣx�;�瑾B�f�si�'��T:�)d��sB���&����z���1ȗ Ӯ��r��"g!�D�r��f�塼� _�jQ�L2š6�����Ŗc�K�'�hU�ɼH�M����Xk<�=�����!9���H�*9X�GG��V�߱~��e�@��c�����0�:���o�p�s���a_��UUZ�g�(
X�ي�y
,J���bo��GP6et��۱�QN��sN���J�CM��(y;�o4�T�dWZ�ǘ���x��#��<�m���ۓ�m���`Ӱ���䉛Tu������t����|�,O�0��t������ R��AB��Lm��~�o��R��1c�Q<�>���T�����C����{��o���͎�m�e�v���ԫ��E�w��B_V����	�V�h��jTR���\���+HY)旞���1�(���3,x�D$�i�������R�$h�IZ�^�s5�� �Un�H�;��CI�sꫢ)o��0�����:.r&/5����rT�.�Ŧ�t���J�)���	�x~�C�1��s"Ag���p�j�0k�;�="$k��_��,*��wb��h�u��^��2ED�9���o�*��W;��f�����±��Z�{"���VM�|��>�����Q�Is1���W�mϸ��"�$��D3(�U�@�2��?���*㪥�j`��~Q��Lq)I�E< �$K49��b�t�+�&�`Ѻ��>���9���Z~n��a���Ȯ6}��0O�#^?$B��͌��('q F�~of�v�Bdzu���&�����N�㮓9�mP��ȩ
&� K����w	IA���=t��b�A�ub	����o\��@���7�i�Y���{��R��oX��q0�b'Yw���hO����2��Z�NSA���[Ը^ K�*5)�~%%s��ʗC��d�q��c�"۝L���;�2���7K�3"7Q/A�V�'UJ�w�L���v鼱��/��5Q�(�d��sAQjf�ڞh7��S5!�au&��6�FH��f�t���O�ў|M�۝C�K?��`�n�,�O*j�'_pa����P���N�k�P���9���p<Nwn{N�K��|n�9m�x�
�9l-�0�eM�*����]���}�wA65�kWOE}���� ��we-�]�h��q�������VN|���a	����%*��S�Z���--ҋGMg� ��ܡ���v�t/>���؇O�)1��M즯�����w�@z���'����4]���`��x:E}E��-~�Nx�؝Wv.�V�<�r擋��,���k��Omg��d%\�d-����6!7�tO���X��
�|�Su��P	GOJξT�Ƕ�^�OO$.�qd��-V�Q�+{��⾇��羉�,�
SFf��8H-����"_�xА�"�`�5��<��*���6Z�ň����n^6�}��*��zƕ�;_³����'�Y^\h���6�K�	��`��5�����WG��S4T	
�����(Пn�4l���UXǌ �����3h��PY���Ѫf����Y���.Z H��A�g�8��?�����o	�`��S�fvU�4UY%W*\ƨ��������A����A��4HQh�м�[��Y9ͷ��3{[�9��]�{�A��%�2��M���Tp[���_f���c�q�}Ĕ-K,[C��R��<�(�j��n�M�w�r��Kw��̉��3:��3x#y�0�����1]�e�YT�K��)8�r�X8���ӔP���1��0����v׻��:�%'�c����M�*C�	j����{�W�%� 6�k��5����T��EQ�BI����s�Q��4R���v�F�uF�b��]��Ff�h�@�AӉI�zfE<&����5*��L��"�.;^��~P���y`q��]+�=:K'��t�Z
��-��P�k���զi{�bX"����}���*�P+Q'�Biálp�F�7�<`�]�e�Mj�/~$�+��4Q����+�R<:��>\Li�&�Ã)�����oѤa��y5qv)o\llA�i��� 
�7��?��%�7�<S�/w�F*d%����/�ߖ�����Q�9�z�$`$���y�[Eܶ�8]�5��#5�߳��Z�7��R�E�.ԇ14�7AO7�:�#7\�t�F/�nM�J��'M��k%� l!�F���f���A-�w��%ܡ�h������I�h�-k'*��u�0x-0)���$� g��C�M�Z��]���y_V]g&S��&���N��lg0�AV"G�Ȋ�/u~�?��`�aEpcG�=A�}a�C��^�� }Έ�#������=ǔ�7�3ܛs��J���y��Dk�s������O��ɡ
��l�><ƫ7��iw��j??��Х���\�3�($f�D �I���YHi���0�s�����p�g`S������� �a�9R ��A�q��5�X@��H�+���[7��7Z��^>��̛D�%1YR'�L�K�Fd�����ۗ-�����v>l[YZ�5*O�baehV��T`JW������,͘��4�26�H#�6<_����=����~�P�o<�\���l�C)���6�#�i�� �dI���Ađ��8�����P5��=˕��,�Ӥ��=U��5$�E�����ܸ#����?�ʦ��#�[`�J��W�K��� T�,m�Jh|R���D2z��� ��ʥ�]�u��&�\L������}�1�9,߮��C�Ed5$p�����.��'<��V�+G�l�1� l�ާB�9��{r����A�����i/���+ �[��A\�F�>��gŞ�5ݘ�����+T� :!tN����/l;�8�q�3�Y�
xQ_�:C�)�LL��Ok!�v�h;��w��}��H��B�!	'A@������a꾜�1�*#`ǹR�9�ײ�ss�lX�={���
TR�/�c���1Yz)������H˕K�E.!P�r3�7�ڋ�F�St �=G���Z�"���H�Z�h�!=�sds�qj��P�b5(ꦒ�K뒁o�W3dbB2} ���ͷ(,]+���W��I�	�]�J��ŮwM%")%M��R��Ux7�я��^?b~�3�>��FU_�^",X�D���*�1��9�G�i��z ��V�Q7�E�C(�p���Ku+5�6C��Y�5�E�AB����1-�K~�哏&�fv�	4�%��Ѳˍ���jE&F�ݐ�[e��S�x�&��~��]'��p�`�3o��"�Mw�&"�y�����G�y�O�l�F����^��B0�:�^����F�M��$Y�B�`p����ӯ~��6���o`zU�4�l������:F�7V��h#K��5>������f7�j�u���/#+��Fƴ=4����N��r��Q�CZ�f�&����zɥ���8i�U���])�;�C"��Wo憠!F�p�`7�^٨�SH��~��oW��B��_��� �1���S��j�{���*��.���;f���x]G���v�� ~?g陆ؠU��RW��^U�;�q��$�QM1C1� Uğ�Ns�iz������t�-����6b+*�M�6��'\Y����� �'�j�H���	���!zg�_���O�:R/�
<��k�����Ϩ^�����T��7Wu@=�Y��RH���(0#x�":��,�K�?�G����>��U};?�W���|Uy�y �d��lp<�H�!�qp'���%|���� ���'9�o<ep%F�@��|����~�FN��XQ/�j$~��G峊�{l�jlh�R/T�1n�^O���p�'�ci;ޕ=$��i83�0>͉���'�@��L�*s���@r;�)9�J�1�~��و�W�Rᓦ��)\/<�9�=d,�v"�- n%�~J�"�w��&N�H������7%�]���[�ny�R$(�}k�xh����hJ6s� ?��4�9�7X�����wF����E�>H�}������g�d�j-~7���5k�k����6��W��.�4���n9��~|Y�̝X8i�$��U�W�-���֫�����QK]�H>*@�0O�e�A���6��aPږ�67��Z����?"E�&W���s�`��S����>vs��?�UA�
�X��Ҽ�4�����.�Pl>?�� Z��>�E &R��߹0>A>ϭv�,d�4�Cyp�M��a�=1�F���7E�%7mǸ��I��2�T��0��N}��A�\}��-ZFlW�?a�h�}�b�֞�א{��3��J���,p`�'w4�d�����	�� �SꈲL�BJO��*m���htK���	Q~��Q��l2�+����.g^>+*�TL���ޖE�ǐ�9y|S7Q�F��IH|�~�i
{%cN�� ;����f�KD�6�v�J6�����Cv�(�
�F�^����T��OQ�1��}�\���N�z�ǃ3��98�v���?�[��Y1}�WUi��;@��p���~��z�����H�Y��E��s�g��=��n���@��;��<�b7m�ر�RI4 V�	�f[�،�ݼ:
�^��$���	�
xiN�p��|e/�ho��,WJ�~����Ȣ��w���CY2]^m+�:�L
��9L�&�.��I��'ۓ�����kN|��5��K7UA�ԩ�ϑ��DnY�����ˮD��>N�@Ca�w4����,�wrV_�`�5��;���i�����O�8f����m���e6���~���燣&�y��CBŵ{�+��U���ьQQt��]�#�o��1�u�G��#����K�	�̔�u�czS%�ޛ���y�Y9�?�Lwi�)@�.�W������+���������u������B��S?�w�P���s���k����;6�i�ƭ4�����=@p��+R7�vø]���Ýf�΅��+�8럁�\�h߹��:*=t�
�qC�aH��?���@�p���ݚ:���Ia?b�{��f
����+�Q��8�&�u�GH���t�������fA���!�X�rgw�q2 ��E?��4�+��fa�� �òR�h�<q�[�0��ɰ�i�M� �Jy�\B?��ɩe��IZ�"L��B�F��-5ċ�#WAk�ta%N]�^�L�����BH��C��<�����=*x�Ý���C@�� ���(��[*�s>��g��a}^�%~L�6J�z�f5�tS����a�1��AH���'o����<�6���SP0�ǲ��ՈI;'y ��B��j�e�^wwj�C/
�N��Sr<�v���z�:��a��_�<��ُ���4�0z�	2]p�	�t�2�_�N�>;9$lm]˳�h���/�o���x�R�%8eS�$W{{�a���Qg�$��]�j��1�q4s��uN�E�rD���/yZ��H�A2��a���Y�z������ *��q���­��&��f��1�|��"=8��ί'w1/|�u�<�y�S`��P���'Ԇ1U���]����X����Ǯ9j���&��2Z�bj�s��ߓ1ylE���
|Jϯ&�>��Q8ĘoƝ����_�c���+�8Iݖk�WS�3���$b#��3v�92`<f?J.Cd�i���f���kp8ꃫ�9��HiQ�Bmu�#�*@%��j[�d�*f�~Um�\������$v�`���jo���� @�l�Ԛ�9�[�D�߸UP[�}'Aؚ#�Գ����U �\
^Ӻ&*1�!�E'��J�p�"���h�񳮔����0e󩵭b�t��^f-���y/aU�C��Ep�S_�|`�+u?�XD�@���J.m��F����~� 5��N�����f�e�Z��Kfi�-I(b�@~4�Z�/|��Y�j5���E��$t����_��X/�*��[S�w���j�>,϶p���R�������f	z�������ڌ���	�|�Ҝ����0јy*+�l"�D�;En�nN�4��{GD�
O0����	i�F�Gh-��W7HI,Ԣ�gX �C���-|3G'�*Z�����|]�̥�h�����wiJ;�tB`ʤ*�F���f�_Q��-3W�_:8�	�U�M�� ��g���R"q�I�xۓ܅(�/�Q�t^4��x6��%x"M��[ ;�z�ap�RB�t0�����S5L�`���7�j�T�}��������uI�I�1]�-[�g\ �`Ď��t��hom݇s尸ؙ���6��nU�{���rr�=�����fܦ���V?�H������3�p�k�Dl#�њ�k�Tl�o��q��Ϋ�Ff|���."U�N�ݡ��l� KL�D�.⺗��ڒ��|���__[����x��~僯�Wi�d�7R��I��Lѵ�J�C����+ ՗r;~�BJ't栙Gu5[�:�Mk��!�r>�/������?�`LX�'pڂ$�#(oS���d@%7��x�oe���i8>�� �y[le:Ğw!�ܙ^e\�8���`�9�8>����h��&GD��i�"�r*���9$N^�o�\f��>H9��U�_RGz���z'l}���f>�_��A��R��ѷggƢ\-k�����DT������G4�GƗ��=�F#�J ;9s�քo#�W�xs�O�N��<��噌�1Cc2���ʚbԵ+��`sI���CH/�-a�>��������pM�t�U��0sFƘzM�kZ���m|n�='�^!~�ae�����Fo��U"���E+���[��R1���U�Y���%�E�k�i���+�q��1����.p���_�P=c�(�1��1���Y�N΍UQ�;�$���4o�7���T��~'�g��=�_��
+�t��"�ܠ	�@��l<�;�2&ŕ��߲A)�C��udI���ѤA>�e�(�-pBO"0���Zd�[/x��*�Q��A��>&����������ߵ�������D�h��8�VE�w������uM2�w��va��y�M�v���l���_�KL�yY�Ed�8TvO5Za�|�e�R�9�NXk� ��:��n÷��9���I�ZNO�њ��
u��M�f�	{�g�G�Òk���j:�c����T�u�i9B\�o��k/kp�c	n�ۓ�Wg���4vO�vO`����.��.M�3t�BD����,_3�^�lU�s�(Do�P$![�|��e��AҲə6!�WOe��� tN~�������'8p���ɲp�����������g�����?Vn1�(b����SlMþ���*d|�3;��RFF���&�w=o�W-��e_�h
.%H�x�� u��=������P1@2(�O�m���K��²Χ�'�7���h��\��RA�RFv����"4�#�V\��X�b.
�~��B�mtjQ�6&�$}}H�0��(Kpʒ�/��v�ǲ����W�X��ch����g~Ȯ{p�#;�T�TϟΛ�B�d8���笚.�P �ݿ�-�<�'~��/6��c��-�֍�l��ؚJ�/k8�_N1?��jP���ю�`V
�;R���`��
,��1�i	�+�w�M����{<���") 0�Ԩ���Wa���ɨ�iP�#n�����O�t`$�T�['us1,C��O�#�����ᇳѢ<g�כ��i��x�$X#|�,Q�%�w�N�\�=[딎ttO�!�ʝ��`���h�|Z��×��<؇#�w�C�͉ ���Ӊ�k�XJ`%�1Ah�Du�
B�������8���J�/{�>a�] ��'1��Vף��V�.�M��*%��1���e�$��E��cO)/"���QS�2�W%�-�&��!���1z�]X����vG��{�m̜�� �c+��w9�?��:
�)-�&!�7�J�� *���#��!�-7$�DOI�V@�Z y�X�_^�0�|�[����޺۩��3��w�������#@/����M�[�v��]�~���&(P�O�@�>8�j)�GW���ɪ��d��N1J1�y�]w=W��=V��q�`A¢��z�p����,,iLU�ӋѺ�T�]s�K�N��Gܯ�sO��3p$���kG�����Xő~�[N*)3?N���5D4^O�k��r����	:���5X���{2�0��;���#�,еA��P�����S;DLQ�����JY�G%�#��έ�p���p/6ۨ� 懿j����.WS�ϑ��o�M��ı���N��Zv�ZBux�W�B���Wn���MK�ݔ���	����Rk�a�x8,K��PΥZ���Hi�ZfM%M�T�+�o�rw��,�T�U� �����d��ȗa���2�*�9fH@Mg���0M�<��d� �����"��߼�F�|�O2�c�ԯ�U\�{��i�X�~9k��D��k���Bp��G��)�K����7�W=a=�D�?ԗ�^��k��8�A�F�s�&)��
b ��N�vǜ�T�%1U�.� �a�Ze!o�S���}
=x�A�6nED��V��h]h��YO��-#�뻴\���2���d��S\+�o�B�5a9F��]��^�zV��
�r�W�}����}��-��k�hq��>\�|��܍�M�I$�,��^Fxt����6o�hl�qb��jבB��f_6vփյCxڽ'$����Ϟմ�e�杲6?����v���[Q�^�Yz:��UGo�wפ�o�>�����z�h�+�?����8�!W�ʠwo,%î{�fwğWP���7ahH�63�����_�)��yVaO���s/Q��1��Kҗ�z�ݹfY�#+b��/J�B���iXkbv2+�d��/��?.%A�I=��	(���m�&Mg����r���⮃XåZ^eC}r��T���	���A�kU	��2Ԏ���r�~gY�q�+������V��
/�i{Jb[�3���6�8�y3=�̕e��+*��JYQ	�68�rxY�=Rt�'`�.�w���G��"8B�q��Z���+V�����`i�R�(D�$Z�9�{����-8��KQ��ݦV�Ew:'sJk���!!�:2 ���c��4���p�ka�iG,����OL��ȭI@9��ꁑXr��B5�c��t=G��`C�������MH�c!�{lw���nC)tƄ�`p>�1�8�z=��3W���H�t�$���ߡ��mi��1]]��F��2lu�]��(��/+.��[��}["^>�2���^>B����`���ʍ�o����@���聤�æe�gg�~�����C/�Υ��o{�Dyr���]��~6���~̟ak>�	2�� ����5a���x�_��W���o?��ƌ[��d�\L/�]U%�K'�|���s�OD�N�ٯ�����iCә��rV�@Y8"l�}Ը����I�7Ƞk�)�/uO���q����8�0�ȥ
|BBS��J|mߝ/,�=���΀1��yg�TkߣE����Z�#
~��z��q�Z-@�rj���i}�K偶�*�۠��ي͓9�Z׆*��Y�t����D�M�v^Z�'(�j�<T&y�H�!�l�M�4��c2!��t���{2a��^�=aV�!��E�H��B5,M�C���3:�*���LIQ�aO�J,����Lsh?"X]�x;;�pA�G'�5�.T1̺�wэ8�d�Z�ا��-�]��]���Ea�_UK4S�¯,�0�h�3%$r���M6�-Z��p|�����a?f�sU�����ѭ�M�Wzm�T��:e��B������*��M{&���${Ϟ�]1df�M�ыE���
S�P��4��,n��>;�T]Z�!XTk����
d +V����XN,���*�3y��G�t�m+��D��(�k�Uʔ�O�|�]g<��L5�H
D1�~�%�Q�d�זC�̭��ᒪ�鴶��P��֪)��X�/R�#یBj����;a�q�-�S�9S�0�Gssa�ƛY2�.�2!����\��*��vJ�ɯ��<<d�n�w:/d�S�3�H{m������A�䝿nF&�Խ����۞�0���y���������n�5a�#}��P���4��׮x<=�C�0G̦�n�N�8�
�k]�#{c^
B���9�ĺᒖj<K 
_�]�7u�"Fm�V�+��������&�7�RL � ҹ����a/��a	ɡ1�\w�_FJ"-�����n���%��G"�q�F�0�2�U�s*^�@��ڻ��Ԍ񔟍��~����'Ϊ�;�j �9�ϐ�y��%x�z$�dw_a�%Ԝ��Ъ��O�D�Zg8/�w��]�Z��-oR�IS+��D_�Zf��h�.R�������¨!�:�En��w�˱��ծ�t��OF@D~��� D�}Ԙw����u�2Q��Q�#��+L��gԶC��&������B�d~Js<��"g�S�w��)JA\L�P���`o���
��!��X��MYբ���8��H�4g�����ƞ���f?Q'�QI}%V�J��(�"L��Y�0 YQV�׉��	���#�5@�w���P��_'�l�hq���5\tA�z�#~�}M�z���˽�~/��ƸnL|	*���<2�9w=������N��]�öI=)pgѯ�S�>��!���\���5�Ct_V��/��ރ��>��f�b�C*�TZ-�}Z�ƮI���Z��C�ϢF�[�H�g�^Ȝ�3�E#_Cy㠡���3%QϨH˽����#��V�]�Z�fNid�!��*��pn),J�O�.�io�:��+�	M��N|3�;���(����pc����_h&h�K�÷0�h�W���=�z��=�#�_��y�]����"��<<:	����2��F&�4�C���mOA�~�/�)�
$�W���z-^�j1꼯uD�Ɠ�#}��ލ���al�8��}S7��t1� D=���2��%����Im,
2LzLn�?̘0p����I1U�:{8e�����>�w�?�n�p� ���t�Q>0���w��X��ULuD�>�tI3/�x��E*�Wէ��n�2����f��T)�#Ȃ:�x�,�şl3�LQ��\�7��ݴ R\����r�u �rr��r� ��q�)�@�1pԽR;�K� ���4�wqwf`���ak�	����=�jV�Ӝ�D��[�gc�FЃ7�|`��nC�ɟUѫ�Y���xm��u�M��).WP>��r���EJyeC���h-7�b�Ea��Cm��F\&Q�~����*��"l�%��$�2Ig�1U�q�*l��D�/�3A7�lE˗��/���(g�M�"� 4����2*�B��yQ8ΤE�*�7�w[�&�5���	I����F"�ر����:O�G�Z+�U%~K���ҼU2�Z�4��+Z��?7 x.�tM�MemOdufn�����af��������ZCy}D�]<�������8q�O��Y_�{��~"9�#y
P�ʤz�tSr�QY�K@e�m6�^�n�n�o���l;vmnW3̐�˃!�_Q��/l�n�����"ļe� ,6�̃��R�5�|\b5���J B�y�jʗX3y�	���l�t0��4�:G����j��0�\{gs�Jg�xH����
���K����L�%�Ӂ'���=!_$d����ӮC/r�y.#�m��^�O�פ���~e�]n�vn��q۔7A���į���yHO[q�gm�;��z�YЪ�2P�/a�P
Fꭩ�����g��O�=��6t47˚DJ-�k��*Iu7�N�Z�����(�g��y>��[�vg%�Dw2�;T�n���:a�u�����w'�����m-�N����c�ȭݭ궻R���i��e��ӣ��CW��2僾;�e�&*��f���ir�� �=�78�P�c�������@D0�-+�P�3��c�J���c�p�+��&ʝѫb�D�Bȅ�GF��4	|��h�Ee�0w0:5}�Bb]p�$ ��E��.k<4 ��X���q�������`R�v����9���.�T�:F�]Jr�-	֓>l#��Kk^�F����8d�'�]Ro���5G���#� �6
���z,���2B�&������j�uƕ����9���,e��� 4�V���Ab/� XA`�$3�sͭf�^����8�z�Mzu"��ZQ���;��ǫC�Hi�y����kO!2��p^хGC"���uQ�]����4���}ti�����V���0Mq�pg��]�r�{�wL�OK�
���7dG�8Y6�9�I^ū�bEU�p�"��ӜQ�C�FX��U?X��ve��>�o��d����TG3�:����(�f5ڵ�����F\$y�|�J'���O��M�)��S�I<X�1;�+j��$��/f�c��A��2�+�M�j�5|oƎ'�WLp8�zF��44a.n;�N�2Y4�~2�Ƕ�*�����l}�s�Yq��er[}�5t��%�b``	��Uhݡ��c旀"]N?c^�w�� ���I��	Y�5��G6 �r�g�����Q�t��3H�S�����_d�,0 L�e��7�D]m�2K[ZZ�e�s����%7��!�l�5 �f�#��~r����^�z��Db���<RZ�(�d h餟+��O>���W0� �I�.@���^>�l��s��@D����C�Hw�9 �G�P
��ׂ-�(��L*Ξ�Oy�����3^Y�eh����_���y��S�m�4�D^,�,F�y��s�?�w苬��=�)��d2ߞQQP�$�y�"��7z��t����ͥ^�[�m���]�aU|Jv^�D�|!+�_��{J��ѝ/�V�{����RQHb&bEK�9	�-C��LR�ZLzQ��L�3u4ؑ5��nDO�HOYL�'/ƛ��l�axw?��=U��P �r)��귶��h�a"ӟN��������)�>?��)��w^~�V�R?�X��
I�<��G�쏾4 ?%D2)�Kww��4&�Ec	�,0�8�k .����$�	���얗�Izh-������ށ(nq����S|lpD�z�y�@�+L	�
h��%]EcG��v0�X�R/���іt�B �ޫ�Z1�a�yΚ|����7ϙ$w�ɥ~��O���lFGd�0ѹ�!�u�bn��"�,���J��N��ƛ��'w��{�c�q\� �a7B!�0A4z^��I��V�U��ck�(/ia	�ݡ��L�>}FޡS'��	�+��Yٍ��Gr���AoR)�+��\(��偋<^ScJls�t��Ί�g��>��dl``�<T�\��bl?tml<{�+�e=�Ω}���я3�=������;kND��]�)�B~�[`�d�hfX"�� ��K�!�~�9�e��;�C��DBp��돳%e��?����
Jlq_��v���<���������,*�ս�E�%�f��u(!�/�3��`4u�$h�u�?�g@��꤯�0��Qs˺���w:y�����2��e�Nsn U�Z�pV�����q{��qa��?��^�7�����P�	���ׂ�vM�XͅEÊZ��ˑ�OSDK�_�ic��0���U,�'�>*�]�m��+�O1`�E���*E�e�@�Q��;>ݸ����U��+dӵQ�x�U]5�a8�����ߒ�\�9oh�wވ��Z���U�&&����N	�)�K�6�N�����NH㮷��l�ȣ칢8k��ZH��5���C�O�q�rd����l^�������"nZJ�૦��;Ҭó�\�V�ss[T�Wؠ�9��5���>q?�Sj��6�u�Z"`�%/qF�r��kF�k��6��fFp�P��ی�{�� �@�� �)~�w<'�R�W�u��;�2�8h.�R�h�dؚJ*4U�-8��kY�r���,kk8��EC���G�%D���Ӏk��yl���zy�����+k���:��I%��K嫪|R�9P��.6��eF���g�!��6�GWU�"Hy�t{�<j�1��o<���������b��֯�#p�J�h�S���*ό���u��klQ��&Q��I�����M�ag�^�!,�Cg:C���s�|"�3L�^0�CKbi�>jY�6T�Y2N
~N	n���S��ӿut�|��B�+N���z}��Ɏ!�z���*)�x���t�B�82���R���Q�bȎ]#zn�jq/�um�VT�	�U	Gp�O�_B�����vtx	G�G�r7J:�B��-ś��ώ��>������#H�����8�q�d����|F2���v�F�N�O@a�G�����*C`�4���}��@����Q�L�����xGE���1ahT{�p�9��Ȧ�k���q�Ob�*Ì`]�s�9�S�k���1�k������>���������m�A&kop9"p#%q0l\�\'ʠ�:��`n=��R�����I��] ����N ���N}0~��.\6q)�iC�L�:���/�B�Ԑ��H�`j�}��쇈���s��-.��|�
 �|�����#!��菭tkW�vq_���>*��^0�HfE&�:Rv����&aD�m%w��㩻(�[��x�7M����m�B��-�<�N?LV5����u��y���{
��L\������q*"I��dU�Z��:4Bh����[������	�4����sN��4��=��!��أ�c�&�q�e%�a���5C�Pi����ځ���!�qvs��t-U�'����Ö����BU��x��3�_>N�`��	�8�95��n�?��M�L����*G�;as�0P'�)�;��̼���:Y�����fopOP�N�c�!�ͯ*����t.B}��+>�%�b�sk��eХz#�U�s���jo�MĽ�p���,�]G��VXݠ��P��m�4��E��a�>�~&�]ƫK������A�!4���m��{j�����s"(`ǡ��N�#z����n�̊��jU  �<m���E݊�3��@�����^a'��{_��n��$��`	��z�������+[{��ai��&���o�����q��ĴHpe�Z���h���<�����yG�1x�~�M�e�d@�xS��� i��[u��v���.�wi�Y �{
��n�7AqG��GAp�\���J��E��Ý�@��{�[�gYa)��ZyUcw�Y���0n��6���W�1�{�J�(��F�%d��K2$�^��Z.��*�� %m��n3����0��d�i���J B~`���K��T�� ����;>�ڵXHrP�]���p��ϝZ13%O(����O]�"�o]�����l����y���b;f�]_6hk)h��&��{F"���/#�t6A"v�]>Vt���:@�T�m'�Bx��^]S�Q �}F=�,v#`�U5F�I!�MQ�T��㼽o��� 1����C	I��-��ڲ�+�y<`�b.D{C*5I��F�G?��Zp�^e5M&��� {0�ʆ�dޟ�}�ʞ���(�K|,,�hxd˸1s���!R���N���*�h!o#��C9=L٪�4���ve����l��/WYH����C�ոˮ�E���I�2��̺�N	�s���2��浂��Gn�*��П���u� ��/µ�%��fX����.�o�c8<�O+H�%�Tv!���j)��qPȰ�$9q�a��_*��#�Bo䄷���]Svl�0߳.�c�&\H��~�A�5�D�ڽ�J�B�==ص��|�D��,��&ylR����!�s>Ih&�(�j���j)�1��?��i1�	�rIs{�p>��}�\�y- S�:�'~eZ��mU-����SI��e�s��*P�c�ML"��V��>���t��IL�:�o#I``W��~�x6�b���@.���0��4�>IG��J�u>S_8��̵���9���́��%�=��9P&�:����A�:��p9�$�`��P*Qqug�'�(�,m�fG$:X������=08ZpB �f��=�@	+���
[Ĉ�M?�"h���¢O�(D�"�/��E\_��弘�.��_���歷��s]������ڤ`�6��z!��)H{%�k��f�]b�E��ө����>�Í��52��i���i`��5F���S��^!@�Fh"�(��n{����ʌ����/H�s-[{3R
������ؓE���0�������)b)�:�=�I��s���`�]��؜t�Ѽ��L��Ff��;74��ʹ���,oUdUIp��ǲäז:?&����\WS���N��,��?9���A�1�no3b��؊�S�@ͣ��^K@��.~ϿO/���õɿ)���9c��=䦞�%�����^M�ǭ���T����\POe��UF�RB<�1��7�2h#KoH�cH�c��]��1[<������1�1\N?��������5��l+��C������m�[����+kC G6,	��e�O2�V�����vz� H1��b`b0*j&v㠕?﹬�ٚ�����EI$-���쓙�X7�F?D�%qJߠ��������Q��EUE����x��|ţ�ۯ3c���e���!��k�aN#v�����5}鎳���K�jq
�pTA��>B��m� ��n�	n�%�[S��s�bo�2����U�-Z�bj�묋����?�8�2b�3�$>�6}��T�����,09�M������m_5|,]����m���I8s�jqM������Njs1赉�s�)�WB�S�	/Mlʫ=�/��Y,ȸ���쒐ɼh+�hZ|"D���$�� 6�\h�#?�m��0i��!��&���"v~�%J�!d�b'BU�db1ć���Fw�&����7G�{!����ٸ�{\���#�Bm�^���g�|��o��z�D����3w3Y�xB��YQ�0,&(њ�S�_۝Iw��:n����].FU֪���Ű3�nM�{_��	�n����c� �O��ET:O�vwm ���w%Ȼ�� �KZ��[g!�HIL��E��� 鈫�ܞ�ӡS�x�g��Yq�@<.v�ݳg3�1��=@��#��r���,='E45� o[��c�7�h�P����y<�����"\��Q��9�mh-��N�s$޽��jf�<Q\�� �Lj]v�[vR�by��uO֝��UB筱4/��s�=j����\����/�)88��HҼp�͊ ��y:ޖ�<K���ܾ��i 
�^��8^Ε����ԍ))�11��`��s^�
�k%���Y�?�+���ழЩ�a�� �챟����+���~X�.��<t��n�y�l/��g�F�M������`�L��ђ���C6�,Eעq�4D|U.�ƖŊ��]x�ѧ��.�b��z��!�9�h����]��j<��=H��G����I��D��aQn3^��\��40�Gv3p|���1s���
oX�I!+u�b<Dr�A�"��oc���n�@��^�7LD/�	uqA��G=B7��o��M;�ָTֱ���QO��[UY�`- ӏI��9O~fz�{�8��5lqt��ye�P��@{��FoN�!��\�F��#���TK��`��F�re^�3Q��Zakmo�?�c�;PS1��	G�� ���3�{k;H1j��������_r���ZB�w�[���
�vM�hM����"����4�Y��I2�*��JB�Ȣ��Gl�f[���9<�Rv����lCXZ���m���t�E��5��v�h��w\��"F�)0��H�h��k�o��ݠ?�Z��سh�Uh�!
I8�D��<�m൴pH��G�csdڋ|�]@l�Mh7d�|"T"K񄣗�D��d~�,��ɜ��)\��g�S:��bx;h5>9�� pѾ����V-��
��c�D���d�������='"ba/�Xv���̃�{�,��Y+�Z��^Bni��
k
�z=.1�?�)CR��P?"�>P�!�+=6^�-V�w&�kh��Z;��])��lA6���m/�����:�£A������!���z��� (�zʩK{ʙ��L4<Yf�iz>��&�>�d�y������4e2�� �q8�)u:�ܿC�)C3O�?����sq�5G���z])wW3�h��U����!OP�-���� �.c�GC��#)D��K�x��?R\�h{ӎs�aw�ͫ�4���L�Bk�-s5ѻ?/
4��9l��kt�vˢ%6��=������WO�kL�6�=�l�%a5����8�٬%���[|�Í,�|�s8������?��i����sr*�1�7�pR�����,m!��GI��.��{��iL��͖���F|n�%W1��������zѽ�o:�B�����"�S��"	�z�q��D���v�·�:,�YV�a2�W�Go�u:��,���3�E>��.�0ċDr+���K���������Zꗗm��0�<V�ѳH�q��e}(K����y��R��cd'�K��5��+/�I�Dh��O�L��� �A3uɩ���
28];.a�w(�O�*ڲ"�/d�Ā3q>�-��cN:�o���
���3�§[H��M���ț�����t����Ag#�i�|�j�b�K�*Gi1!��FD��^d�`<5Sβ٫�|�:nFnB�U�%��M�I��;�O[QS\,	�{6���ิ���^d�b5=����.���1̍�h�Y��_֤�H4xJ�{��
��~���#��� �^#	$P�]���񈺐��3 ���Ќ+��y+��S:��N�t�E�S�V��Y쩤6��-���k�]u��dǴ/����)�(��3Ƭ��c�K'J��l���ʴ��r�2N}�е���+�x��^�k�8A�K%֓>~!y�RY׺��
ͦA�j*+��}4�ݴ���S9v�}*�ߢ�n�W5y�N0𼌬�Iٔ?�H�pQ,54~n���j�|H�*vC�C}W>������HXI�伬p�L/�MB?nU����l��3s�ъV܉�4@����W��GY.����{� �D��^S͔"�_?��غ=��=l�x���⼰������㐦ɺ��[|��ݴ)+~#�m�e�8���B`�^��9��*r��W^���h�\9�ٱ?��{N"�8�[?�|l�3�Oc@`_@Ҟ.�1��y��YBPUW%h��/���E���|��"�Q���c��ddа-y�"V���<f,�[�OJ��aT�;l���i�X���c���e���u$�UC3@ζ_v�� �y��D�,�K�ך�D�r��= ݷo�<�笔��I��h�k���DE�j��y�[�:�	�~[鶳 ^p)�Hx�Ң�~=�:?�ᅅs���t�	a�
E!Zd��wQ��z���q�h$I����H�O^� Oy.c�.�z�$ᑄ �(�x՗��ݔ��˙	^e�����w�$�#�St@��|��X,��0���ᣪ����96[���t.��>�]b%����p^3"}b��~���C�n,�h�=���ErE�
�)�w���.L570{R�����a���?[�v�� e��
]`�@[�h�&2\?��,a��0�®����� B�����+Q��^�)N� Afr3E|N����}T
+�{ry �xz���T)���D����n�v�U�d=�shAt�:�I�]��ߑ_:�J)�X���}p<���x�O�@j�n��_)�����"1�; �VR��s�������Q痵yQ
0e��L��l[|O(��_vu�R�Zj�7а:�8�5!��cU�}�S�o)�?81�	�5�?)륫Q��?��XlW�V�b.�B֥�^t͞�Ȯ��T��y9�_�c�/��N#\�S��:];�r�+[[��!y�E�%sMVD�`�T����Ůk�b2$yL[b8�V��T��i'��ʾ`ߍ�t_b�~�����'i�x�@�v��i��{"�bY�|��Y��VC$������V�h���x�_h]��ɏ����I�"�v���"�}Z� ������1�%W�l�By7�F�=��D�^&�窱���:��i�������	�㺛���:!�w!�9�Sa���M��&s�R�YК�D���q�Uꖳ�ġ����v�3]A�`զ�S뿆|1�C�:?w�ߦ��VITuT�(-c���ުK%��]ֳuv2C*)YC��������(���+oΞG�?�!2�ˬd���'x+��q�g���;Ϩ<&�Wx�s�/�s��:��>^��7�Ɨ{E��ʈޥ�5>��B�� 3��Ⱥ�h�*T|gX ��7���Zp��⚴r	���SN�ўBr���!V����E}U�0_�=h(o)p����η�`�ZVֹ���h�q�aLw�������lD�X���X-��O~E�'-�y#�i�Ą��`����cܲ�S#�dA0���d�?h5�3�$&�ϙ9�}�f�O`Jb��n/�&2�=(�l��)8���n�K�O���&րF�4��<6_&���F R�wVV(n�r�+���O�I�8��i>[K9c��3�i.���&�;�l6�5v�o3�w�ةN�Q��Jۨ�����XӎX'�b*Z��M~�[�K����O�!�4�Oky0J�D �j��x$�=�����+�0�f���n��>o�`�t��3�ˏE.���]��o;�t�wc�2IF��'�@M�k/A�w �!�-�y�k%5��5�2��<�5��_�z �bl�7�O�vp#l
�NR��Fz9ߍ�3A4Œ)9(j��Ǘ�o��4�ܚ�|7��X�����Ԃi�e�������!�`�U�*X��v��!@�/����Ηc<�kU�88g��!ވZ;�R>-aRo�]�`�RX*4&�Dǳ��D�@�8�$�B�����M�K�y�E<�|��E��&�w�Q���'/��w�N�+��ۊ�Ӑ�쁽uoH��KÔ��v2����=�$0����;�ť���`ړ���2յ�WM9}�Iz"�g]&�,�`�����y�0�=�3��z=�vbv��T闟!�W8IW�)��3 ��r~l�K�*Kw�+ݡ8�X�FE��ƥ�͐�J�9�L�_�t�&U�#�EJ}��2]���Z0,�)����u�5���:�D���a��²�D���-v���3��؈�J�������DN�)����mv�W�o�W{�k��S���&���|o��=��s��X����q��7�=>��(~lIF���H�BZ��x'����} ��$_S����Ua�h�8���V��A@�+l�>�u�U�FJ����D�ˌ��KWa�o���������]g�@��	�,�듧��տ�Z������b�f-�&��	��4��k)n�9�����)34L�W"����Y�D��Z��{^;��~��Ɨ���v��&ov� ��H(j`�Gm��������yi��A���M2-��Mr��j�4��M�nw�Mi�te媔�0h:�����I:���"6$В|��M�i��K�)���y���W_�Y�Y��!��q��H�F&��/ ����ɢ�90�A�(S�z�����}�o<6Ȳ!��G���Ds{� ��zk��&�z�xTϒ��K���S������]��)C�+��ܝ�fʐ��ۄ1�$0�E"�Q��\�M��.\{��7����W+�C�!ͅfu�����F&��)�0pg�e�a"J;s�,��(j'��Y� ��� �Y;E��)�N�Ӛ���LKt��. ;�V2(cZP�uN���61�B�dj#U�����v���-���)�)�g`�j��X_�q���@7���X��[��.�B�յ�<�Lrm(z:Y|䛲�����P�����H�t}(���{Q�lGb%���7��_=����Ds8R���)�gZ*!?�B��m�J���L�V�m��`���^Q�Sn��g��B!ab7�﨨#��|�-AA�2�1J��@�f8zpp8�ص2��h5���I��@�t�eXW�Df[�P��Yw�̴��ڲ��a;��D�Ѳp�����O ��k	��*pǎ%�3e.���Z�ym�_���N���ś��<lҒp�_@����X!��~4(�H�$��m����|7 ԏ��K�;������߃�s��u��(-�����;�l�u\ϲ��d�-���b�Nv�9ԫ6��OO�#q���Tk�;6�E�Ǧ�`ʚ���(;E?(z�N�M����RV�A�\��bl��)��y#�:
n�C��r*V7��
��k����2��Ovs�ن�?0����&�$�0�I�&�0�U�����Ǧ	qa߼���\T���o�|�0`/3C���Xt�rכũ�$���k�t~i�D�8�*%�|���uS���ꎽnQ��U`''tO0 �0�am|�2]�Xs>2]0'W��/�佇�޹yfg}���@��w_�)��������q��2���팮�Ѡ��["x贘j�G̕�o���'�h�?��� �B�ٙo�3N�T��?Y�����,
���|��aP��>>�u�y[�:�#h4C�S�"H�f��c5�I/�p9b彞vl�����%���$L��B��bU���)��de%K%P�s�n���q�>����#4=>Y�-V�n��|B�ͳ޻c�,��7��F��W��&1Xʳ~������3Q��r�2^�\��2P�#���qL��R0leP:���:�?R�G�b<�Q	���"�H�y!��C������񜖔gY)N~뎗߷f-}Psn�����.�Z����;�m7e�5�؋��ú�O�İ�2�}似�+�'a&�w�u���bHB>�W���K�G�m���ւ��A��V���r���������ȡ�}QDl�?�(n�
,0�s�fO�K����OP4�'ޫ����#$GX�5�f.Z9��#1Xr3͊�3�;H��*�����:'�i�Iwf~�z�hJwg�	��%.㒺UT|?ފ�e�bmw}�(�Bq�n�}ɕ�_{ʹ�l{�ƴ#S�fs��W��\����=�٢H����&��#�W<I����c͸�;� +
�ՄU��W�j��� ��q��}��k�]�|�i~�Q��4��a@\ɳir��/�.h\�!��!��t�c�:Q�̂c�|�=�s�b<�Wq��8��D��C�/��C%4�/49o,5�Ns{P	]����llN8� اne9֬{�V�#����1��áт?�u�ժ��	m��uԬ���]��VX��D��o��G�d%f��E�G�"'�N�h��T�~�up\ᘲ���XV Ϊ&�+y3���ypЬ(�g��ʔ���ݒ*�Ll?S�fb�t�W.t�+nK��a�uC����,�!�x���>�z�k~5���aV"#8�RqZ�4��b�CU�:����� ��&�ǈS��&)B��#��ф�2/"zxm��Tj����婘h��k���;=[{��j�`�8�W�妙�Ґ�,�|J��0��ԩ�cY�#�b�m������c����Y�Z������քUKS5�QL��O`���.ǧF�;9ے��՚��ߛ��uϋ�sL"8��gA*_;F�(e�\������{��O6�׬mhj����?��
n�寥����Qa��~@�*�۲�@�%�9p~�X�:��s��KR'��g����糷FY�.����1�g^0�X���إ�e���rك�I�4�Ǫ2��*yٱ��e�N�`jO0�\�8��&��F5d
_�2�E�^�z�m���Zyo	Z��u�LaR����.1�m";�Űn�b��Y��8K��u�,P�\������B��a�wY?U��w���)�d�nN�[q��K�*�Իl�@vUYA��YԲ�+�����i���M6�zN�-d��C�ǀ�ެZ�cXD��<M�����wFG���ӿA�V� L�z�����D�^�3�~D�ˁFO�2yg��d?��.��@&8�*�mo���S���-0({�$D��,Oǲ��I!QD�rk�hY��h�Ë�>��΢� !|�^ˀ٤}�,�+��C?��6�ˣ�^�Ƴ@Y�v��8ڷ��^��:2�������}Y֭@?x�,��)��.��5| �sˣ�\\������Z>���x�M���/�L�*���&6��tJ�7g����~���P�hb�,��z�=A,8�6��9\�N'FQX,Ѭ� ?��	�z�u�^��I������<&���h<�<�_�Lf23쫂���ϡs��$^0���~1���z(����8���+^�Z(/�f;���6��~�1/ԷzL5L�
���١�p������\£ض��إ��a�Wf�fH�@��|iV�������f<�K\�Q��䗣�y�&n8����xx8�UJs6y��Ln}�!���V��P��ɓ��W�r2�
�6�l����[�l����O��	��H���K҂@�
��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�����uK~YSokj�&�9ȼ�P������şd�rU�gb�nEg��e��`�"9H�bLr?\��F����H�;�&Emv1u����7�^K��1�u�ڜ
�4y��s�n��S/�������s��ai�T�V�6�H.�X��x�O���H��s&��,Na��d�V9���|���:����amB�Rp�� 5����$��+h Ϗ�&�-�.�~�
P��X�Y��+�}`������9�~�m���_Pآ�{�����W� �j?��1��M2)s�?�Ng��Ї���B�F�]�;�y�	-:a>v�'�"ܸ�##7�밼����di���7�m��o�a&������Mk�[���c|F�v'�-��,j5bu�����\�;a�Wg1��d�-m�T��M�{�a��d�/��%���<��#��`��������;C��~�70��\M[�[��E���S�A���'�^�*���+��С#H�ȕ��v�.R��aZ������Db�#�29DfE,��P��L1N��4�k�qgT��@�@��9U�Pp���Unc���(oͮ�ь�v8�@F�n���^ZQ2x]]ۆ���S���~d��"�#v�ǖt�2/�0l����'�˜��ro5	��m�̏N4�Z=At�ѵDr!ݨӿ��}��M/�127;���^��#��<���"<�T+#NZ,���*߹��4����L5�6�5�Ob�eR�n���N��ͱ��]��t��Z���*ˇ(�C���QV�?^�~���gAA��^��K�'��L}���n���aGM�c��휯S��r?�W���ۏ�>+.M lƮĽ;��Y���&���Z�bT��8�Ń���I����:[��/�_�l�W�+ٰh+���E��ԩT]�;n^�&o�r�|�*)j���#�`##7�n�+����ȈP1؜�K����t�ă> �#���.Of�tX=�w�t2�v��$�0�Y>��b�K���'�C!/�+L ˋ�f��N00�+ͷ��
*[����-ȯsp�A,���2���\%*j��8���ߏ�<.=܁}�j�*B7?Ől��EeCB� -�m�0ˢ��s�)��|��RR�'��MPt��qfu3�v�o���곭q˴�:�-J�0��f�/s�U�2Ճ㒓���L�1m7�ڒ��J��!��6h�@j�������֣�����)N������SP� �p���]�>�rO���{3�#&0�]��H�Ϧ��i�#�\��M�b�z:�َ�됓g��k|���і��h���Ej�p��6�с�ё�m��(&�(p�:X����Aw�d�읓�7q~�"��J��2����$�����q~E[���$>~�C="]���ý%� R���DcTv��GU��A���t�VGJ�~�*o�+�ڄ��N���P�ZX�Y��XhjW�x%+��,��d�[vw_׻�b!�P,����~J$GTw[�sx�"�돛do����2��/M���֒��'=.vhi �Ǔ�1�\�X��>IO���3B�}Q�����@K���h��5u���M3l��r浣�r�ކ��.Z����C��?B�H�1��dz�
�I�~h/��T9��T�w�u�}=��A���N(���uH�W;�������R"��H�o9�{����#{�<��� �׼�s�u� �`R��T=��iW[u2e_8I!R���{.�-�#8�*�W�mJ���S�{���~��j�BwA$����`:o��W:��m�N�MX7l�yFji�9��,O�ꞙ�a�&lJ�։���Ǝ`�-UJ^l��y�j}2�N�Glt��E,��`�\���T?��	�DnȘ/1-�h}\��y
�R���h�P���]��,���b��6c����W0=�V�W�k�w����RD�����7�6�i"��ܻV���Mr2�ro���$��4���9�v3L���Q%\�Ma�8��BZ��dĞ��t���`rc�b��ܩK\K���Vj���Z�F?J�8��{�3Uv����m����x�CE\}.��*��y��o��t�?]�E�f������ǹp�,�}cr�j��ڕ"#[�4-)��'/�s�l��M�G�l���� Z��|䉿+�4�̽Y�%w�L8�E]���?n�u D��+sZʝ���G��{���@�$�+���������e�Uf� ��k*Ę���P&T_ܭ}⩯�L�F����U�[�~<{��>l?��Y�8���A o��D\]I;S�U�r+XI'�.G`��,�;�遠N,��͙q�qƉT�h\�&�!��Tְ��n������s�%���`�-�[��Ŝ�&*@կ��=��<
�d��IMYj���"����x�qh���ﴕ('�	�b��R���7��\o�x�����p
Y��\��@�qXc�~��v��"����V��Dm�Ҙ�PPR���*�e_��=20@�~$k�?��p���z�l�촀��e<4��<�u��o���6[�-�b >���UYK�FM��Q�R��h;v���0�@������7�����l�ȳ4���g����sdm�

���dkxw�iI*9<�G	$zE�<?9��
5��@R;B^�*mf��QS"�����A��ƥ����q:`Й��,�'�~{s�R���e�F�}�����=�S]��@P����gJ
Ŏ:�l 2�� ��;�A�|])��Q�|��G�ݿ~��7�����b���)CJ�(Vқ&r��ȕ��5��k\�v� ��𱴳��������S\�C}��c^���bqքl��=���	K�,��ɂ�9r)=��S*�^Y�.��_����$����ϕu��A�ph���ĸןV�ݜ��lы�??��fb��=����vF1}��?�f�w�=[���گ^/���[,��7]�F���¯���t�A[�@g�*ς�-��މ:a���B�2�M�U��Kz����">��Xa�^�P3�� S�49S2��(���(�(�j] ʜ����Q<'�o������d�r� �jq�r��2M��Ţ[���^t���LNk�$�꾍�#SB�p����@9�4,��"X�*lT~�0�w��p�;(������T"C�	�M��T�;�;���nc'Z�0��;Sβ��5��x5�������V*7��;*�G�����
�������@�]"�qNz��J?T�QU�i{ �'~�'_�]a��Lo�@�i�Al2�i.ީ�8�8I_����tJ���B�p���$��r]�"{����B�gyU��+��-��Ë�z����mۿҷ$�V��O��?iusk>���x���g�c��ެOa�x����s�~���=Ɏ����?h�2���*� ;��G\(�>t��y�zi雛I�������W�~�D��2%��VH8�0��{���93Mc|�ӟ"�N�<\{ ��:�yɿ�$P:�����:�9kl�UKem�%`��iQ�7�7� ��?�㣌O�hBE�Ǟ�����0DQ�	0N	��"��ߎ�*ګ��+�H�v�K��ғ8ş�Y" �{ʓ���1��J��r�X�c t�b�^{S����W�x�o�AJ����P��E�`�ͅ;��D�M0=jx����'(J�6�t���v��p֭�����Z�����>��\?|���5�G>�G����<�*OX��0�p%��� �I�I��aa����h�`�ƛgP�7s~�[8dP�ϯ��S����)Z����s���J��#D��[P�2Ot�W�N�[�s~Cs.�*�ƃ�foLh�եz�e�5ȅ��i1�����<�{g��,|g.%����wM �$��#��Z��~�r��g���U����_ٰߩ{��9��S���vAuʫ�Z�>�JT`���VYi/��S��_�u��zw�qP�m%��c^@ڌ�L[`9Z�t�(�I�I�v���~T5*����B��+���;��]��<M��#ұ�F�E��
f(l ��y06b�\i\fVC ����rUT���R��,����eP�Bw�L�,�zö
e�s��WsQ��9M��]:Uz5�=��g��:}ϩ��o��X�j�z��tD`%;�^�\�S9����:����"�F@J4Wڸ�ݽ$dQy	<	��ga��J����R(����%��*��*�"�َoC�80z2�+�OrZ��W���Ju7����uh�2|�l(=��*R��`�D�ď�CJ�+]�$V�R�Kg�/E�N��{�Pq_үW��yP)��W�#������Ѷ�]�H �]��X7��=���@?����	�%"bk�M	�
���{��0.�8�-��J�j��]��$ua`	F��i#A.'j����%��K�����+<�\��:���K�Q���V����ߔ�$�ShH��7���,�GzVo�1��m#0���1_�o4f��I��7��t�	�-�u{��=��s��(p&=����]��!��v��%�g��TX0���p�����q����q����+|X��<Dw"��k������Cm���W�l���C!�t�
��~��g�Y|J*]��!�ycoԚ
ʠ�9��Et�f��" P�
��û���*C�����y�A�%����������T�1@���g����+s����f72,F/~�Ǖ➰�>�2�#*�nTt�w	�$���F��"�e��6W��)�����om���Co�ԉ����X��!����;"$������|���"p���?�N��GV
@�FYY�MM�8��?��4OEz�p�E�h��l��\r����G��
�1D!�U�n�r����L��E��� ���䗝rU�g&wY⎅���.�eg7,-� ��jX�ZҔ��B�����_W�(���F����� 9]����n�����O��
���>��
x�nS�-9�J����|-�YCA"��,~gX��b�~��Qo=M���OD����3kI`�G�s�o4E
ʪ�Y0��<?����d3�+���)gW�Ml���f�TV�������:��m����B�r[��o/�ȩ��ii!�ȴ��M}dA�����&�&�2F����"y??�Q�t.+A��%�򏋢��"$9or=T{��>.�m�� �;E* ���<�X�q��m����bn����ƨըc��=Φ�a�����v�����d%U�@�`�����k��LQ)���!��=�A23Θ���6u��f��8/)�Z`�/N\ l���zi��"-��u�j\�% ^jB��n��/�zͮdV3�����A���3��|E,C��MM�?�G�F�}~PT��e8�T6R[���V�>�0�����.� O���rh��
?鐉����I�95��R�`!��9��Z4&X_��ӨM�*i�Gvi���3G���LՎD١�72&N��Q~y<@3���qMa�f�Y��kF��K׮��I@v��Pi�A�:��"^�X���x�4|�Ĭ���I-��\��Z�s�V�Tk'��&�^q1'�I堻���Ȇ]#�d�SF��(�ɨ�����HR[0<C9�a-��0�� TO��aG���zB�t�R�Q852e��YY�6��l���:y_j��&�P4+���]dc���Q�ٞ�����N��w.�%$9�®-H�%�t(d�l1kI����eU2�%�ii�c��w�,'n��m۲�J�m���Kq�Ϟ �3�P��7N!�B����K��9��'�0�q��,�^�I������|0��N�v��	%O`Q$�e�Z����UT�Ťr��HW�E_k�4�4�-�a�}���&�n�ʋ��&���G��4��D���*s��(m�fJ���(�Y +�c*��L��:�Y"��o�^���!\O���R\��"
�`-���x�����]�p ���Sy%�	��\��>/�&o�pX '�G&aYe"�e�S��@,A�O��+~Ds}��t���{�����%��e��$'+F�h:T7��.����Rpf_�7V��;��#�h�c���P�1�?�"9����%�qW���X����<�=��&���}�i�X�?i�ņkS�}��v�sȜ�o�:�b��:�F42i�!d�dl �/���/�L�00Cb(K���y�0��b,��,f�	U(�$�?s�d�}m���T�����@�Kp�����?S+���Q�����V���"	E}{��d�_����'q�j�G�o���F��"^B9��3H��	�ߒW�Q:�g�V�R��E	��$FEe�]�W�M��I+}��n��q�e��m}�T^PRF=�'�f�*���2[�h2���=V�S�3ͬd*:{�<�2c��wRЖ�s�]r��w19B�/S@K�?&:��/Z��@9Ys�N應\	�YL }y%�^O�-sC��pGv�ă�r$Q �ň���2l�z�/ik9�n��X��VL�Ƭ1NK�a#UW�;���LxĮ�f������Ԟ��Ŷ�����������]�E�u����ual�~Wc1*�9�֚M[��FYl-.�G�ݵ������O����oh61L��=&2�O�v�����9Cꆟ�������v�[�`ww`�W�F�;�p��d&2����� ��g;�����$,�{	�P�/{�rB�%�6#��mBx�E+���g�qW;G��V$�)���Ѷ��l�uu�^���z�����"^�
������?=���]"29�j24�뱐���e���`�0]��G���g?���cV��Ȍ\���U�3��TR�\�:��L(���y˦.ѷh,E;?�O�_�1�%��qm�P6�w�~��`fA��к_o.�S�V#����R=�$h���ĬN��dM�n����-��U/)dDITA*�b� ���@ă�5�yS���X������Ӯ���6#�C�.�?�I��C�ƈ��bf2�ЊN�Nk�dc�a��%��sO�gzڛg��J�f.�Y��pF���p9iL�/h;������}�V�`��"u��tw5�_9�wjセ��DG,B�������땫�H��r��-H�/?ބ�D"��[��ŝ��y��b^�����dz�T&�sW��7�;��� ��5�� ��n�[x����])h�+�&�n]&���[	m�Z��B���Ɋ�A�[Yn����$��c����Aߘ�����C�G~C�e8��#"#�׻Aw�rb�,��{:��Jz�ԿJ�L�4��Y��q�ޅ�-I����)��/��� L�)�����1�V�$|&t86 ۫���u��y��P��[
14��^��6E����%k�c�Hյ0���~�V��7v8�8�:�����};��!��&���˷�����u��x�ʮ|kLeL+n<m����,$v�
Xg(j���nO���K󗊩���<:��,�K�6U��/'_�41!���=��v���C<�^ˇ����/e����{���[O$�踐���y](��}�����]q�͸��0�z��X��<�g�Co���P�@z I�i��`���߼�=1C���W�)��}]���ʾ�����T��-(bc�f8}��a�=\3|E�zY<1���֝2�M�:���ؕ�2	}T�g�YП���]�f���i��i5��<�$!-����C)E�t�
��ד(�_M'?v� �=<*"�C}�Fk��]4�&�Ca
�~f�࿅��C!�����b�~��L�jʸ������ҩ�T�Ʈ�P	?�t��:�A�>t�p��L��}1}jH�����_�w�يD�5/Tdݑ���#���Z�0+�B�ڳX^#ǣ�3�[�HX�����]���I��HCl�1O�L�T�B=����J�0Ja�-�4ቇ����7z��D}.�\;`Z/p4q��:e{O�VP��PP�+��٨�C~q��,ӵ�-d��8�C��q��S �; m�:�f�9�:^��|n�H{�HoH�����%�I��Gф	+�e:�9x<�4IL1�����2����<�d��BH�Uo�.ي��0��jy��䧃�bn䙎5�<�1�anS�ڭa�}3SS��s3Vj��m���.t�+%�AȔ%]�y~��C���Q�E"ΡC�:� �K�J��Aj_���C�>I~��_�n�i���g��:n��ߔ�f�܀ݞ>��Sp
�}�fR���5�e�k�.>����Y"�5�uY}.�Ҿ(�'����:i���Q�]JM���j�O�ّ%T;�BKLj=���]��C`�	r�C�y^7��N,{YQt���dDY,��:E��0N�J�ca�G��g7	 Z���"w4���� �4�b�`����A)�qw�j�@�f&�:�m!\Ia�������5> ԫ�G��zn�L����ӝP�j���p��OIY����VVr������rA	+B/�|�B�u�7���o�$�l%�v�+ڀ~�3�6�?���rf�Єmu	=��f��p�w'%�6�� g���.���p~�S���c�6ǈ��u$�xőϣ��iQ���o��U�����Jhr2�I�i�\3��Қa�@�B�c?K���;Q��S6�$����[:�(֪����3��貳 ���je&����G���Ȁc�Byjj��x����a�t!�����E��H�K"��b�q�!�&�g�ʶ�\�η����֠�'�4��� �5�b��q�NT%*�n�a�H����H��v檎��
����я���z����b�e܇Q?�z���q��?�����-�7����yW��m�7-�w�)z[������"ӻJ%2�D��K0�P�<&v�z,��o/�nx����*�F���įʋl�=�K0 ��^��1�u�J��,1UC�NaQ�KG�[�	!��5�����e?�b��ȭ�9��N]�ؘ���mt'�!�30�.�[xe0A7���P��ݹn
N�A�J��R�{\(nC~�(����� �ZCL�N6�&�;ރ|��7�e��v��br(N�^k�%����Q����?��z��DoJL��l.��b��mŠ�֞��\�Q��h����l�9��^"H.T���"�&s`�+�=��Y<��Azu�eW�\�k�>��	�`�n�J!�s^4��9$-_ލn�n��'����q�0�J����l�p3�d���
�﯁�
|�x�4���J�)3y1��6VT4�P(��*M�xJ�$�*(Y#�jCgѐ�Yrߡ'$Խ�R�W����(�g� =��!e���sw�����iH��`�?�;�I)(�M�,u���� ���CN�8{�����#�$�8"���$�-%?ۃ��]��r(S!�����c	)�|�ޅ�I�~Pݚp.�0|RSҦ_�´J�g���/#�E(��y﬛�5�o��oܫ������o>�/w��Wp��%=*�����	�&�ο!�o�z�	ց�������-�[�nK�x��% ����\4M�:��l�9�\ы�'����vC��L����#Kp
���ٍ��8�}u�^�tMn_�H6�_j(���,�*�KOI6#��$����K_ΩzB$F*���o�W��GIK�$��a�ZxS�tۧ�Tձ(w��xim3��pэ�)�>�9'Cq=*�V|�%hT�H
���vQ����q^aP��p|���!K�vŴz�u������P�)=�&'.�8Ǖ�4�S��$Em�����bo��`{����q�����lS>���`����-U�t�PZF8f.r�8�Yn����b�8���,@sG��+�AS�cL/�̬�&:������t�k3�2 �s����m�>�/n2ql]z�ʘ�pb�+�迄G�9-g���.���[��,H�1
���uXQ�I��E}���jTn��B��2J���L���4���uL�WmT*P ��H�o%��r��n��?X��5g�X�͂�D�,Y/���b'�~��ᣢ��yu�ɘ窨[G�;1j��B�c��R�"�K�CU]��OgT�،V��+����q^Y��uA�@Z英��!�J
������̼r[~\����7a���߫F_��M=�3T��z�\��H�@�5�\0܈�q۩�ɗ�#�����Taݝ~6#���'2���_��cd�5t� �_W*�E�/�lr�tƝ<5@=ro�x`�F�(fc�	��¸Z�@ؚ�#�����T�8���IK��z����+�`�8��K|H2�?�a �YH�c�ߠ��,�4�\��1�_u��s��w/����ŏZ��b\MH5.(��k" �+�V}�D���v���-������.�9�hq�+G�_������w�%���g����2�K̿���v�j��c���"w!Ƒ�ǅ~L�H��9XY
��[�A-�VV��e���gͨ��|"����,%1W��;J7u8��v��4�bvk]�+�m�:�����;8���a�б��1HԺ��~���!cx|T�lk�Gg��ym�Kt(Du����.yOҡL�ģ i�\�e'�/��1�%�Q�B�,��L�v�X�0�(���U��
{䁟��%���{ɱ`?\���o�t(��B�I(v�t��Y�����;�-�L�W������;����b�Q%�ۿ���s9�j)3s 1�����m�)��	��Ja��7:_%+D�>���B.z׷E��ᬨ�;qE��R�Um>dv�e�>))f��1a�)��2S��$����Y\ch�5u�읭=�$�%.)Ne�1��L̸k�, P���L�r:��s����kϥ?l�Fj ��1��]]u(���7���^!�ݦJ	�п�lz02�|���1T�}���%���;ڒ.v���۶	`�?�8������*�P���َ��bD�n����XK�#�U��w&��������G	y9X���?�9�ʅ��0�� k���a��@J�� ELP����������=��n��dT,��B��Y���>@�NY�UYdE�����4g��W��R���2�d�WȎ݇C�R��KYN z�x�������'���3��N&Ŵ�����1�
�� ߨx��J�0��>�p���9��Y��W�k��p]'�^Jys�(4�NRY�����uə��d_���o8���瘯.t��� ��~�NuW����]I�0,_���h�G�CV�e�F����.y¹��w�D�+��z�$]�b�$5 d�q��|�G��.M-�C��!JU��C3��Wn���Ԋ6�d�c�����X������&"��cm��YL���J:�D���&��f����VUEt�-v��P�ݷ��1 ��պ2c�����O�tN�|t��,����o�&��*^u9�WJ��U�
�?��_a�.	��wPNN��4m5Z���͐i��v�y<��'�n�T	/acz�=S$Wf��Q��2<͚�'(�޴�+��SB*����X��J�<uw�|�P�	�7O�����	����g+"�*4�a���v�Ɂ�$ؙ��^����wL��Ӱ�dՎ��$�,wJ�J�yr�n�&u �C-�C�^I�r�goeo_���]R�+Gb�d�F�9˖������݉)��39RvQ��#�6I���a�ړQ����K}�],Ͻ!k8L�j�$>�U�mg>�"MV$e�s�hD�t���B�̅�DA�X.��ۈ��<{8Lqe���!����~w��c����]�Z���D��"U޺sjHY�]����꿨����cq賬��Ѯ�otv��y�JN��K����� �wSR!L����$�c�q�;��0�����U�`d��a�K?��{C�Lq�e��3M�)�K��w�
��z�#i@}�nP$�&]9q����.��C�k�¡g�����%�=��j������}��"��� ��v~�]>�qST�����)��q���l
�@��p�Z����d�s��T�U��k���@���0s��[׃�p����h�9��f�GJ���`SƦ+˱	��5�x�NM�x*J����!w$�����R`#Fuq�Fo�@R��q`����DX��Q[�Q*1���fм3���.@ղ�F�e�S֪��Z���-1u_r�4�Jº�0��u�1���y��Yl%jg���A�i�R�V�I+F���p&@��>�j_Z�ܧU������hӇBi�
�9z��ܚ$��!3V�LފA��e�)�6����չ���8T`�V����z3Q]�Q#�|h%c_"8�-��f�wZ��Y�5tx=���=�C��C����J ��	�x�Sf�׆ӧ�k:NGů��E�d�?��)�6��-�����T����J���"Ш��,�ҕ7
K�D��n��6%�B�URv�Z�E1%>��q��_ ��\�h����>d��IXϣ��A>�(&)p̆&�D��<-���N(vp��[X\썳����dM��L�����كҪ�=]�Й�Qh(M����~:��]��_���X5
;���2�<ɘU%���{�J�v�R1߷g�H-���NO��&�1����Iq����ѿ��kJ[�YI��2A���)��|=�+�����e�)�>���������Jv�\������"S*Z���Y�6TvN>�slT`_>"�L� ��xU�e� +�oS|����yj�����E��EF���J4@e���b��CI����y�06�%"�Z�t�J(�Y�����FQr�b�m��J����np(١J�����/ݢ�1a����ZQ�jQ}�c��ڽ�l����'�������x��N�>Mn�T{�@OC�%\7���ICD�6�bE�f�v�,]�$��'9S}�'wB b|�l�©K�W��j#�|s7��y�M����o��?#]M̤x䓾�Y�A+^��#d���#����?XW�A���Lhc乛�0X�WD7"��$���v9�tz>q�>#֠��@���i���@�g��U��O�uz��&���^ �ZG�7�C
Qr��5��-g��z�,x�{��k��PK�q���8:��Fʼ@M�M@���q���GWm��:$��	�ɿ� ��>U���zu �씀1N�����?-T���@��c:��@f�N!�Y��*j[\>�r���c$���G�a[���QR8�֨�e�PpC��8_O����P��A��:$4��D��)bS�S�r�Q�qE1КVDͱ��,�@h��s���@�^�[+�/�n��$z�d�-C�[��ݯ߫���amȍ���j "P���Qe�4��&\w"&��v���C������}0_P` Á�\��/��*\q���i�]}4�'����9�E�D���.<Ω雑�������K�y}@��>4�_�r�9�`$eB�ƣ���$[�R��c�srA�i�߲����0p"��n�R;��@��;@��Jq7r�C���H���(�諬���݁Ĳ��*z5[�4����oxn�n��W�-4�1��[5|]�������x��3�|�$�K9���T/��	
���1�Oy�E6h�
(=ȭ�3p�Yݮ�B
A T��G:8Jk7��>Hk�J�Ei6B%!�[}�[�څ�{�yW��^�A T�xp��?�NR&��{���V{��|��&T�i��q�x�#8L�L}�Wo�:��SK=� ,��]~�����?������O?�YY�n�����3_ �bh|0��Ҳ��r
��I�����AS���A]�L	Fe�,����M�y�*����!�p���m��o�i~�砺�g��SEF�k�א��Ƌ�����pJ�F8 ��l�-�E�}�� 3��Y����u�%���_��>����Җ#���7s�=F�̤�2�1��̽�I��~��w|J�uŚ�<m�f'>I\�p�2�+2�$(���5m=���$G}\���=��(�����	~����Wt(+H^n* O��g5ڶ����h};C�l�tىC�o������8���͔G��&��n�t�?i�D��W���QG�z����H������^�x>{>��چF�P�|6��*d�����dpĔ﷟��CTP2~X�Wh�޲�{��,�^k"�Ja~�2h�'��rت�����W��$�;;���)/��2��=�>�G 'I#_ؿV�����'��L,L����񝚢�/���?tY���^.,
�nK�B@k����UaS6�t4��q��^�����\�y�B���J�*;�-�-�El�5���̂M��q�����B6� ̃O�,���S�pA0s��i�Q��m�<�-,�����@�	H����R�4�P�m��=�X"O��:��"H�2Ԥ��E�\�v�'T����G��p��#�QYU��Q�=�p���Ų��S"�g���m�nr"��h�����x�wr/��H�*��7v"�gQ�ٿ�U
D�����Q��Zs���f�o����J%l@�3��{�̸|a߁@o��Z2�<IWo�=.�E�Ga]�Y2۶��ȋ5���Κ�4���J��ŃI�%�T�l ��,h����9Z�/L��_M���G�XP�kW_�W0��:DVɋz�t42��3n~�6�H�BhM�	�ZX�mK��u
j�[mݞFm��3�ƀ{.�V�@XPA9C���`2�B�'�D����cW���U���dE�h^�uV���%؝��/��E�j�����U��n�V.}��[MR�S#,��l;�$'�}�Th���\B�Cd�a�� �\�D�}�,�4�՝����A��l���]�}zO�!���)��r�n(za<6=�ds�ŝ�@D���wU5ɼ�(���cQ}�E�?��~��Ma���w�nI����OW�}OZ��2��Q����N� -0Lk��Gk=5����$�G�)F���C�A��E��4	��<�OӡΤ>vKjV!� ms�h$�:��W/�զ:9&b�J0$2��1�-^�U�"o��`#���7��ņ���|g�/a�����K�	i��{{-l�j�W�E��W���.-��\��0��e\�; }S'5��5�������l�H�Վ���:���������x���y�?����ǻ��C��][��� ����� ��٥VR��L��m"�7p2�ܔ�NT$���F�,�ee��LT����#��󎆘Ex�
gx��t�:��k�n��A���d�N9�[Zd���j�� ƬMAu����Ue.�
�?�V�Tà��l�A{�r�kF�
�6Q��~�ti�'�&�#��h���Z��1y��>��� �<F�v�!� Q�\�D^�</f�~�������`�˫L�l(v���u-�O�1��� �,DNZ�� �����*�����*3'X
3z}�gՏD�)z Obu�V�\BkJ��4��j�]TOHb]t����L�"^��s|�%d��t-3�(�u��=�T��'���g�gP�J�|���m)Yu�^K�;Π{����h}��dg�j9���̕�>iT�J�`�,�.׆����-ⅻ�C�4�P]{:O4YV~�u��a*�O����P�uּy�y�^��<;+.X{�Б�ZB�����`�q	��Ӌ���j�:�V�)Y��Ix4�煬GS����CK��I$�nȽG�sÐ��0͓��ifҵ����hC�ħ��s��� V�}�J�L%#P}�T=㓓5�E�`ߒEh,��9����܏�,,ˈS�Z���_���c�%&~�M7����O'���\��[:_(�l�؆�q�L�$|�;���<GU������
�D��a�Ӝ�R\/ǹ��C3����l��2���Z��Gf7m��N1��,mCƟn�8[��F��!�3�Ȓ�^SѶso���kA��zZ�����hg�j��v1�պM��zl�����G�ӆ�	e���J�5CK�7\Uu�i�y��ف	�\�G�o�-:����q��,�m[,�j�����;5��vt�{L�c\0�~�8��l'���y#�]�����RC�r���p�R��>D����f/.�{�ռ<q���w5��uHvXtQnq�<�lf�c^V�;m�����bXv�gu@�.Ry��
�����i|��fM%h��#&SR����gͭ�<�+�3-�!��R��w����k��1���
���Ewmgi`}�	�e������<�w�FG��5xJ��~�jO7�g��q8IL���\) @7;[�f?�4 �X�]]_W�ef�]���1�-���)}��ȺR���J���,J�}~��ݠ�<Λ��W݊�㕔~��B��CU��j��|�����E҄�TF��>簵�+h����@F��a�C�D�d�6�d����l"�����L
�A�u���@�&^�s����9,py�;�y���'9M�y2��X]sbCQQʽ�T��<q�ᶨ]�|���g��"F!��nDnߢ�]z�N�j�!�N,?ƷI�.|���.˾����B|Y�Z�&�{�1��6�h�K�<�ܰJ��=7j��Y�ŋ��*��zb=]�1C��P����8�@#?
'T�U<�pȂ�Y�#�0�L�(�q���~І�6��t6D����Z��D�Ǥ�v�4���p��Ņ�0߆�i�I�� �_Zt������d�H�⫪�g��B<���Q0��c�Z	d���.E{r����_k����V#1j�L���z�)�[��\  �O���U��Թ���uHC���4i �o
du{�%8���U�`������=�dl�!�1"'���И?��� ��e�|��FF�x};O�+me����-�d�c���F��R�����I_L4.�H���l�ٴ#��!��G�aդ�Dz� ��-i�H?"�����F�����g��3Ig����+l#:�6����'א�QD�Ն� %���r%�Y^�E�)~L;>����=�\f�s�ؔx���q�9^�V
O��˲B�L��󋾼M ��'�^F����~�^�2aV��b`�����L=�ƻ1�9��k���%�\��z��h���oz;��߉l���Vj��JNҺ�c�q����+��F&�����߼|��G=�C��p������!L��:k�o��sN=a��)m�bS�1[�����c=��"�~��;p���C�q�$�� !��G9Ghvo����"�O�2ς-�=`�2c�3�#��bKJ&�bb����?�1���B�sz�Ԅ(V��3?�!~*<؟&]NMz8�Ӵ�b�O��������Dѱ��՜T}��1���έf�w��OLRdud[�T6���Ԩ�7ī�_���:��i�������k��>�.�P������Yf�<��;���5ȊT�@�F�T�٥x��G�>����ZQ�����$�3�)�=.SR`h#��r�g��Zߜ��i�v�{Y�3��;���u����6&����/�u!�����܈�`w�M�CO��Ng!MT��_o}Ti�T8^������R�	�0at�E϶�}8����ò�!��y�L�~=�����@� �%54�����]��H����6��;ȩP�0E��7����f%;�~�� ?�U{A���
�Ň!�ˍ�\W)��7A���[<��cPm���6�o�[0��t�|�HD��G��(���KH���b�wu���s�N!�sֿЏ��l���;��T�)���5 #�w)v	{�ȣ��W�(������a��z��^�e�9��J&�} ����::�hv����=�t:�.��b:��[�X�e�&(�x�n)DY�̃���� ���:h���O0<��^6ף̥�+u:Hi�X��X�gf�t)������Ք�xT@य़��Oz� u�1��R���9>g�.��P��]�E�Ī�8<�H��9��VK�B���`q�#TD����!�r�V��������0O����V�H�R8)G�M�(�rނX��s=O �k�(U�Px:E�:����޺'�Gg�_�� 搉��^xl���������]�/O�3�x�6��31	��$тn����w	8?�ZG&�G�_�o�W����4^��
����D?�5~�k���S7%�$��X�WG�g�o(�U�[^�So�c��='sc��~5o�Q�1�-�"��f��U�վ���R�9��2�@�`�J��o&�Y�b#�u�K��凔ne�nluvr-*��-5����K^:��p��0|3B��{�}�9��ٸ��M���q:��`��ZC�T�QhX:�L��Op���|�bq�Fs�i��+���� w<'�D�u�3#G1W���ǃE�d`T^}[w�f-�0HpR��ϳ�������i���Po��� ֬0R1ҍ%� �M��}'����/I���E�IA�Hrj_��FN$bi����Z�[s�䚧���c6�J/�[>��Ȫ�H;�L�W�&�{�/D�Yv�Ӛ P5����w�F�k�h��!~\�x�}�I��?�~R,B��o��nU�R��I�-�:�״Ц;fIPd90�W,i���"�o���L&�����C�B0)�O4���J�>�$+AֿJ�W1a40����#>����VX�n>2 l��(f��*`PM����{�D��p���6�J�^~���$5k�b?!})\�脮l�5���mVԄV�A8���E׌���[lk�>����޸u\���L���o)
M���mie�8���,�H�y����[7�z�b�=bG������,T�,�D��i����ἾƁ�">C��:�va_�X���:��k��t��n�g�X�%9�r�6��a�%�r�'��}��Hz���[�;,tj�O�j���n����%��h����衱�����ww6s���4���	W~�����}�|E����5���5w����)���r̘����k�.|��ی)��@g�L���Z^�� !�Q�c�A��k�?�����=k6mf�1�b\O�w�ޅ�v����I�N�������a��?]W1&b�l�K�Q��2#:_AY|\���q��a�#O���22S�_2�C��޾��Hh���@�����;�v�^j7��ʟ(��EmjNΏV�}��Z�Q��\uu�ueF�!k���=�g+x�Cb��
y��!N{^�D|Z��P2t:�*��T{v�+#ٗ�U���f���j����0��T�
������T�.P"��������9�ʖ�y��eCh.B[��S�ī{9�|7�\&s���~��zWM���Q���u�78��[S��
�0��;����Z#4�0�;�sw0��G�eN���,^<�sx�Cn�uW	3d:T�P�Rb�����s��éF�f0��L�)�^-�x� �x��,+�3qHe�f�J<t+;��④��(9�o�q��/�\��xXd]nՅċ�z}v%��R�0�I������!Ǆ���� )��_��|�	_(c��t�B�w���B�`Q|[�B�j�۱�w8�-��Nۥ�-�61`t��i}�ܴ.O $�d$�/���b�Gc����,���f��h
v70/Nl`��y��+�:υ�����+����\��,��,��Ƹ�wt����H��K�òV�5���2�@A��~�dW�W�y�vS6mk�hC�I�-�s�$¦ɽ,ԶE�|iG�̓߰a����S]�lW-��(�{\h�5�|�`����j�=>C� ����UN�w��B�~�,U�I˳�nmK$�xپ���e4n%p6V��6��h/u�������@���N�HR9��O9Q�"���Z#�.� �o�T�Z��̪��?�'p�V��L�h�Umb,-N�*��g�l�P��9�-(]lF�$l���vu��ʫ��L�x����k�a�����?�20��N��0,S7���+6��4�JML�C�S�%�ʹ��o�x:�PD���x�ߨ`N�����GUQ�V�I��z��ժz��vu�&ά���T�0�9���w�dB_֒��;H��=�=�:b	���(L��oa�x��� ݏ��9m����w ���{.�f��[A�ۜ{�3�1�l�:-}Ԕ]���UO6�a-�C�1:�{����l�����&���%�Z#s���DZ�]�24���$��%�	^-@Qu8iO^��8�gmI�N�T��<'M�9�"��}���xwLP��ڸ������.����6����B���n�BTH����
Ew�%㏪ͥ��-Lѻt	��%
ؓ�U\j���C�Z ����pݧ<M�K��s�7뢉Z}�-︅կy�M�f�
o��%��"�N�-��_�m^߱޻��C~W��#vo�ؐ ���\�9[��ʎ�G$���ӎ"�V��ψ�gs4�.S��Qw��a����o�ý�V����smy�{��b�j������}���3kmϙ���+L#�A�}�~>klrt��u��$����U�x�[���;�wbZ�lm�	pϵu}w�,Dg{����`�U�*���c�eL��3�>B�ا��s.�Wc�	x�ꥫ*
�(�-ps�i�{$��c����h��y�m�":� �+!�L�F[,�%�{�vG��"2���h�;�m�;��0
ld�m�u�d�t�������{S���n`{&��b�
�>دS��i�b���?'\���124���p|��w���=y"<ljecD�~ԍ���ܓ�n@+���J�'��fV���~\�0{��$�>雊]߃�5�� �����:�Ӑ��g�������z��?�۶���"�S)�@���}G��E&��c����p��}H;IF4���01�R�b���W��q_�H2���*�QWG~����ˋG(�[�4�r��gp �~�}Wq]��^��AC�B]��E�!X�w��A�X��a+�#@�&�Z?ѿzڂl�����	���n\��F���}Q�dn:_�m���'�/�^��JCEa	��=�ېi	:��W����-�"�Z`��v���8vm��a����g=�\��ȟp!���,d��X�Q���y��܂Ч7"�����K_)��\�^�_�0��E�ִB�3�膄�~���7w�@>�>�T�� jNP�r
X,��B��c�e�
��=D �;V!Fh
�ڰ��$��%*wCWX����.����W�_�ؼ}MA�[��ۺ�1lu�=����O�@���n�#sqV��_uH�NA�Ǡ��������M[n�~��l�ˁ����5����<mR(��{�9��g� ��N����9�F>;�JU��;�h����>R��o���SN� b_��.�&�6������W���n32�Hk�\��(\s�b�kf{��֗��]"i��*q��250����|;%���d���&|~.��FNv�"��Q�_��ލ*�l�h�G������'�F:%0㠵�~j�W���;��L���\}�D�0H><kM���)r,fQ�<t��	�`���^� �34 ��ɯ( �Ut9Yl��� ���?E0x�ND��q�ӟ�
���CT5�F��)d�늙=��v(d���A]ky��c\�C2��"F�Nv��^���'��ϳ?r-���H��w�w���B��k�^��-�"(ty+�؝��Yw��M}�(�~g������1Ҍ��R�����r�nM�N�q22�A���ƛ�(S8��R�2���� ]�����3T���2@�"c-ü ��O����8>�+L�9,'�!2�O�d��8�i�?����Q>m#z���x��D��E��nQ@N�����!�B�̀C]��L���v�m�@~H�y1��@
�S��+��d��������j�~��bgsqsY���?�ԝ�@�6t:~$5j��MȪ�� %�z��R~ɩ)و.C�{o�+�ђ/��Ԥ`�X"n��i��)D ������eyY���77���z7�j:�>?�x���!X������Y	�v�̷��'׃䯱�j1d��s���Q}��l�
�n�
���"g��p}%@}�=�ڮ,�E늗 8��yv�]�����x�N�Jab@m�RCn�P��3g�Bm
�\���"ٵƅ���X������j��3H#!;Ѷx8zR�f�&��u:��N��#"y}��
��f�c�u}�U�^yEޙ������Z���RvB�T��VpҎF��Ε8�ڿ$�j!+�6J�n� �}��cM��'�=�p���f�u�����d/��h5��Y�p�pRe��e������S/ǱU�����8ج�bp�	���e͎�!''T�?\Rx[�.�ֻ~`�9`܎a�.v=�|�&��t �Ddl��g�$����{��� ����79R�e@���HR�5>����*|��8q������A�$�*�,��alB�z���%���)*y[Mx��ts���1���]��jɎ�y=�չ�Wp��]���e��D��N���㙄�Y��%�<�E�^fd�9�,\Z�TUk��Td�b�E���v���L���);���B�Y���m1|�Aō�RL�đ%uQi5�'KA��	��s�T^��ĥ������:T��ի�ǹ��;��=��+6F�J�c�6L��j`Ơ�3J�^�B�U���ږ>���bFl�N��N�z�U�Z�9!���zL��Ҷ!��?�2u�F:�"I�<A�i�a��1A#�ֿ��,�\5j���xŒ�.qZя �����0p�{��(�aWd���i+I��dii㋊���\�Yi^!Z��
��M�/Ė�ρ�wߒ�i����$��/4�W��bc×�ހ�n*T�$�%)�xA�N�S�cB��ʔ54wIo���l�Af��Ҭ[�rȴL��uxL��jO:��<B�Y��R�\�
����t3`���E�hJ7�eđ�ƪ�^��+k���<|:�7�z�>1 5}�?F%�c:���Zm<���>�`��i?���HcC�.n��\c�q��yB^�1>,&ЕlwH��J�W�����/�+�_P�?3Ǧ-���w�'3����j_�n���3Ґ�, C�Q����+��k�����_��̅��Q�����J#��c�����<	^ϽTz���>!~P.�lt�6\R2F�[��Ki��JF���Qi,���S;~�y��I^D��L �I���4�0Р-<���i�c������
W`�6�����w����R��I�S���	�Ϭ�k�@0��g^Vi���n'��% ����]t��c�s�W���DÂ�Gm��!L�s�o�h���F@�&�(*�sq+%I���z$|��hC�;+Ũ����J@�	Æ�3d��#t"���d��[�h-��)m8�]��a:�x�@���5��+�(�O��V�3g�Ěm��6���ow֊���J�&|D���ŋ7N�w���<���vR{��qn+i���n(2�&�v<'J����v5�����t�� <D3��+PHؔL�ES>�7���+n����Uޏ��*r��k�~"N^�*��4P�w�RI���I�(�� ̓����N9��1�k�+i��.�I��"cd0�z�ѱ�$x�g�J:��xPiatҰ�`@sm�j��Ư�:_�����TB:߬���&*����{��س,1i�9U�,$��ΐ����唭yu
(��m��>�s����T�B~.17/��zl��0����!HU?�77�P�tֺ����9�	5�!�nA%]������g0��
�ӱ�~>�l+��^z���%��̶���������֎��,�QֲAK2�_�}���@��̼�Q$ȗ~\"��ϰY+�~�Y	��i���x}���8��,�	�O6\�1E�R����o��4\�T�����:������ݚZ
��5O����7�H.�g�I��&�]�d��3M9(�JT��I�-�uS������9��a�z]5�`�m9���#��{$(�O�>������;[��ӝ�*��{�q�s�8�F�&}�5	WH�~��1^��U�=�����=Cנ����g$EW��W<� ��i���K8xs��z��2ol����ݏ-�R��g,����3l����L�
��1#��mˡ���N=g�v�P�ԥ�;�V��
#6�44"0��>�|P%GQm�3��v�Ԣ�r� �C' x��?���dk�ڳu���/�*���@i/.��=�;ژ�y��b�e&�Nָ;�ۯ�+U|�� ��@G�R�k��s�Z�~��_��j������`x�K�;�k�ʘ%Y$CB�q���"Ź�EY�{��kPɎ��@�[���¶���B�����B?�e�,��:�?WʦD*�'k������a?��QX���w�Pw��{��j��ҵus� 9^S���I!�<b�v��_��ja_w)��s�P3�b["N�΋Cmm.�&*��#D� mf�9/Ѭ?v��Ec2+LǕ�3)�_�HYP�X	�7���1p��Yg��јQE�d!�,<倮�C��A�d�<믶�S�d�kT.�-���Lt�Bi\��G�eB�������<�P��ᙻ��moփ��'0��r�DmzZ��/B��dO�I`���rƓ0�$Y����<�؉����A^�«X���tv��:���#i�t�!V��gs(�{����
o���5���F�+'��.>D�	�^����Y�E�	i�%v���Y�G�4�VxF�CF����\p�H���_pz�@!h#�	�z�7�eq�uI��nj�lIP	ǓV����R��~q�t�He"T6c$L���� ���.����n[{�x�X2L�ϛ�u>�ĵ��:�����~<�B����bede�O�+�{�U4�R�\���gx���s:���s��*9j��}ⱍ�!UE,�X@�U���[A�������q 1 Hr����m1 j�MCO6"fX�oO1[f���uo�� �X;�ݗ��^���}��V���MR�<��@���V7+��i�[�1�:������Ro�g�^|�R�t1�W?�0[w�g!\ݎ$�0F�q(�Eo44ovd��ȧ��p��O�&M���yH�����X�z���vY�-{�1��)A�l(��5Ug�2<qA�oF贏�.
v�U�G/_�p�]�Ǣ��!�=��jt�syw����!��(�pW\�P��;y*�4 �
{+�Z�h? c�.��V�	i�?�UB9��N�S����~q;@��!�3��
�F�\�mS�����;]�70
�.�G/�)��a%��j4�Gy#��\0+��������mPQ�
X�h�sܴ*���{��$����ܚޜx�qH�T��E�nS��Χ��Y��%�8+�:Wy��� a�η���GƗ�f�J?��q&�L����<����P�y�Ȭ����<gtw�V�#��Z� ys��&*�l���B_���Z/���(72�w�������Ϸ^$��������`�p=�J�oow���r*�Ӌb�&�3��Ԧ.�$jMr#��(wW�Jm:u>��^���:�%Af�����ŏ�0��;>h�s]��+��r]W�*>;X>ڝ���!�G5�����瓗��oY:�GD��ژ0�F����f�[�%�itLGv�#1�@�w�3��X���A�v-�����7w��"�����t5\�O�3i�*��S��X	�`
�8�1;Mv���6�3?���PЈ��R!�h��{0�RU:�$JO�?��j(L�{(�۟ӇH�����X�� �(/�> ��ݚV1�����a�<�9Ff�c�'�=��4���N�A�A������THy��#�N���� ���5�������6�HpNG���DIIR���Џ�~ 	�����^�}w\N�m�_��559����1�l��7�f㺀�����7�z� �:���"R�{���35���:y��C�-�g |*�w�Hm�9Rgh]R{��V�����x����1_�V<�!���i<�W٠4�/�a�%�,�(ijど,�ϥ�w��l��3w�����\6:�|N�m�����$<�Q�w���4�G����!�c�:�T0姤��I�������#8Ȯ0�4�JL�[���!�ӄ�y��JS��}�
���V뢠CT.&a?��}\�Fl��C�?�Qw�3��s�Q@��$KP�r�H��$���.�n֫�ԧSO�)�:�����<�F���=��@$)us,- ��l���b\�G֮��CI�������Ε���[6�ZH<�����v�ͼ�S_:�*Qߒz���%z`t��D��W	���t!
�^V�k�m�h�͗��+��������?x7�)�/P���@z�Z��:�%�������XfZ���\P1@�dI@$A����$�)�����aF�#t�ԱHC��3� ��9��:9����������s����z��e�g&t�ef����d+'��3G7�7�L1OL��|��|_�i�%W��\���TV-�.uj�N�O��r<��Y�d8
��9�˙��Q�w���.?.��zܽ��0_��K,i������%=�`$,�����5��@J�d'�I9o�T��B�{E�����>ܬ}��m�ѩ3ta2+�ğ�+"��K�����Vh��{�u�t��GN^�Eݢ}T��L�
����5N@e�MZf��������x���x_;�0Zi}'��7�� <�XkZ%�BU%��n<#����S�xe�3���6�{g����l��� Cm;9���m)I*?l:b�ͩK,l�X~�&��1״��))�!Q"���w�At��o�g�f�So�֡�U�I�$�.�Q��}�ƛ{?lRǤb���H�hÌ%	t��U
���~Xe�9qi�E��M��5����f�����?E��nmf>���
���aӎ�� �������7 �G�4xf�%�Ii]tN�V�c�yVya�6�DԞ����\ޓ�kc,��aL�K�GOʐ���[�l��7���z�*uf��\���i=O ��j8�>���҇˨}^�'�u�FYI��M�Kj���)���!0��+����x��%}�49Ǽ�{��G(8�����u�����~�!EX�8;��6n�ʱ.��������2����~���$��5ݰ�"ږ���F�SN|x��½W�<1�,�5�����%aYRJ��ya��÷}CU�g��\��ԣSב�|��2����L�,�Ak�y,%���ǥ��PśA�ϱ�����e��!�<Z�:BݞX{��N{���h�V[w���Fۋ������Z;î�Ls�l�j�<��h�����5���8�y*).���1�[�
J"#��#	�n[ȂV�|�l�����<�6�\lk���T�1�D�5N{F2���AKZ~�k4���S>���M��DT	y�M�P�Z�UV�w�4�\��2y��-��R�o��!OF=����Ӭ��8Ȥ]��������gӱ���� ��.���B�F$��yf4���ZQ�8�lP}��M�^�iRsu˹������Կ�g��9n��q���������@=�QK�T�;I��a�5���7��X���Ǚ�����pR�[M�H�qL"��̥�p,e�m���~�-0�n�n6>���e�%�@�=6�G� �PSK��pr�
j�
61ʗ�������U��v����n�ȡ԰���U(��
ӗ%�����l�O䶨pp�m7w'�ֈT�G��D�n�g�w�h�+&-&v�iC��վ7�~�kO6��Œ��Z7-� �UW�<@�Ϣ��ك�&$�2�L�����ę��-%s�Z�
Ѷ�{�;jB+v�� `6A�V��3Ҹp~�����3}�R��L�ռ�fE�`
�������iir:%)�c͢���K�ѕb_oJn�X��'s��Р���?�Y	�p-�����Ɍs��o
	�4�D)���<,v>^�rjS�o<�K֝Y%�*���z7����^�����˾��Ϲ֫t<{�D8iw<[�Ѩ{R
�f����7P��ۦ<	���~��h�ٳ(��Jbgr����Jr��s��9��4�x�_���yL�ю���]]�&��Бr������L�0��q�/�K�ܦ���9�VT�G�ҹ��� ���lv�馧�ٻ�FxИ@���u�'���pA��~\U�rc�AD�nrCn�t]��C<V���Q�}�,nI�������z�:��O,��;]�;W��/@��c��u{���N, z���U�\I����	��j��(�(�� kz$�\�_<���6�)8PO+�%��N�_�޺���9 ~�ee���;��ڴ�����:nP̻FAKV���~R��;_Ϝ��m�;yÕ�%6�W��6k߫T��:�<�亚�7� (�'�(�!"��!cM ������1u�A�W����9*�w,��U:gQSc6������̵b�5N�~#�;)\��/Np]V+�p�.G�x'�P����v�i���xc��a
���q��d���.��s�����-�ٲ�$u)�j��]J����:$��c��l�_T��O�2 8�9��k�.�q��|���''�q��3���O#L&$7&Э<��A�>��by��e:�F���ۗ?�2袧Rܛ�Ȼm�l�[�����R;��|z�z㟢��vK�a�(2o���V1��_2�J���ɞ: �Cw?�J�D$��|�`�J!��M�Z3����2�����350���!ʣ�ir-�u,o�(�ѭ?-ĤK�S4�%W�dl�'�:ȥ��v��;�@�N^���=\އE���������=V(r���P/o?�$Lz(:��q�Р��	�]3��i���IщqB�}D&\������]x8.K>ʲ���ҙ;Mֵ�#.b嫳�YM���zY��R�o���즞>=�Y����T������,	�&�|��o��MΛ�g
fO06����	})��	g�ߵO��+�K���u��!@��o���EkA������; Y��)[�2�{K0C^(���亾"c_vB�!��p�`�V���E`�f(	�O��2۞�~p��� �[�q輕�&	�����޽�R����;Cֲ��]p����r+���������H����alAq�%�ǒ.Y�P�#I�>�)�|�SQ$���1�Y���^!�*c���;Bbb{��W�.~��4�H�����2B��&����E���E�x�`?��~�֨Yp*�@=���ý�tY�����f}2�����ϖTY5�~*�\� I7���Sp;��-D��,ʀn�-o"�q N ����k�t&~|m�>=|�T�5^����s	��X%��=Sq��h��7IH���q���
�p�ba=xS�ݴ�EC+��\M��z��o7�[(��V?�R�D*���d�.͞�{LZ��Z��õG��x�Ƣ/��Pq3�À�w�v�(��B��\k)G~H�V��Ļ��ۧ�����z��!�,�F������ͪ�.JѴ},�@�O��p$&�O;s���Loj���J�Fd�x�)����MX#$��k#���"����S�0I�H���a�e|������\��wJ9F@籶P��!�{`� 3��� '7R�m�@?�tO���ʛ�et^���H�1ꝷ�B�n�t�����mşbI%�ؚ �47 a+�o"�
��
X�L$��"C�t�$���+8Yi�8Ԛ!�V{�\��l�q[�/X74%䭴�f�9���|7����7Y���臊��Q�/�a��zzA&����O��L����cq����n@���?=���uՆ�,�XU�9����^�d�3�H��}�1	���<�Fg�݀��OG�
W��� ���z;�B�t��1�z>����X'ҷ���2������m���\iK��5l�;I���a��M��bj��AZ�- �dmsu<zw�>x�����g=�'�{�:��x��q_#Ώ>C��w��c�ˑL6��BǛ� ���B�8�ς �c}ܞ��"�M��&f�h��>�M�	�Q���{���
N����MͶ���q�Ԥ{���{�YX]־��|��s����+��e� �pڦ��
�<&'T����%I�h ¡HY!_d�$EW��eL�I�?vp��'W3W�&��X�%�M*��=�����zP�]H\+��΃ y�5:]�.~�o7�=��-���&B�C�@l֛�5�X�n�:Y��w�b`o��}�,�D�z�QD�ɺ�����Ơ��x�Y)v�EX����X�v�ro̞�hhr�M�f�]%�+L�Bw�%�e�itQr=z,n�ƿ��_c�jg��4��|~}T�>Q4�͠ܟ� f4��/"�WXK���E������|�+�*:�H��;�R@?(X@]�*��c譸���zBt�Xvb��
�ߡ�F�ZQ6Y�J4$�g ��ޤ8h̨ۡ4@7�'S�Y��Wmեb\e�}�Jӌ��)a4�������XT<Ep���{����T�&�����o/t����8�������E�~h~&I��۷>J�p*���N ����G$Fί���b�R�
AB'�FB�����S��U�k_É\�nUI�O�Y�"��s9�:_)�e6�{����ϙ9g��|�gσ���� v�M�v@zY�D��3�'ŀ����$nZ#6ሼ����Z�ւ�b�%�*ɽ���d<�ޒ�Jؠ>�G� <������:G��QD��M}��D�f��t1�}�JG�8�ae�M��땃��{	+�LBm|<�?]��8�2�|�v���+t�C��X퀎\�?�n�p�74i�}��W�����������AS1�I��ʑ!�O=�S�T�`�ʾ/��V�x��ї�j���:��J��������HYT3n[�jڔ�55�1n\k���Տ�ĺ�/ߡ�zF���K���l,���i���ﴧ^��@���G���ӭy:h�oZ��m�1ȿ���&��;xz�QI�<��C��1��vb��Q�֌K;ƚſ�F�*2���ĩ�d�A�#3�Cs���>�%�`l,"�5��f�CAx�a
'�Q)��4���Ϧ�%��miSA����𪚽Noy�z%/�"��efݥ[��zJ�W���A_�ߌ�le.��g�ua��i$w]zpm��?A0�`.�1:�L�m�?�3�1	[�t~��9D ��6B��M���l)�}-��}X-��I�w��`r/�pg�y o4�S��djN��ə�޵Ǽ=��6���h�C<�����`^�pȘ��(p�b������!$�[��� �;-ٓ�:b�v��נ0k��bU�����+ȓ��D���߅1�0�T��}��5i�hNMK�E�-/1d��Ĕ�ًqX�-��ȃ�JU�>8S���5%�f@�\�4DY��T�2��^����Y>Ѵ��{ou��~�F����\���lj�:�!���i��3��f��fH�׽SmvY�-H\Ϸ�p!�H�����	��92�=s���e���@)Q2��~�Vu���x�{NC�{���|��!(���<U"0���� �£����n��¸�,���cl���v����a���܅f��Be�8昶 ������4���-���tG�|��C�(}�]~�w��؃U+5q�:�W)���bj��)s*���d/���+��w�¼�n�~��}Yi�]}�k�u����8��5A��N���1]s�1��2v��b�{!$PKvN�(�ܥ�5C�;�^q��,E�����Ĭ��v*�����2�ϻK����J����&)�>j�#��:�E�6B��z�gf�Ѵr��-���9�N�;�A_pR�?�Gs+�K4��s��L^:��/�J�Jϐ����J�تj�b��8Y�c�	�<�O����D�ⵥ�$|��N�Y�iW&���W���:(�c���������z��h	�(��<�4��~�D0]��� 3�X�5�p�"S�:̬v��(�q�%vJk1��t:��u4�[���N��J���Oޡu��X� ��#�ܮ�������!)J�g?�
*��n�r�|-��� cz
�f׆���zl���\�t9��n���v!�0��#�@jl�K�!sĊXfnԙH�8�G@6��w�d*ׄ�E��sS��,���W�[}�r��VVP��W��<K���=I">���a�G>}�lv��X���'�����eVc:��_i�o��]y��@>�5��_a��� ���xJ���h�!h��E����R1G+l��V��W
d~7�Z#�:�lBB��Kd[����.�:����k��oZY篿��;�sR��OD@)�:2y�ȇ_|st��ī�}�<�D`��W���y�nH��dJ��_ȶ�i�/�W��{Y�����&xҺ�D�4�U{��{�����^?�ڈ�|'�m.qn�vr��1�s�,��d�,0\Cw Y�; ��jG7�����d�@}�<Fƻ�~�xvn����B\�n��<�<?��*�H�$D��j�o�`[YR�;L���W88�q��O���?&�P�Mv{��:�}���u[�J]�2��[�ZƤ����#Ӂ��n������Iik h<K�&i~/;� V��Z��BW����T�j�MĬ�����la�8&x%I��/$�s�l(��7����^�DY�kÞW�J ']��p��)�D���o��V����D�M�n
:N���:2��y
�Pb��� h �*�I�v���|�܆7x�M0o$�<��P�P�HC �5�u��e� $Sx�~M�3Nl��0u��� j�� "�^.q�K\YA�qv���:�����D}�Y��Ӏ��W7�����!�w��N�I�a�{Χ��Vy{ۄ��R	��!3ѣK��d?`/�Bh�!KaY��G(O{0(�_��뺌�˷��V�Y�a1'~��=L�:�u���w#����~�b!����%Dcaٍl�X|�'�\/��[í-�!W�5 ��nut>�5=@���+�w�!]��>����~ض�����l��k�O��q��05L��駎�M Hma��T.(�|��$��n׆@�<�x�
�+��:4_R�w?�H�*�p5F�9�rb�v�1©$�o��N��w K�9�ˡW�$</���Jp��n������kN��z����b�RO]�=I^h�WQ��2t��A. ��=���u�� ھ;KI�#1i7�h� {��p��-����"{
TD{wWi|/��p5�F�λ�3;7���AL�\���B�h�`����1���bcw�������Y*a�y�V���S�fL��͊L6Y�� �5;����8���0*L�4�-��Cdă�..ǖ�@J����X��^dv'c0��<�J}L�omܵz��[�H$=���A����:L��e��/���Ww�;:]�/Z�����gxn	Yư#[ѐ27S�v�D�DL�hLV��`:oX5z96`�>��F>�!f�(��y�-�������
� �z��n���+� ���H#����s�
�����[�H5N욣�q���xؚ���(�W7 (?eh����<�c�+3�T���b+)p�-A����Jxƞ��ݓۡ��<��d��VL������/�!�ܨi��8ٶ�rd�Q�:WL]¸��n{ 5*���>2�M�gZ����y�69�
��[τ4ȕ����O\WZz;Bi:����Y��a�f��d�R�R��n�:���l$x�8���1W�.����N$C�OKb���)�������[�!� 
�Ĉ��.-�ư�J�S闓��x/�/�+/����i�l]�7� ���Q��j�T�	��7���_��<���?�`��~V���**.��/�kL��V�x�j�.D�)V�<!�����薛�J��P��fL�T��y��L> '��x�V����O�s��ۤ�\�[Cg����;��]2�m�^�v��w��K4����4�F">*�ڄ=���M-�>�Ȭ��K�	X���~)0D���Jq���o82=��
 IpG�.cx��hX����I01�S�!��
�� G��hT�����"ۭo��V� v�^-�O�-T�|X��h۔�+�컂W����大F���O)���31��y���y�dMɓ\K:Y ǀhD��_	l ��F�H�Z��N�>�l�s�ذҙ�¼�_g}�L�$��6^\鱊|�A_�u���<�A�4a�P��Z�,�p�{>}����z��7rJ���	�����L��v��,���.c�$c���ڿ���p�o��jiXI�����vkjz�2h'�8�zMz���ٮ�o��{��^s �ځ�K��-J����*a�=�>�辂U����/`��'��3�P`dO��W
g�@G����;?�
s�ۖ:����)���U<Dߖ�4s�|����4�\�P�ڟ�E�&��+fTS6��@2D�xq�b�����>M�'��|�������c����'XA��M�dpV�w�tv�aX����7��췩�.��_r��M��	.]��4Ψ���������nH4�U9F�Tg�hi���kѬ
��D�Zǝ T5�Q�Aۄp+������B|�����1���/Q�p�����>�K�
d��>�
.��r>���C}x�WY�{�NNI�L�������⠈�B币�s\��ǔW��O��y�܊��ud���ސ�?�]�
~��$�����)e��f����wO>2����p��Y�<52ޙl��͹�u��wl>�1�)�˯��1��8D����P7P�Ls`�@���H�p��fi[�Wa�6��y�_�?u����Z��{li+�:�;���j9�^E��i!B������y��K8(v��h?�(���5c��7^�):#�W^��=Ȇ��A`6�����q��6��S��j��������՚Nr�6~c�zH����4%���xS&"�:��:2i��玈�6��sFn8��{ \����a���_���4���6�zw&g��}	���[�i�^�u����.Y<+���U+?B1P����'��5�����&��sl��Y0?�w,�H�� �E��Q�XAvf�|)]��jqQ�Ay�CNj;�}b>������ty0͏,!��}��eb��y��u�R��o\t�u�������߅�*ٌ ���������{�z�c/�(#9�ОU4�á��G�P������`ɿ:�������O�C�=�̖����LS����
�A�A�B!�v�W��ы�h�Z͔X�uH�w�k����\(�
�;E�p�uV�� ����}A��&�#��x�Lǋ��, �w��=��b����!m��YD/�IK�?����d�h;�yh��&,�Q~��2y�A\�:���F���q
cX����sRJ����}��z��I�(q �a7�w�J?DB���Cȱq-�U�-dV��E���#4\�0��<{��`��1�l�j�����r$1�̍U����mŴ��Q� |�8�BSGj�n�|8u��7#I�r���ӥ:<a�#��Z=b� `�՗�
39�J��nZ�h�9۱��K�b�~�VW��ZԼ��
��[3�bօۆ'����ym��,'i�p��R��	nddhd��������h"��]U7��P%(_������194��oƽ�0T����;y�J�,(�
ֶ����_���rt*"/͞E�0�-�+,��Q�ggǀH���o�fb�3m�k޳Ƽ!��J��S����e�6�ܵ�[���� �,�,��|ѫ؜��GX���1+k������p����?YU�}e�߁vM3�E��>��CT�HhI�_{'��{��)n=?Arf)mj���㬑�G�nߣ͌RF���kt�4�=�g��"�i�:�׾[l0j�;	N+����Eᕘ�|�����i�5�B�ƱM���/�&�� �z����	"B];�
���~a���V, b,{K�?��`o�Pb��Ur�ì�Z��?~�j�`��9BzH�$�n�[<��`���SN���f7�8z��n�����>��Ʒ��83�����>�����>�Fo׏��B0� qݔ"��	?s�i��F�w�Ӧ��һu,��̵�F�������M0����G�G?tq�7�]|�ᰘ��ii	Яbz��{�?%K1*N2Z&�`�xt�}m8��F�a�6,���j���l�am9dm"ƷJBs[(�ʑ�/����_IA?���8wV�L�I½p0h?� ��&&��4Ⲑ��+~
$�����,�oC���y�!�nf�ډ�}�<��c�u�������p$;&�j5���Q�mL�t�N�uyCW�x��j�7H�/G�sG��@�Cg\S�$YX�Gi}
�ЖQ�甋 Ƕ{Мj_�� ȣ��X'�h���]n�Ҥ�q� �M�E��(}Y��X=�a0j��1]�SC	C����/�1R,\�;�:l<=Ʈ�Fm�06_� d^���N�������`FB�y�����Rh���i�,����42b��r�c�$ZQ���ǎP�T���<!��8%����P�~jW�lf|}Ȼ��a{Cc ��!Q��{a��e�9/E����~��-ѧݵ��w�%��E��:8�	�J��#�ًX^�����0�)��}
�P���V׹��Y\몸3@����	gG1�$^����Jw��O6�	�mΪ�0x�A~B��7QP�0��Yc���ъ�tY� U�.��q�:�ʵϒo����<��x�NdFኃ�Z���O�UԞ�o�8 ���?A6({���|Y;ɞÁm���֞�q���QGJ[ Y��z��/w폸���e-�#�)���C�*��K�_���<�P�����E�r�`���
nT�(La`�bg������oH�;w��υ�G�{\���[��d���3��4	j�l0.pĿG����Z�"�n�{Ƕ�yXR�&�:sۇb��0"��J;��a���)��pQy�Gb�]�����R�H#|��|��_*񛭗wa��q)y��X�.��q�'�M~�.��V'�Qi��X=�
���!�5��T��8�[V��#�/4�A"d,�8���_���.��.�(Z�L@���P/�:���%�ǭ��c����;�c�"�g^��,G���bU�tT�$���1�������
����+Z@ �>IC�o<�n���1�k[�W��=h3��Z ¶�
n>���x���o��I��2Z�� �P5v=�ޏ�"�ŭ���)�?h�&Ԋ�D��-�G��7>e��8����ѹB�����'�jy/m�F�r���oS�^�F/T>��r��N��~O�ꕄX7�;��ْ���b�3��X���(��,#�Y�.�:��(B��E*r�l�I�ćl�W&��t���m[��V��s�|Db�K�T3�P8�՟a��d��\ܹ��
�#0�t`ރ�ƹ�e���|ܥ�b��M������0�"�m�2��,=0.�����:-�*m�Ξ�T��Vϖ�0vU�	��QT��-�9äD����|�[����њ,m���������U�]8
\J�]�ϐh�>�m8^\:��*�ub@���Rm���"�%��|'�U
Y�N,`lL��7y���8�ś�iQ[Y�'F6���j������Ȣ�[D�(\(�,b���OM?�� �f.l��]�2_R�o����O�X5~y�㹭Н�5B.m�d����ٽ��XEX��+J&	�-Ҷ�8W�g����� 9��Å����V�GW���Gt�I����	ۦ��;߆��$�.�{�-̈�$��O%�g�����y;7P���nnn,*�f��Ĺh:om�\ۏp[��n� �ϓ��m���M�-�3^��4���#8��C��G
-�t�辛o0	s_,���l���&(	=v�`*�gL#*R������+��F�ܥd���-��V��Z��5�L?9-ɰ�Ld��8��%�d����&7q�,|���\̍+����/��Ņ#X�M'���eE$�S����P��C՚4��֏Sq1W�泛���f/?�p�_�*��<�$��)P_�z4_��؅k��ge�3\���ղ{��-����
H��qī&�Ɍ�>�eVd���z�y�܁/nؖ�dk�"����+UA(�櫲>��l1�s�+�82�	k�R�5SC��E�Յy �dp����o����&�j5��a�"d��RJ�Ô�Y8��h�]��j�6 �~VN�R�㝗\�	�܂)�6Ѩe�[;E߄��r��EXZ�q�����O*3�y���B������.�V���i+U`����
~[M��D�����+V
��݈�d��z�?_OG�).�ӟ0f*�#���(�2}�z> �{�!p��s�#�	Ӂ˰�Y��T�<ɬ��CS;G��2��Tg)<B�2��p�L��n��$��	5��y`R��j*9a�bL
7!�C�q�o����A�_��g��2o#�j�T���~2sX�l�?%v��uǈGiRÌPNz�[Kug�b�ɬ�bl�)���a����+�fN�W>�,�\T�&�[�Oƀ�Bo]0�Iu�ħ:$i:!�>K<��Ԋ�u�`�ʴ�v�j��v2���B���k�+�@,��A���jj�.dc�P���i��L���l�V����E��ks���*
K��S�f�-Ԫ��y?�b,�M��������h`�$,����Wb�	L�lj�C���2ks���07|���O�I�잰��\� +�V��>�7�vV��S"Ĭg >e���/(<~V�����7�'�� )���`��_V�v��;������	vBoZ��& �[�����"�������h��)�A��@�)��m�"�@:A���M���t���?���@����b�Wc�Eb1���ǽ5Z�&��yo���#��<ʃ��#!�P��;q]��h��ng�Ud#ΟRR����>���2J�rz[ �#Q ���%���� Bgp�X �s����o��HB��vk�h%��
��H�-~�aɹ�n)`D���֤�2��\�)�<�3o���-���C��_C떛�rE�=Gx��l	��Ӗm��� <M��O�N��s�����=��#��ƨ+�m��{�����#�/d��a��� ��%��~�Va�'X� u8��6� ZQi���X���V����L=�ҹG��h�X��Ö�,���O�^�">�O�y%��A�Sf��Y����܃�Wh/�h�_�o(���P�9�F���X�P]��3Q�ٌ�{�JP���:i�tqk�|)I��3���}�� o��= r�	�CCnT- �0�(�)8Su�x9��-��@�<�Q
VVq��UE-��"�c;�mEu�Tn��h����L����~��>� J�܈�V�8#Nl��^Ȅ�����]6ZH�.q.��V�u����!^1����o���Ry���Л#dU����7c��30It���2J�±�F�+���R�qNn��|@I�WyH���G3�S��>������l�7Еp�-6�<��_�GV�hmw�?�.M�(�	�Vԕ Wj�lZ�;ß�hԘ5Hqw������/�|:U��=�^�^��}��>�OD�'��)�|��xr�u�Y��I]����5u/*��3ky�X>)�"�0�ҋA")��2V�&�����
ܟ+8�B~�3�u���""R�Pg��9����7���,�)�W�>�k���3���M��L�r��>iY��l���Ӄ�V��8O�'C�2)V����/��N��g�R7ܪ��VgL}Ut!�t�P&�,����涶���c��ȟT�Z�cAA�k���L���	�����d�u�Cu�Q`��#i8&u��`�M�r�o���<��k	�c�g��d���s�&��0V��1:h��q�)���yc�����ۇ�e¤�~��͡j�O+�m b�3��WM�Å�Dm5����N@��s,[&,p"�VZA��d�������Z΢����{ɖHO�ː�~kql�|��Z�S�UЧ��S�z��n�@��_�ʃ2u{ֻC�u�9��\���U�gE1+w�d�����ج��K�FR�"7���h͐,��خ���~���z���9��g؟���)e�*{���QR_�?@I���R4��~E�깛�ۋ�u�V�+���M^����U�'-o��>D�]��S3���d.{��ĥ���4��?p]��?b�e����1����G��[�{c�Lۘ�&�Yg�B�Es8��!�5�g��c��|8����=���;�&�K̨��b�ySX �l��?syC��ֆ˫cӮ��0L[�卮�w���='���n^-���ۡ���y{�ѱw�}Z�J�b~� żV^�ޤy>���uKb���zƩ�N7;7:,���V��ΏU"��,L�7������:+��_	RÈbG�V��l���)�>��� ���[��퍠HR��\8��&�d+�.9�ܯˮ�0�������k�k��8�.�H�z6�������*s�q��1��1$�3�i�e�{����	-!zT8�`~�=��Xj���Ȃ�ݝ��=�����Je�t���f�;ӤU��K�v�K�4;mM�.9�R���S�!�I�*%r a�]��Zqƫ�� i£�:+�MlK�}%L�^MJ����=�/���!LE��(�����8�
����'�ʑ4�U�@���Mh�=���ʬ��rg��~=:��.�I�ض��y������=˽�%��n�4��qcY�����4�~�(�<�bFN������W4�]]e=�a�ԏUт�:�G,ūx�o�<SpP�Ti�q�md9�Pmd�H�����7�шЃ@���CVՀY����K���a�>����a�~Q)!���Ņ����O����btUC	/Dp����Op� ��Jɀ�[�Y�CN�zjG���]g՟���q���������+[w�)� �s�	͓�{@NQ
�;*�M"JO�k�vm����Q�v�x /�8����_
Uq�d���\�.p�ʛֳ��_uj�1ג��1�ȳ,a��wԯAMC
7���mV�m̪B34�8���hJi�ш��W�}�|Ϩ�>ߖn�"j���Q�%��v�&��_��^7�tѧ�.���f����+��7��YV��� Oy`6��O���B�-���˟�K�	��kPT�i�Y�J���J��� �z���A��Kv�Lߟ�R�0���G��'h� (�pt+�����b|�
	�]�镜���LGB-Ȥàw�N��W�Tc�����=f���s��W�F⭎��������9��Y�D��������na��N��HϮ�K��8k�-W�RM�3�p�R���a[���XZۢH�*6R�Rk�"�U�����d?�}�Q�aב�$�Ol&�~i��|�r��ϝ�i�4�����(�Z�cV�r������R��Dٹ�c����U�߹�Yi�Ġ������)b޾�X����d��}�6�C����iŷ}�/,u�)U�ʻ��V���]ךz��7v��)����/l��0�A�ϯ�MN�V�TٱW�V:�����G�����ka��mDB�[q�{/Y�n�����iM	�^NԓY�1�Xc'�FS*H��tm��x�/x��4��%�F�rJ��q��3]����{�h��P�|�K;i�\�W�@�.ԣH��@s�+�Q�;��Cc��̯*���&w$Q�C��	t�K����'��_�r`k����q~YifT�,l��Lc�T�n}�Ռ$�YJQV��|��e���E�v��$sr�W0O��N�L���!�x6S���� <W�x��[���Y��+� �TR�7�V��&����_K���KL�������"��_���}��2Lv��F!�&�O�r�ȫ�t��Z\9
	[Zj�{S�`.w��b�M����HmZ���n��bo����L
0S���zR(_7X�0;�%�ֿ��ڥ��MY.��pڊ�ˑj�$���8-��ӝ�k�{٫ڑ�ђ��[֢(?��@�>�mpB�υ]x���Ǎy�;2n�<d�=ϋ���YǴ��f����a��7�E⨇��#je��zV��S)�O� �A*�Z�����b����a��n^��d��$�K��;\fb���z�g��l8
��丏�yM8���6����H��hO
��l��B�MI��T�_PU���ş�*�Kr�d[ڶQ�y�O�`k;�~���h�}���r -jX��ٶl5f+e�g�\�����ǂf���<�[N} �%��C�8\Ȝ�Zp��u�=�c �B�Oq���Ϊ���a��{�|�P�s�\��ڵǿ��(��b��2��z�%(Z������ǟˉ#��.�/��>����?����a�ii�q䊤V���<A��u�>�c��Eq�܌"��*UT���,@���(( ��2�昔���q�u��Ƃ�R��i�!4�XK_z��{w 6�Ԝ���`�@e�3�xo�U�FMV�;Nc���N`p��N�� ����#̯���ώ��)�����dtz����':	+R�ې�8"?x�8Ky��1;ޔY�1�V@1���)ʂn�(���KCG�sAa*wN�}�܎�㔗]�4ҽ\R$J�4y�����Cl�a�|�^}1��6ɱ��1C�.�rD�U�m��}=���D����\0�-w>x��}�3��D��)�,���q�4�h���[�s���74b�h�D��g\e�
�I�v;&�";U�H�5��a��)VZ�
��/ȁ+P��O�S��C[K�w��#����MU��cg����ػ�j�Oi㴹_�ʚ��4|����_zvp�����ʷ�U�M��}�QvW�Gum�OV�w��j��U�T{	��wB�6f�ԖR�'j�蔗j��[-&�j'���cU�I��O�z���*���C�Da8Z�������FaoeJA���>����-�P�$B��	��M�f_�!���c��zU�`�3t\�W߶}z�
XP�}W���L�>X'�&�L
��x�&��
�}����U����v�/G�"��� ���9��P��{�Ew$���T�ϭ��im�.u<��c�?ų4V�L�*%��%��,�-kS�����T@Gw�B���)YŔ�	�.j�a89�WZt�W�7<��҉^���|��z?v�zO��gF6U�Ͽ1S��H� ��\z`��<�;����	����(��fnmU�(�ʮ��z��kJ��a�SW�;\���˫ݐ
7N�ы��T|����)���\�+E[0jM�\�\?�	&@��Ճ�{�ɪ����	*wo�xr��}虘��@��T3�+1 ����op�56>����K�I��3�S��*{]��	�vsɤ�%���:G<-���x户W8��n]e
&���d�$�w��M����RPl�O����L3�Ugo����]z5b����Ώ���Ƽ�Z��:`�N�ÿ�u�LP��A�`-v#����l��c�Ni��rc� �Ѳd�����B�x����Z=���Z���:�DϚ�a�r@0��{`o�O\A��®������p�������){E$7�x�����'>��v����,��\��AH����W,K����#�Av�=s�F�Ȁ��L���O`�&A#��}�U� }�X���E=C%�Z�� <0�C�&ZB~rl~�+z	��|�T
w��q�:��7�e0�a���E��a���T��C�Z�idR�[3�hV�O�}�u�!mZ>�Ho"}�Wk�mI�����#]v�����������|"ӟ�G������IfD5�1��+X�"�&7�qP��4�rlK��#
���>�k2l�y�In����7�8z����Dp
��\i�a��i�d�8������q�c�p�PT�_ <}N�����M\�%h��l��8d]j�j���R\Š�T&�L1��j�䤲�(��G��\�q¹���T�,�)ـ��{�'#�j������}^R��}֬��Ulc�
����``��f.�q�Kex������D[���2ݤ&w�6��T�D����|��@�Ï��F`׏0��y�z)Op�aGa,Q"�������(���x�4��QfM���"ِql=�iI#v��5���4s�V�����ox�#�NRwbL��Jg+�t9*�����kj<��4�4HU|�xv:i��jrR�Po�AD��?{+@��yY�S*(��S3p@��7d9w���^�qd��E�m׷He���i8������NG�/����ǖ�B��#�>����O�=M����jz�~߀B�Kcs׍TU��i5��֮_�W��g����� �-\b��4����	������Gs�J��{@�<K�W�.�*�/UH3��Y��b>��pa�o��5�f��
�e�r#b|o���O���������R��p��z�~Ө��8��r�*�,B�3�����c����j_�ԉ{-����\�Zj͸d9)��%Sc{�}K���:N���(u���������+,`z=�	�}���S��:b"��1bo�/
���-X�=�92�RhZ�VlW���3f}s���w��΀]CP�.�r0%J���T��4a��Ĺ�:��?���$�T�{�J�r����-ഹDɭ��
P�E>K�5#!pp}CD�xɲ%\�*^(��ު(���ƛr*ْ��S"h,����#w�Q���6x0>����h�q�ro����$�%,@zN��J*����
U4Dr	ӝ��č�fF�EdoңA|��gO�P쎛��*��ag+:k_Z�<����Sމ/��õ�A,�1M�XH�7D�1��w����Ae{r�U��J�/�A��Z~�R��Pݯ��+O�/���7��|L�����`vxW�dU�PJ&o���yz��kL����V�V�@�0�ͦh���%Z<ퟧ�����Z��}">�	���v��J[5.X6�!Fӝ7��<�ee�1`�@~-��Y�aןX���Az(��C��Jk���5��B#7H��Ҭ�e���R�I�H�6�I����Ki6x�MfA=��[����l��aW�pn6m�6�%�6B��)��_��1�0��Ļ�{Ō�O�_�}�~�u�t#��lj;���2�����
`er�o\��MLw����x<�4-��Ï�4<�=r|>؄�����<!�谮j�?����nT}(�����Wqi�,O	s�����4M��kkz����X�m�P�x�O-�vp��˦f�+-r2y���q�0�>g��swo0+�}��%����=y�l��t��+�f
_����X-[�^q^��|�&���E8+bf�#e���{kk�6�	����oǨ�4���6�',Sb�ht�!�R��`���A��q�;
����7�f�sN%�:w{�&�2���VWw�o	�&��v���2�wl��B��T�gM���z���n���ˊW�������W��)�`�@9����迄K�j�O�3,)ް��o��b\��	~9�1�#�	U�'x�!����V����������_
ޮ�V���Ӳԡʷ�{��T!�8�{����R�A٢��\�r����w\m��
<R�18�D~��:��4y�I����B�6��`}	G�@�-[x@��z4c�>)8��RI�6Y��ϟ�,��T2��������-�9���8���T�6bӵ*=�J�U�>�:�oEĘ��:��,�����������̊��˓�����Pd�6�&���nۘw;R�Zm���rN�r�=-������<e�>ft�Y�ܠ�`�=��U��c޲��v�q��}7u	S�5CK�]k��p�s��uJl�`!��&M��Ȑ ��d)��˷�������FN�J�����L5�b�����tʒӝ}�����f�&cs�����;�~j]�8�iI�t�����4��*^E	 ���<%�}c�,�P-�rtr]��-[�=��������VЖ𝖩���UO�ٕ����H%hs�Eh��g�FSɠ�x�V3���S� $&<��"!���
���h嶣d��3EH0K�7���U�q)(����r��z@H<E�3'Mg�����b�_��5/������Q#��Cȥ�~�pםmg٩Yp�?�C6��֎3�/m��y� ;��x�\s���!���Gbn����(q�C>���zS��.2Q�c�ͯ�-�>��m�rIȴY
�ߊ�O_	��o0=�ؑ����z/ߔc��X��7G�jh D����-���Z�����e�}�e��/2R;y$���1Ё�r�VoX�g����L\�g��M��o�ńJ���1�!���V�
��f�Ȩ�ʹ1��`F�&�%Ź��RT��~�]�5Ht/�q��]"&r�B5��Y��:#�{{�Mab{T0��P<�+Y��v�$�{���� .i;��z��qB6�sL��P<B|����61�u��t��B��T�EU�� z*dQ2\4\������@�U�U��#�l��=1�jb�wA^7*D��%�)��ďf#��YA�qa����}P*}C�]:���'���j>{m�����M2�KvFF�<��O�8���JZ�׏�Wo����|,�'b*B�	�j���<K��0M���+#��B;���rV�H�d:]�O�M�����9R���x�vB
S�ѱ���DZ_�p��)E�>{I��.I���S�ќ�����f�9�y�B}i=2��dt�V��\(h���������5�=*x2�X������[�|"(|�{�0١�[\� X�u���DD�]hk��s��Z����`��]<VZ��(o�O�j��y8y�Sb �A��φC�hF��KA��J�爤-� ��Z�;��������S遅A��5�N�i�)@���Oh(��H�j�턀�yUBߨ@��=�7�}D3�|`~��by�θ��|�z6�<)yS�β�|zC�2	"��x��X&��\9q"�w��@��� }W��a�� A�S��,aEh�J�����`R�=Af�N�1T�-q`٨�r��ލA���w�x��X��Q���`��~bL|܍�4UN�]��3�3�	�hp݋�[�q�_�	{xNE�
]V�)��
��z�z>..���V�_��K9�1�gG����Q�����>��!�=��*�- 2s��>l��ZB>s-���#�l���qt��oÌ�q!ox`�Q6��:23���й=uŒɅS==�6��l�/+6����Eۃ"�md�Ns�~�k`z@�9UБ����w���e�_<>B���N�l3L�������odG�9 �=r"�N�uI\ia.��^H�X
��}��CȘIS�`��}�儺 :��&xK ��Z�yq<�a9� � 5�ɺ$~��E��	�b5��I�E.��#,�O�>~�!��_H��۱b��ǁc��E*���Õ��ñ���=:Π�|&����pyʙ���䦵�@mnkrV��lGA���V�tS1�O`&k����1�ل����#�٫M6ٕ3���K�78�B	�8o�NIT�鈢R��}��m���8��H�+��	��fA]r�w��1"ˑN��Ҡ�M�����]��������Wo�y p�N؛d�9�x"۠�OĽ���g��)�ȅ��	c����ag��Zm�ʚ�	�J6�]T��S�\�����c�<�i��D� �b"��ET��r�$��2���	Z���f�1��Z6�|��]N.���l������J,��z�y1[�������)�Y��,s�oU�n���?�T
=����z$�pP�W�ݺ>P��&�P˥13�&�TdyQ�Ʃ�.]�,���R��t�W�\v ��n��+����O7a�P�����s�i�����H/ ��g���f�9,~=pϜ�:����f�髿2���1N�_�c����y4)g@�7�f2p��U������6,_��*e?F�y��$�-EH�W�k���<Ϡ�Mf@��|v��=�������%�)ɛ��Z�
8v%F��h�CX��D(�;H�(�#�r��J��t���$��߹%ٳ"ΨM��w�O+{��?5	�n�|6�+�2�Q�d!�	�yC�Ԗ�_G�ʯ-I�i�{�!�zՅ�\�֜���:��b�|]G�N����Q�b�*��b�|U�r�2a�E\J� �@���ѐ\R�ĺ����T�u}ȓ�0%��&�x�d���|�[S�:�VǉyW�h3�F�ՠ6�������N�w?�o�����aj�C!�2T+Z:|A�G�:��&�V�ÛYZ����Ɛ���eju<)"�C^�� l�u\0�_��l�r,<1�5>I�]�t�5"���w�^X �����ɢ��x�1!�/]�-�Be���ԅ��{�y6��@���`��O�k#ŊT���`�p�[gp`�O�^4�B-��g���6B��*]��]l,N�#�Mt!G���-�"�`>ҼL<���;�"�q�F���'p�S%Pѻ���4�ƪ��H��5|O��+��1K�9����JR��j�����>X�1��_�F��s��o:�2��L�9�Bϧ�,]�e����wG����{K�Y��Y����ϸ��<��uA��Ϋ�/�{Z˯k�&���_B�g��L*�Ⱥ<�_ �,����#�X�1�n��;v�J���F��啟�3���%튜�?����r%�{�fv騙��à�L�4J!3�#��fE1� �D�A�����H�4�g�F��X���l�T�I�&���x�ϛ�mb1(?����SViy�!b`��UNR�>�����൶FQ�o%�܊����8{axB{F��C8L�����{D���F��G�Է�,M��6
�f v�X��H�Ӥ N��Ⱦ$_i`�����G�-�}/m��e�٠��^�>��"��4��:����f֓	�C����lU>�ro��H��SC�����Y&n���H56�Z �«`jy�'��9���/��R����0-U[��X)BЩeo�L���Y���&�_�����T����ҙ��s�^��HV��>�g�n��k���l!NW���nO�����1�O˻M��BĊ��vjT�O<_��i����G��y��?1�~�����+�����ܧ"�G#��hS�0����!S���M�#-�
p�[pg{�fj�����(�S��YI �6�Qd1���r(�\啐@kA�v��9w�9Ĵ�o����u��7C��~7���y[�^66L�$��%��5�o��J��l!�Xg�ᨂ�� �=nf'��+���ۡC4*l��ٓ�g ��I�+^Řj̱#�1`���O�F̾9x���=��fY���<tp����h����%o�"�G�_�HR�ed����#:�m��f6?�7W��qʪH�� ���q�2z�͌�I�w��v�Ia�"�ԩ2'?٤<��Z��C��.�"����0!����b��dUP3�D�u������1�{�U|��r"/���v<�|yZI�Ff6 ��o�ދ�_ubN��s
2L{y�m\B�����H�ۡ>'�л�ME/�۾�܃oD�0�-��{�����P�U�:�\�5�S��s?am0�fk�c�\�X�Fe:����X��,�X�����?�*˔��t���}�έ��}�80g�I��p�ć��ɄW>$��Hd���k5���l�°�:=���SW�0�}���Q?;ɚ�k[4
.R�1�%�('0r�M̎t���&��L�s�H��l��b�4(��M��Sg������'eG��T�Ʉ����j?��G����&f�X��+�^q\�}r�Yҹ�u�����A��}Maw1$�74\�3B׸N�O�[@0��tj�p��&�s��[�U����L����牤06�Ј�G��;�X����B�n���zj�k�0�ʚu2�gM�'r�!�}���);���u{όM[��?�#�V%LNrK����Z������M�|��GB�jڄ����7�F81#���D5t��	���l�z���"�6�t�۾@bg�'�߄�����έR�k�yW}����j�V���T����6Cg�XI�M�i����d8M
US⠾�������/c��XiCv����&lx4�P��*"EE�
����8�T�R���[5I��M�%
CYҞ-,���nx�����3�.>T���ڱB;��=����;>M`J��[mC��[E�vD�239��|�-T�BCVͥX�ߞ���ɦÏ(Ì��N)ݩ�8[�BT�7G�]D>��]�9�MGM�Uf�FK?1���C'���叧�g�Rwj�J� ,�3C a*6Td��2��w7�u\��l�9DT��##��X���9P��RQ���am��S"ʩ�T�q^��������@��z3P���Q|�x�5�钡�-d^n�fRQ���4bT�U�y�Q�������{`
���<�̑Z�
�A5I�Yʺ��:N�+KY衤lØ�|s�3z}�gR`�}�-Ô�c�a0��ށ�y�q�]�f�;j����se��$�r�>��`����ʨ�/;'��4Z���o0�����J�cD��y�����q�r��Z��J�E?Q������>��D��l!l�v՚��˓.�$.�P��Պ߱��q4�h�8���a��Hpd����`$�<[B ��j��EbS�F�o;��e,�`��f�vT�q@�$��N�Hf��������1���2�g=�`>�n��q},6G�q�Ph�Ad�mC����	� w7���76��1��ݟ]����,�e�jѪH�95|���wy8�`�[X}
n���~d[KɄ�Pd�s���-�n3&�1*sN$��ᎣC����{C�
��5�H�*�]Ձ��6[��Pq?/�`�`-&_\mrhn�DG��%��e;�ĝ�ib��z��JiK:�E�n����F�Y�k�7ʅ�[����M�Lq��㲉):�TV�ܨ��aU��*Uc׋�Dz�p����Ϋv�ӄ����Wt��q�0y�o%-��;��3G�v���G�h�+�2�����s�w�O�Qb(�|��?��Ag�N*�s�tͥU+��m���Kh�L���.���|��nZ_�6]���`	�gK[�o�,�H��X��ݝLX�E*NP�y�������+*�v�17{��o�m�����sC	�Ecn�������>3Ն�~穡L,�����6nɥ���(�_�^S�ݷ"������[U���WJ��mi��'�Ӿc�l����t�ؚ<�zN$<�Y�Pf"3���0���S)�~���vN(}�%�x��z�R���P���V��#�J����7�;��'lx?qP��zn��(!�h¦s�5{%m+H��4�F�� {�n��@~p�`si�{Ƴ��[�#v祻����̯�#���D���3��a��{�(��qN�yf��;ʐȐ��K���T�4&O¿K�@W`jFP�	x�Ep$������8���m��JE&冸H�q���+���+����C�E����(��5�e%��N�M�"���|���'q�!(�$�|�V�/���v��>�83c�`b��o%@PKz� )��I�����Ip�C^�Tc&��X��H�(��eV��[X�4b5mr6���n�)>���V���$P�3�I*�*9��LX
�s*x����,Y���7�4�66_f�G(�����R��)8�FV��d�����M	=�Fx`WS�|�K+5�ȼ��ߎ2��fX��D�ɟ5��V���'��	�8�a�M�UAΡv�%�_{	��Mv���Y�'(���v�4I�*��Oy0�*�>l"Vc��\�3܃G�4��H�� Q���d�`�t,R�������f�j�\��V�$������ߓ}u��ñO�G��k�'�x]%}"�Dg�y:��h�H�Y֍��mX*��6ϏRO�;ׇ�����?LC^� �S�G�
v4�� ���#���AFd�	��8*-2��� aeo�y@$ջ��门~�l��z�bǺ:�I���x���{�&��59P�A�Ɉ6G$#v�fю���(��|O�0�4A�
��=���ۉ8?�z�%Y皺������[ƾ��(�6��� 2G�+���t���F�O��h	T�L���E?���O�P�%���e�>u�ٻ)Lफ़=�S��w��ͻ��բ����� ����a���W��f�,�Λ��$>�lҲ��td�o��K��sC�Y8V�g�;�(�2C�������;��1��2��Wh$����ӫ��@Z-�L�4�
��8k'zyO�@��٫�܅��+��|l^;��s��l�8��;��E�l(�o���V�gL'��|�Qt1�+{�Ϸu��ߓ%��f���sQ�<�+~!��	EY��V�:ԏLR�w�Bu�rp2�H�����^&ne4�3�Y�Os_/Dg5R��z !Ø���v�!�j��K��^$O�um�[|�8��H�2[K����6p�ʨj�>nE����~f' ^X6PY��㟰nM\�u�����������ӛ���0P�tc�嬗����0�Z������#���reI�}ɈnDp>{�N"+��WP!��ܭ�\�5�%(��s��o������ ��l�W��wA��7��İ��=�^b���w�&	�N-;{̺{p���LFv?5g�p���$g�_�&8@ ��u�Y��V;�ݵ
�Z�����SK���:�R�n��ޝ�������L'�tQ� ŵG�H��iȡa�d�&�9kl�G�����g��I�>S�T)�'>���z��rO�@6o��"�)2�Q����9/vL��L,o��+���� MN�h������,�z
kӣҶg-o��z��%��/D��v-V�Κ�CA*8�J��l�%�h>��z��7�F�O��W`�c��q{h���Ti �
H�<|ICu0��
_�z��8#�~wn��<:�-R�ļ稣��z�e�"�{�u.;���!w-�/�I������������~]j��T¼vc���3��ؑ4�]K��~�MD̔�_u+��k��ܘwt���B��am����h����aO�%G}���4�k{9�S*8�ٸ�Kc�N�(ޗ]�C���>�5��$��Gc5Zf K�>f�%�qؽ-cȅ%��!T����LkZCk@��c��G����~d�۩9b��6�H'�籦�6 �cU�r��ʯ#����9�̴��[�$����²I���UX�>��D�ݹ�5|�}W,�PZ��5�4���S���o+��yE��?ٷ���sB��_�?�r�b�y=IK�7&�����s!�|&��9���W6b���E�gȮE��������iN�#�'/�4ܑ��9\�;V��Ju J�r]ݞ`��eX��%pv�5:����b^�Y�ML#P���J6�n���!�	�&�E�71��+�ԃ��%�Y���@͘����	%�����΂���G�i��*{�^�����!�&�Dd����|��ю���ށ�ֱ�6`�������3�`r4U�0�L(�l�xʪ[�;���1U��9B�9mS���U���(Z�~�Hָ�<����%zњ�A����&��ƌ�g��k�L�e�����<-��#ts��+yVPx%�0+�?0)�	���3n�?h	,)IKn��!��4��i&������A����4d���ه���ژ�j1SSM�����dA���X��u�I�F�)�t����V�:Ӟ9M,����L a��$�}:����nހ�b��'�㞥[$��	�!^t�O8}k	)%#��m>c3!g���'2����o�v�����$�V������ [.d��Y��n�UAn���V`Eބ2����|	o��D�3�w�sz�-0����WϨ���ӱj�k�{���
��uDXf=2���P\��6�f��N69��ޏwv���`h��k� �Ơ4]qi�����e�먑�i�
OU������a���{���V�Ҏ�S�c=�ѝ���D�{���)��3�W��<��C�~<�n�c+��ȯy��gu컨�P��F���Y�[V�F�%�K�
Q�,��i��B���@e�y'1�\$�Fǥ�­�_�{ `ju��ʙ@�������u�R�K�>Gn|�x�y�T
uX]7N���e���9	pw.�rҔDC�����7%��,�5} �������8�,��bmD��K�� ��z�v�� 1�"��?/㜕�J�D�;]����.^&��Ҕja9�IAұ��^Oc�8�gL?�z+?I�#�r����B�k�L��d�[)!�ڟ�)�)�����YIddIB{�}��0q�e��*��"�谲:� ������<:!n��;֛Tl�LA�k�Y�ӥ�����̞K�	\K��� �bM��Q��!,��P�PО�4-xZ�\��9)ؗ��8��D�׈�E�����PkS�pcփ��y��#I0�wQ3���5/vF��8��Y�TR`����?O�ժW#=�~q�s�U^�Sx�9x���~�`J�%�^���dL��q�h+�ȪW��B�'xir,��\�DI!��s&��0��VV���W���*�Bk������5��bꌝ�%(l�� ������{yטp�ր�dj�';2ba�3Us��`�#JgK���KC]�O4�����V:�o)��^������.��0���KE�W���9����ʳQ�ylވ����0������hF��m�8��j���͐`R��x��Pl23�D��g�pg��[ܡ��C�(ay�c����"��;�@���$b`�ſJ��3�귛ܨ`^������#�0�E*Zw/�U�����Yb�a��	q�IB�|չ�j#e�p(�Tx�����섊�*�پq/z�.�d}7��@&e��:�н	uXU�L�(d( ��U�{{20�[(ԣo-����mT�k6�A	1	a�=�
�����$-&�B����5a �����X��K�X
D����t�̏�5ғ:xB��Dq�i�B1��iق'ln3�����3�8�$��Q)����Ѕ��y1F#tM��X����p��C��@��;�	R�{1�� �j��kc�6�Y�,�G"X!����ޔn@�ZZ�	ҨƄ~B�{�&��:"7���!�M��*2�;��*i0S+�dٗ���I�%����^����	���ąV|���;/�q���s6_Uj�A�U�1;����mYY�c�����j��A�����N��!#����;Z(4����TӁ[� ��!p֢W����o�ҽ��5|�@B�\�g���y��P+�q�Z�4e���֯��4��x-3!�_�:-�.x����<+�K��������"c|<@sڒ7f~u��N�ֱ_H��o�;���_�E�]�T4Ϻ�s����υ�Q�2�t�o������a5��gV�	Q;����T*�h.f���r�y4D�衴��I|Iяxc:Ag�%?B�|r��)��� ���6�$����`+؏`���
.�>}�D[z�ـ&=m����C��R��wd�>�ӓ?zvõ6�+:�gf�t?s]�a/��|d�dK-��a4c~�ǳ^ѱ��x�<*�_������Ε�.I���a���D�YFn�=u���C�9�����@�_��۶���g��U��:5wDTă�t?�wJw���*->˜�"����a=!�ɃOQ�Sy`e��oY�oX���Q��W2��K�����r&������;�`�')�~�6=<#e����O���Ġב��}�M���9_<�i/u!�Y�����K&���<?Ic�͔�
��E�X���?��*�S���$�_}���tb�yD��Ǝ����q�W�NX�Qտ	��QZ��7�LVCm¡�;�%S]��ԧ�\��#G$�ɿ�Z��K!�\�9���#��3�0�����ѻ���)1{N�q\�t�ϯy�$��}蕬G�O*�.T�ְU�]3� J�s�27z��-����W(��SL��N)��ԑg�&� ��i���nr\�E�6noș��7
��6l���'�)nbY���y77����ًiK�82	m��:��j�$�F���@��ZF��NY�,�ޢt�4��r�u�wڝ0�$xZ�JG�ch{vBv�Ȣ�/���e�A!�)
b�Úws3h�*r�v�p�?x��!/���s8Aw-�Ǡ5G���}������\�*B�[�����w�FT�6,*���a��Ej�����w4�H�E4`�L�h���=,���Ʉ���΂+"b�ط�����R$`�Ѯ9cOY`��^���4MZ6����$In9�􄊤��� ���ȶ�A�x�rc���3r1�3Ǝ)x)��d-fv��$� �9;�3�&n��lק�՜��Bl��LT����%x�A�e,0H���2LK���Ot>��q��MK��h�{b�:x>���3��&����箧�&&~�B+YzPT��T!&Mc"F?=@/^ꖫ�ޭG�=�O�LPߙ��q
e�yO���8�c�ź���qd1fE�y�����5i��L�5%,�4^�ʶ�`Қ���3F���1�O��a�P�_sQ���0�_��\{��0o$O��Q�$N�T1}D��%����P��K䳊��N�>h<1]ak�a�(&z���y�XR��r!�j><�늛>,��<�p��kIQ<���P�����je���4�!�EX�����W�4g6 2!%�D��l�,^�:jOuhg�3� �U/�:N'�	���К�'����ձ�����c�I�V���������%Ҷ�+����3�v*z��iÐ	m�1��HSo�@���"�i�MPu�	\'����YZ�T�4�YW�rN�Ew�<"�r�^�]4�2�I'�ȉ��9)V�ΨM�4<q�˒�m�{�w2iVi�ľxw�r������0D�e{M7��b�Y2e���ۀi�#�Ka��Ù\�w?�I�'��N��/|)0� F����x���u�tYY���~3"z�&YC�+6t��Y:��|���5D,�'Ѣ�c��
���#�$������ʪ8\gu��G|~�"FxΤ�_~�v(x�WӴ�H	���u�Y<�.��_m��ϑ�]��沏8{?�	�,��6Aɺ����Sm�b��(C��٨��n^��_�9�SبZA=�}�߾�����6�z���߰����7lZ
aX%��4o�B�y(�� ��]	9�E���&��W��&�ۚ@w����4�Ƥ�"���}�@v$�#� ���{�P�	ơy����19}�B,���W��yhF���0�r$�{�AcH��u��4m{���� [;�z�}��a�����J�%�����9�X�`�w9�j-��˴�]��R2����$��*���?�)B5�un��2.�n�g��P���E�Fp�JA\�X�)�����vy��&u��B /g�Ȉ)���l!��BQ +v|r��v��9� -+�-��[�� �M����5r"Z�cҍ�j�j�Z[�in
�A�l���7C'GYk��(�,���̒�Oh�`���$OMH�0jLjzX;e��٬����פ"��d+֋>�z���o��κk�������K�Թ�c=*˥f/<.���1����'C����	��V��(��-1��d�(��|m��w�����#�h(A��^7��ټ�~!B���O��0ѹ+�	$�˃�78�}�;�n������s��P�~<�>cK
�����&`�#ѕ�`7�r�~A]v U:��Sĵ�5�
d~Q����u)�3�j
O�0�v��8���"l���)�@9�g�'BҪ��aGm�8�qR$[��@� 6iJ��UӐ��e����L޿?�]��t۟qO�G)�u��v���+i�R�x�h��2�^�@�n����h8f��-�-�T]glF@j����W3+9�J�����)D����̶ڣ��Du��NA\���s���8�>��7?ܜ�/�hYC��Ml��6�F��ރ����y�V�������؇<�S��QRo����q�a*0�+��&�=(:�Ok�Z��q-�6�]3����0o�v���..��I뉚�۶�G�H����$�츨��2��g���!0n^��J��I�`'�����P��nO�N��V$:.�!������5�Fx�F�w��#�,�װ>�+C��|d�h�-��Sn��N��>�1��+���.���#�$x��>og� ~� �+�2�ג	��-��WtK��R}������9Fr��J�I���� �i)��j[�C)�E#�2E|�[jҲ ���j!.y����}ex��ak.!�k�!�z
TJj�֭߱6�b��(Vt��\�:��$q
,w`9��z�;=�\e1��!q߂���U�6��0���G�~wZ�!q�eW�b'zzl(�	b�e�̟r��v��nі�X�N(��<�h�܁&���!�%Z���	�N��J#�85��˪�>����a�ɗ��Nk1��q�n�^�/����	��%��Un�Fo�NYo��e��J�ivF����8����Hf�X�'J���'�3i�>�@�bf�	�o�}�pCi���C&Z���Wq��������3���)R��:�1��_=\o4���C��e�'�}�C���g�������_��J�b�m�����_�,�W1�>-W��2�J��k�v��[��2^,�=X���Lx��ym�	)�`Qk��sH�15'i��^�"� <�%Wj��a #9Ӗ#QF9����p���?G_(�L�ΐv�`vB3��6�f1�t��Q�h�w.zf	;H�~�ζ�*b�4��l��K2�N��lw�Ř�e��1�@f�c��:�\��@�T^��4V;O�̟,i##,��ˊ��A�*,�K���ݣ�L����r�&/� ʁ%j�˪{^Ax��U�nب͙�\c22���az��(�z��W�r�A^�}�i�:�����t�_���$%Ux$�����㢔�|6��jY+�;��X�T�=�ƼhXCTN��o$ѹ�n������T�
.�YHt����
�JA>'��N�&�l�%�0q�ɠr�r'���eo�m��f���<����!��~�s�o���Ek����g������!����c�T�Şz_,�l�h�0lq��d�\Z��r*ǆ�Ѥ����q��3q��;���"�oh�YI��4���/r���V��E��\&����d�`��}�a���z�MWT@�p��%l��Ҋ��x���[�E�멳��[�#P7�k��G�.8���r�0b|��8�ް���u�$�~���æ�u�"��v]��?�yd�Ka��g��ʇL����=�P���U����J_s-W0.�8��p'�a�,����;$����J�_���॔�W[}�����1H<�Ǵz�:vu�vO�naA0�vv*0�8����Y�-d���-AJ�cy� �4�@�.�{:R�tvTg������\����w��jm"p���d�4He�\Yv�z81-�[��J%z"5S��\�	��&=�sVre���:U.'m��yi�|�f&�4.I$/�"��£HZN����2�q8�j�	"�?��K���z��i�����b��A���|dNi,2��u�lq!�0�׫WU~�xeR*��#T�6!�N�~/ǹRO�W�V�L��1�@��Y���Z�����
 �a��"��L��T�8Mp6�����4�d�:��P۝5�<�`�'\�����Q��Y4���]�O�')�J�X�C߁��pb���:��tV�ʺL�ۭ�La
�� �+���/�l��1l��a����͖-�:�˃/��d����| 0QǛ�
�v ȍ+�{�.�N�fT�����GbVNW0�v|�X�ќ����t3��al��"�{������f��
�?�
��������I�pp�^��A�h϶Zw�1�|��+.��jSb~���!ݼz���O)r:��Z!�u����8�[-3�0&��C�����D:@��M	�MeEAn�B��4���ZQ�ï0�T(�F�����Rݿl���H�Nl �g��Ӳ��e� xHIFɃc)�^Y���f�;!b#'N�ܕ�<:W^�����( �*4�(&b�⿼P��� Ψ���?�QoG�}m ��b�l��o6�[/]\v�b�}TY/�Fs��xW�m�m�l �D�h�=�Q�!�ԕ����7�"8Z�h���mn��G<�wiz jB�,�;.t��	M��bۥ'OY�5�,Ԋ�g�d���d�l�{�e�m~I�U����A��6b�Ē��1Ib�����AFb@(���~����Z��MH�0��pr����q>�m23�l"l;�����iwP�N!*M��m�?G1r���5ާ��N\C"\�y6rʼo������s-�j�MO�[9�e	>$���'���7m���^d����Kf�A�a��է��:�\���%�}�fI��V�Nn�˶�R|?C�L&]3\�.�'H��R����-��p����Ł޿�y��Ѵ�����'�(}�ml��;~ݲ�f�]=�7�@	ۣ�+_�-�/����&��&�}�Y
�1jD2�!ڽ3RM~�.�~����B����6�1�"��+�9G�X��>(�W�T��rkf�4��#e��F���{�sZ�-��� 6*ܛ�4p����~�U�dχ��=� #d���:�$������R�v9��h��g�֌������YA��4�¿�Zش�w��#��ѹ ��%��x�Fj��U���E2�u��|�O��<��K���w0��6>ٿ����d�^��E_ �n0K�k���V���ŧ�6�ƻ	�#��\5�K���e�b����pw-�{����M���k�"ٲK����c�u$C�v�S�T��3����]|�ܫ�z܀�i�$=݊}Q��K�	��nƍ�4'\Q������@��^���Q:�,����jvQy�%τb��v�����j����0�l�k�c�6�����]�����2OH�������+{��`ܣ5���f'#����՚�QyتS#�!
����LM�ڤ�ͯ+�f�f�E�#�y��ES���U�[Om��pL%�]�\5��5S^�p�o��2L��>����j�{�@;_��B^rx����Y$�n�xױ&��$b��ㅱ����}������!T�o�ѓƵn^N@��$=P팦R~��O#�L����ↅ����2�:��� !/<����6�bdl?�b��W�]�wvU�K;%������y��ތ_��8��~��F{�<��iPŠ/{��O��-톻���b�el�½C��@̑뢏Bv�G����	���I%#��N&M�1e�Q��D�ya��@�jR/�&�ō&�����y���1R-E��a�4�p���kR���q�N�4��'sP��u(k��@��p Z����C`/N1F����z��V�~�L>�}��[�J ���x���c�dw{���l�����GjK�^r��:(J�7p�b]1�����@�+6�m�����Pߢt�SU7\=#A���(U�%��6�z��h��N]q��_�!�����3���]d�Dr��G��n�ԭ��t��7H�����AN�ڲXX>?a�뗫���ʖ;�7���_����=l�m��!������[�>��{�!$'|���C�^`�# 2�#�c����ʓ=���ؐ����ң��yo��B�d���К�(м�U
�gB']�ls9�c�ɥ��fǜ��깥��NP��v�'Th��:Io��9������1��(z(�0�C2eFKS�z6�Ɲ�(&�����6�����LZ���?�t�L�[���k�F���%���B��g��nc��!?��V���atK|s��y�����pY�3G0_��r���t�����r68�����Nr�w,R�#*4�2��-���y.Kf���!z<��NQ&ޔ�߯E�م��1�pz��Tm����]ź3a�QM\�k祽��)a�k\_z�v�rM�f�>kWIuE7@u�s]gs��	���lk2�]O�*0f��0��!m{�s9���%��7��g
�U���+�w��#�y`�L���L����֣���:Pe�c){�<�$;8S�Fr~���-�en�v��zo2dqLN�չ�	
XGk<�8�ۦ۷563C�ng�Gs�Z>OB�U})�(���N����Z�Z���1f�\8X�䕏#�Q캷�E��b�lE��(�.q �[E��R�4Pc�b���Abj٢n�#:�$��3j��Ǿ�i��Ҙ�B��=tL�� ���g��	m�6TD��&w�ξdF(�� �?�U���Q኶^�P�sD�AS:��ɧ
�!�	���Fh>�[�9�����!�Q=��oMZZ<П�9�Y����{�n���O��$��ై����#�2C���j���[��TH�����.ڋ�Yxĭ���e�^�j�#s��������x{��:�k�)D)�׸� ��C����iT�0���o%�0�(8[�*���l�yR�m�[̯�F�f������$�g(%�$=U��M
��]�ug�b	+�=�UV�%x�ܜt��}��#�gm�+�8	����!�so���N����3�'��f2*��")B����'L�7�mJ.}�X��X3�UG~��P���
ml�r���xk�dҩ�\b�E�YS�o��1���uŝq����	�^�����{'G�{�lmRFI����~Y7�f?t��>�H��xC�g7�g�AX�6����G^�B������_��?Q�\������]-D�{؃m˫�~��;Q��
!Vy�:�V��/&J��
��+�'��d��&���C�X�kdx��i��|��zf/cb���ʑM��^2��&=���"אy���LL���p���7���H���p�r��I���H��!��u&�Y��XSd���RA.�G��mg��,��
d(
N��:?�1�wb�=����}����#<�����>�9k�b��VI��	$#Z��1ew,f��!�Q]sQh�DA4nE��s�屣$�Cz홊���d���m�0��r�0D��oc�����7��}��9Í��:�Qo�1�دh7���^�|��Y w�:C?@�X�"�����V����6p��*�I�Dc�x.s?�"�l��gA9DF�\)�P��>(́D�4��៖������0z�P��]�Z��ͅ���S��N5����\i(=z���5z壹0JH����P�,<)
�'���7/	�xP5��*-� ������N� �����rE\�}�bрo��sY�Io-֯���P(�yP2�Z�W��MB��_H.ٵ��Ҥ�GqgB>�!�(	�[�Vo��U|_�i��i<k�qX�ʘ�? �"�(i݌��N��3>�2��R#�^���b��	Dr�s�?٧͔�22.熞>xJ�\߁>���R
�>�c<���(O;#)�)aX#��K�%R��ߍE��}���N	�?��#��?�=K1p Vk3')�*>2j�4�U���6%��Ү$V�V��Q*��g�:&5Rx��!DAx�C;!�n82��������FN����j���O��\�AI�k�C��6%<��N���L�H�|�41�����^���X�vb�d��CU��(|7��_�@�]�4Iۡ]���O -�9$3�c��Dٺ���50��%�=�P<N����ǫg��P��ٚ��%�8�3[�}�,�<ehx�8�uvl�)��A7jK���*N͇4�)"ˤ���C��Gk!6�[�h��W�����t�'<-�+�B�p)Hsa������ܑ@U�3� �J`��Io�)�M�X�/#��$���D�?s��	yx�'5������8�
��C̋�VLX�#z%F��P���r�So%�����˨ɿ���&���2Bm���
>���ury3j� ��Űr�K?��g�6��K}j�̳��n���/÷e.�_�-�J؄?T��H�ˬ밴�a���Q��n��*O���w*��OXE�R��,��kb ����7���[��}��/���_�S!?WU�^+ �.�c4�Qの���5rgbg��@(q!�Ժ�Be~ն䵚#+aJ����9�H�B�)='�L���H$f�0�جx7ǜ�4"Q�w�(gĹ�V�o�b�M� �~�����W���T��2"�]��;�kO�H�GK��6J�������D �U+[������D�Q��/�f)HT�����n����jc��t�
��l�}0�"��Y����.��Qjz��[:�jͷm;��ȩ��bd@��&��X��ۭ�Ia�)��)�&n��X�6�2J�t[���F�H�G�g��l`+l'�Y�FyW��#)m� �sڲa՝��j�#舲��� �b�~��ϩi�9ր��{r��נ��8})F��FTM4�T:��:.���j�5oi��X{<���Uo@��|�n��-m^E���l����5d��݅�{W!��N�)XF��\�=1�&(��V"f���I7�p�<��u7�)մ:=�ac�/]��-���a+����C���yi�6�r��SG$Q�r6�����Nk��>(-nb��Ƽ�C�XgH0���ק�<;����!|�aR� E4<�k��02^���W��m��y�5L�q���(N�`j^�g�W�2c��o��Α�������r�18�W/�yk�� ���qh�2ǣ(�_#Y��7l�=H�	$wp�G��Ӳ8��u�#j�ڛ�1ʛ�(���p�.EwSB�nr��ju(�M0O�y�K��71�`���؊��Y�E�W�;��k�L}������+L$��)�t�HkLm�7��T�pp�ٮf���s����ޕ����=5XBmn�Y�4���C���nZ�S�z���?��>}	�&��W	�W���|,`S&*�9&qz��Fy~m�0o`g��h4����p�jF�=DΪ�1cɣ=�I	N�_V��П�i25)g��C�頻H�)�;C�y`l�����[Ȳ���;r���S����Un3�x���I����n:�Q�>֬#%�%z̵w��b|o>�N0/�1�6$��=,E�+FӪ�� ]yA^mM)mmJ�z�W���K��!���ϵ0@j�Ua����BXT3�U�j���L�SJ��*�F�nVkt8�N_8wj�.�n���i��5<�刂�v�\���JJ�B- �F�כ �x�r��v���V:s^s�ý��pf�@uiK�Vg �Z��Hk�2�@v�	vS�L����;�����䅶��"y��$�h4�H����.@.m���/�C��uϔV���r���]([�Bm.9���55��s�L1G���i�^'�n$4�_dY����x�qL� "����t�Cbb�|���߉�8{'Pll{C�TgpDȈ8�
i��Z�
N��s���n��7�Z���^{٤�������s�@Z��_�R{�.�5���>z�2� c-��F:sQ�{]�� t��u����eG)�?:adڳ�:��4^���N�ah�b�&���IV"|ʧ��mO ,Y�]�3��,�{�,���s��$\@YH�C����z�&�1�!@m�)��z�&T�$k����~�� ��T�����:��C,^�4 �C#Wa[��Ng��w���e�D�y;�w�|)_7�k�ɧ�.�Gyo�<��$�J�H��w�e�Y�eGt,A�ϳ5KY4�����HO)Bhw��tQ�x:���1�H���Ǔ�RJ�����컾��<H��?%����`�Q���h)�˲ǵ�sQ��
��)��j�fe�m˽�c�\�AݓZ[�Q5�P�"��I�*N��&�q*�<�P%�_�Bh����tP?�
�,?y筵FjW����@�,8;�2�u1mPhۭ&�	���ws�*��?��Ђ󚈰R��f �0&_�~@�4���
�PoU�Qg���� ��m���iG���ں-4.�㧊�GUD+�Y��v � �:�W�]�q��y6���*�2P����,D+Y���N�r4�&0���=-ĥ@���[���g,�=I�Ď����˩��	f\�[��D��*����r�+�@�.�8$����ۭ�&Iy�`ʨ)����b��0QȆ��b��Y�����)J�R���І:����o=�����M��#�8�Z���*.��%h�f���,��9�GVQW�U?�e�lǐd�����y���|�{E��dـ���<U*�\�g���i���"��w�~K��᳊�7}TV2�<�2�"�LIv���%���gfi��T\�T߃��`�?���̭2�j�
�����U�+�|�4=Jβ.�1�.oL,�"&��$����:�:���m�˞�5�󆔪9M�S�Rz�C�����H;a�G,�������/��g�'�/[U�Q�(B�E���:����E.�|�O�J\�͂��+��k�o�������E#]{v
#��Trfr�7�i��jwr��Yg�͟�(�a�����F�r�p�p_�i�h���z��23�B	���0�$��T/BX�I�
u��|ا9_;L+/�2�=���S|��z,-��/.e8�T�@�ط�l������I�9w�c86H�p�n:���^��BWĳ5v��p��G?IY��ϴ\��J�j�ȳ+J�� M�e�5k��rr��&]L�M`��m�2����
X��1����H�3�~9ld; ��h�--����7F\H�X����Z?KY,ȕ�$!6���͔'�d4Tf�Q�JS�)��I���+��������� ��(o��S�������2*3"��r(bv8ja������J3�hHXs��"����g褟;`��/ҩԕ�XI�N�c@&��w.d��0KJ*�7����ȝ������6����p��Y׫���I�k%]B�p�Z�.}j�2\���S��Bw/!��j��̰k�����᷶ʔ�I|��^6$�Y�����6g勬1"ܩY%���U{��<���ꓵo�	�(��t ��f��s�[���0N{?Z8Q5��s1=�
�bo	�z��L��C��D��F.FW�u���^:>O���l���~Բ��Ze��p	^�8D����<vć>3,T�\ X�;�ۿ��a���q�����C/�� �"��(��d���p�3���-���ƀI#�_![�]B��*2��=�z'M�Ϟ���Ҥ�^�'(F8x��q �V��!���v���v�3(��ǉx��୏�z��6F�w�	*r;7�B�uZBO̶t�ŷl ��V�(�_P�,=~Dv9h�דy��g!��(|�z���9�w�G@j���U��F6�vhJ'bŖ��-�%�,M����l!��|����[�Sg�ѻ�J.w�X�|Pnn�Jam.Y�pkk�j���ں$[�!1,8k������b�i8U�T�I��=c륈&�2�a�oʩK,o�7�����Y b��z`��baB���7�0�&��l�
/:K���p�
r�M��Fp���%[o�i;��텛�~&l�ժ�>`vv��Nj��fHJGF�����|U9�@�%�jS�7s3LjHj���eJ�]����,zE�M�/?M,���������{N*���a�\}y�,A"������y���,B\�ԟ�3|n|�ː�8�d��#����W�4�@�V�Q鵛��)`��@`�Q{��)Sx���?����TNJu�G�-s�:�}*����׆�r��F�qR�u� �xM�bT :��W.���>-��H� ̎��5�> <L}�
�!�p�H^��'Sj
�����S������XŨ3�8L�s��sʚ�����'{��rJ��:{+Q�
��.�b��T ࿪��N|�`�2o��r%��4X���r��֤f����GZ]�a��Ofq��=�)�RJ.Ci[������5]h xۅ��;z��u�m@|��e˚��])1m�:.Q;%}��� �M�,yxWI3�촖���Q�� �B����.�F��E�%�1��c���*艄�`a���4r���_���˴pm�KZ�� K2�J7%YV!�Ĕl���
�����0�^��v�/��_�pz=ȵB�Wv������D��1��&D�i�%�
��o�*x�Ս�{#�H��ߺW�Ī�xv�v���֐i��7qu�K���Z�`���y�d?(<�1}f@��Ni�%)�#	���  �mb�J�ʩ$���Y�	�^1����y���l����·[Y�������h�γ��:�M���z&_ ������^��Ρ��{�srL�R�������3Ε�g�FL}+4jm�7	�QlgW���-+��O��	���cC�v�{�gU�v�ѓo3���	cM��"��՛��3�>:��e�~
u��7�&�����H���<�y��>NC�?�#A?��L��G�P�.��@X���So@\���}��t�!Uwڼ��{��i,�Z��R�k�$7]֌��%�V�JE��q�I���Vǎ��q��?�� ن!'pO���	�E�+h�`�U�8�67�nM���U����'����e�̪s�u��Sh<��m��ޟv�G�C�G�;�����F?����FeKQ�l,�yl�N(�'x�6�2Ԟ�����b�����^s+�̾^�_�{�E��r���Sa[�Ȫ���Ņ9�FQ ��|�v��!j�\���(�Y�s�,���s���2�ZC�(T��·�����zS�y����#1��(�c�b��aV����
�
�j<3���;���A�a=@�\����$EϤ���o�R��4M���n��va�������fVd������eJAдB���R�� �62�o�HK�g?��r�}�z�|a�wY#2��5�_
kln{�'��#v�N�`��-�����-{���Ysi�M�?�EmGx$�۪�Of�L]g�e�-��XC)=�Z7������)����d��n�3����m���k2|�F�/������ǹ�m��2<���6�� rP�닗�����qgq�]�S��S��s�����$ت��o�u��<� �[Q7��T. �_Kt�*�U�i��������d�ٷwy{�*��Vp5M�Gq�m�'�
ٌ�	����~cS��_�őY�D��j�&��T�s��!Fx� y��F!�.��I�~k���o���w2�q�Y&��2�B�>��Q��,u�z|��zgUQ R}���k������XGf�9B�?ƕOD�M&��QA�dL�8}9��o��\ a�~��+��Ha��&5�(MD�M5!����'km�?: 1�[Eqa9�!Ξ%���=����"lWp �D��9I��k������� oh�(#�%٬bMV�8�&��Du7�V�ڇÆ��ව֭�3&9��]l�2	�4�?���,u���B�t�.�/�bDØv���"�Z,\=R6qF��0�H��&p�|Ii��ցQ�t��62D�ZJQK$ْ��v����vf8�͝Z���j��A���=��p
���r�(�F� �Q�	���8K�����2��*M�o|D���_������:�О� Ff��4QB_�c�X삙7
o�+��7�A^m�[�C]�_�Ʃjƶ�$Ο�̆)�(ܯU?Q����u�!S��D?��G�*������wJx��<����B��KS��d4~�R?��i��k����f�.�]�3�������N � �В�_G�wu�5$�~���	^�w���nW��N��T�\���u0��9>�����u�q�/��5��xh-�n��XE��<�I�V�i�k�'U����Q T ������YU}$ac���9ߔ6=Up�:f�t������������ƭ:ds	�t��Sv�E�%	��dQ��J�������N��|TO���F�F�]:��9
�����f� qBG���8��om�q��ĢNV��Mr�9��M�b����}i4?f�i���q%�S}|��$��q*I��Z�o�Nc���-��<S`P5�##��J�l:]	+z�wr:�rԡ쐄'��^^�R�jY�90q� D7�ٶ�RB/z��{N�s+>���
��zgB�u�l�@��� 0G��!
U������NK�!Y>el�������{8�� /R�H���ME�_�2g�$� 88��*0�W6�F̵}'�;�<�Q��mdq����.m����R���,����Nڥ�M8��"!Kػ�⼸w��)�#���Htј4�.7o׫�k+�l�%�l�#�d� ��dl��!�I�K��$�$�����[	���xt��V

��I����o��/����0t<�f�A���H@�[&^��9m;(��iE���)��](5��֨�����+��A��^��-�>��T6�|���o�ʬ;���Zn�����X[v�%BBP2k �t�]<�"jRq3�c~�8��iXԌH�.3��~$�^�����	}lU��3Z�Q5��;[�ul��-��-�5���g��r8�wY%�6w��ꏐ�����Ȏ��'����~lި�44b)��%ٙ=���>9�Kٽr��a�H|Ab
J��C�oWd�2RK;+hO�N��t�I�|g3�=U׶>��q��}�?d�[��L���k�9�VCAn�N��?��f[�9�A�K�7��L�r�~f��<��N`Rɗ��7U>�V %j��#�˳U�6�Ÿ��#`����c3���T!�#�}�-����\	��Vo�U+Š���{WA�XFoy%��l5����VA,qm^�!ԉaG�pN�n3 �[�ۇo����𹠹�ｌ��L?V���5�/H|W�˷��q57_�oߦ�˨-�:?��6^�AhM�?>W��/\�!*�`_����G�����+�;2�w���{�v�	,�b��j�5�GZX�V� �6�p/���	��5c���wt�F�}G��-��ON@���k8d�7��}�kB�����(��Q�]���"�2B`:��1=)�Uv�Q������s,��*X���2z�tL�
� �'�A�i«ȅ�����t��H�˱|�o%
l�3��3>��������=F5�4�Wl��ǵ�S_	�z����#˝�Z�՟��W��Q@0�D��� � G�b�&3k�U�=�]�t0����rO.�?��5��#����0E*�J����Q����(좔{�{�-��V������hf�ˆx�U��Hr[�
P��벧qj�{��(Ʃ���M��*2:�3yp���hʖ5-+g8ե�s;�B�!�������[�)W�lm �^7G���ٞzn�@�+6���U���dP���K�Y�A��SG[��o����Ƣ),��z�,6�Ω�Vt�뚡
Ъ�j|�E�z��2W�.���A�)�D�ݰ��F1�_����.�~xtgW�r'C�,�]�<��Ģ�ݝ'���O]�z!�ާ�o�@Ūu�VEl���֖g�U1�~W��3��"�~���#T�T�D�^��P�e��f y1n��Uɟ��M��F}7l�#A��Yu�� ��m��M�&���`G���1Лشn�w?���
Q����yY�U�~�q3��u-M��fL��ߒ_H��r��XE(<���)1E�;ά~&nK�c|#s\�c��Y�̕ܒЩ�E9q���	ѐ��6Êˤ6�tuH#���cKw�#4uG�4�I�4�fd��G5[S�+)ϩɇDe�p�
s3��ui�q��s��ڡ���7�J�~�b-��l{�>��E̪������ V��?�0���WI�q�#��\)�>��l�Rٲ#ٹ����z�l�u�޵b%��	�%�/�o$*�:G�����TW0Y`7�F�Y�����.�~a$�e*�/���,��|�9��>�wR��?[l�1��a�pf$9H3p8~�.���^�Xn�u~z�w<��FZ�>�����P7Tu�5;>�z �>d��&8�dr�>D���[$�O<B��ܪ���nI�VL!ݙ
�Ub	X�����!�,����佼̈́jk�
�\Tѕ�R�=�.�ö*�4���#�r�|�̠�պMz�~ssz�<d$8��`'�m$3����w��q�w�I��y�p]��uv�1�����K!�G�Ȩ0�����ZH�S�b��|�a�f��͒� 6F<Ϥ�Z��H3���������X�r+:�Dԣ)�����[Ө������苁��0�D��'6�N:��-?��R��Z
�' I�ΠN�n������1��4_�R�0$=�a�w��!:I��A�󁰆6�P�2#���~S��H�p�X������K���O�k�6&�TJ8��Ne��PҶ�m�J���O��jm����f�pR��2
����}R���*����T�W����H����4��&q���.H8�2��G�a<Y��xމ��.
4L�9d�(\���	л~ �wA��ř�,�1�"�-����%i����~	|���-1Â�mhc��3��H���(6l�o��=y~�B4T6+zx�0��I W �D����W�:��]L���K��w��A6�����wN�9K/K��5��"��:p$
\v8C�3 �b+�[�Km����k~yK��PrwV�(����M�ʚ�����'�O�ѵ��z����6��+�^~�+Eok�>@�0�#�Ad��J���Ǩ]F�uo����lmu��aW�I��.�T�A��s@	��J|��FOa�޽��M��R��m�q8y�+ƨK�Z��x;�E6��ٹ!���:���5�c�Y�7p�*"���%gvƀ0�	�B�̡^9�p��Е��ƪoe�?=j)嫷|�2�}g�`�ΙU���F���c�׊֊"�rͮ�`$���� �s���ķ��tN�+p_�oD|�(6���ee�(��@{�P���9�����`�j��)�WK�'7��>��`��'��l����<.M�p����5�yC~3M`�6Q^B]`~$�&3��i%����c�%��{y��l�r�4U��<�w�o9֦��$�*��&~:�?MA[Eh_��=�gll��Y���.:9����cd����F���܄&v�v��)76��*Q��I[���&e��ߤ�m�U-�m4=Ћ*B[>˖�'.���!E�\#��Z���a��7�W��p\ɵ/����M�R�BN�j�C��t;�G�Zi�?�ۻ>�K���S��H���?�K��"ѧ�HBu�?cS�m6d�y��ץ`^���s��ʘ�k��Ct���%��\,-�<���9fb)fsx�1.��g�ѷ9�Jf(��\������6� w�s���v`B`�L�~�z�6�8�F&S�aط@|I������D�!K���R7F��+ߥ��ey�ɷ��-����>�~���4_:���6'��wi��jN���ȶ�},(L���,@1~3h'p�3#	��̝�2^�H�>�6��0s��&���m3����󥀼�j�"����@i��b�j���]vޣ�F�Z��
�z�������N6S�DxOp8Tb�G4㫀��pF@e�G�*�^��X����U����;
����5Q!���ζt"�1�U��4aIT %4��l+�̸��`�ЁY�$����;�[ SJ"�`B#��!5Ա9�{�vO��uI�o������#N#��]hF�d�� < �v���!}[*�
c��y�p}c�Q���6��\����5���D>-�8l�pV��s+��Jm#���e�ANm�{L�G�c�lO9�����V�)�t���$�A�.��z$���P��<���zt�.#�4ۯ���>��]M	Q3��̌y�s�A�Q���B�ӟ*�=Kh Z��lv�w�A1`��bJm}$`�xC�� ����Yr_2���#B�8� &{�ʞ���2�>�?s�;�V� F`uZ�N1�
�`��²�ЇX�*��2w�*X�8P̴����;��̘��d��.�&��&a;VN@��8
�u���a?���Vw;�7t!� ����P����t���`��T]\Ǚ�C	�E�W~�g& �φ]���
���q�w}��Ɉ�������3����K��p{$=zֆ��7e�~�l�$Z��~گ4����|
��tė9	�?�W�@?`r�t�3�D/����d�h��#��������4�(/'�XƟ:�{�F����2��]�:iB�Ae5�s�\=1@'�=o���������\j�;ኵC�؎1�-b��
�拯����*��n�#�I������"�$l�e�voP��:o��w�P�I��"�f8.����5���S>0ek�����Ĝ���� �����l��MC�~ �o�ٙ@=�"��#����L��h�f���=��&���~Q1����@F��q�p��-�%��-�?H����=W��U�L�zۊ�}�p�N���	�[��2����apqc���scVtM��a�6|��P�:� ��4b%���-�نy�w�)w(�#�k� �-E:5Ko��ŗޅ-�ԩ�iH�ȯ����h���r����oԃ�f[�~rYs�WOCƟp럵U=�VGSyǮHMGW���>ֽ�����a���b�#W����vM�;^s�4��4���C|��>���V*�����y�eD���1�+���S�r���B�T�Z�ʣ?�Y� ��4�P�&�:�XA�,�y8Y`��7$��%d�f����N-�2����N3Rt�]�n5��a��/;Y7���SR�1��)�V7��Yqz���*���=t$�(=���=`aY5����S�]m����-���fp������4sn���l����Vl�GwpciY��ETFI��3����X�R������q#�#!�⥶������O�{=�nj�b"$�1J��o�_�Q\�*�P ��x�Y�V�ܹƷ�Wڙ�v
U@���6K�No[��$�{<{Ɋ�Q���ǆW6���)3��0�i}��ct�U���y�]��,o����~O�'�ʐ�~�Z�{�]UCIr�~+e�Lߨ+�$�;�VK|�bc%�c��H����%W�QMz�cBK��vw|ˤ�#�-�^�u/1V�u�R���к�m<%ė+.�4U%�,13���R���V��G�7��I�J#]���Og�����r��bޘ�|�E�t�ņ��_gci7ʌ�.D�pR��+S����e�O�'@-�4}�S�L��F�f#�y��;~��>)j�n>z�AS��39�0�|aUX*�����bf�x��X�1�2r�BK��;N(*P�#�T�]zl�N�lݴ�7�/�(o�����"� l�SK�^">���~�,�]����2ZJ�Hݏ�\��Y\T��T��O�e���jZ�8#ַ,%){a9h�cU�1��Ccc�F�%ݏϓ�o}�1�z�W��z���4�[��h\�	��9n����N~/�'��P�)��{�D��K���A��ff��c�-��5�	���\��W�9�G��RgL�˜9�ϭ��19�4x�`��O��h����g��avC�i���,���j��C?͚lH�i��iP��鏄�L^dC�
{�����H�SnF4�7�ģ�y.��q�UM��*
<|<��X!�b��>��q�q��S�n\���ų3|�:Rx���m���|EN®� �{�,�Jh�eq�� >+�	����L8����<���v&��5��\�c���	���d��i��,�e����7�t�%O��~T���[��T�4�qM�"����� ��f���J�iO��N��&#1 *��^:���3��U���W�b��&u2��L�� Ꝼ=y�FJ�a�֡�yPS|������'�4c��S�������#�	���D����Y��������Tp9w�I�E4�a���������˒6<+��Rk֘���!���m;@����{R�/#U I�4@�{f�2�{�TG�E����%�F�ˠ_��~D�ʟŖpB�p̐*��w9b&������7 ���|5�:j�8Ʃ뽻�\a)�ړ�g2B�=>�N>�x}�iD&·�|g*+�M�O�d�D��%*�p!�QZ�䔔�Zy��@*��K��ͫ7៓��7��_Y�lyi>ԣ@H�m��{��A$���nwo('�M�#1vy�v�vΈl��̗U�1����>? /��@8`��w����78�����ipH�����}kSuE�go/���*�E��B���B�\y�k-�Ab"� ���^���صD��'���RmDG k}�y��%���/Y����+��5�F�Jj��N�;��h]Ų9�̾�����禁��\p��οBDB����*�Q��ؽ9��G71cCЃ/Y�M�W"f$�n�x��F����'��UH�T/�f8�8ˬ���A'yC�p���`�s��<v��rW%R�t�&=���s74U����ԙ����i]}＇�χ����J���vcY�W���Aݾ����Ԁ��hVI��tU����@�2�U��:8��� ?�v��+uq���6E6'�}�)�-Q�N?)q L�s�UBPe�KK���d&���N�N2zL/��cJR�T���º�}�?�
?J����<]!a4LG���AH�}�?r~�5���C��RA�h���9�BAOp�A����R 	S�=c��h~�z��(U
��|}�5P�	����]����,4�>$�����%y&e!�yt ��.5��9�5!L���l-Fc���.)HF�(x���J{OSx�����E!e-N��<A��H8���0�k�{�b ��S��Egx.6m_{�G^]/���)���֒`*Mte�k���m�>Oj���)`I�� U��!ڂ��I�3�֜�j�������XI�&���/�yV-9�����LulU&�}��[bP��"^�ȳ[�/I�0��l��O�� �|�]Ҙ#��j�4��Jf�~�}�v�*؁d4(c�������LS�Nn���=$&t,��`}��6�-�Bk ��a���C�\�Zl�;�]<��P 	���w5��p(Zɼ�u���_���aM�X���`qz�o���lN����,P+�cS9�T6t0}��{���zgt'6[���/��1�:�X��6�I�F�z�F���2��%�j���B#J��p/yx,-��X�Nê�mV��?���f�1A]����˳�;K��fɠ��utZ�����)@��O��_�c��OF���,�M:=#�2fg�!�A	3��m�!�c�P��y����LL&�4��X$�[�N���v}�?����wr��1�>�U���u5��*���ؾh��iaχo� B]�b,k�'�Fo�4D����
^���@0����]w}���)P��a#Hv�h��X/�[+E#��ei�P�R���d9��Rp&+W�Q8�i���A:�5�hbz
T�y�B�(D��Fqa��CÒwۧ�ɽ	`ʒ[c���@���J�9�=>�mO�Y�ye�9vkp,y��J�k� �����QԳ4���iJ�W8��%7V�7���Pq4�*=�2��t�
�[kr��л�{[��Yߚ����7��
x� �pG9���G՟x�����}�M��D�%���F�e��v�Q>ó���%�3*��ޙҽ=X+B���xeF:kv�u�~��W��U��l���֛C��=C�L��+�����aZ���� ,Q��x��VE���r�]P}�K�����,b0cf�Tz�Y������o?t_͗�Q�AD`��KZ>B7e+�P�]1�ZNW١���B�Z�� 6=n6!��P�Q����/c=���6'���g�2c^o�[p�ΑW��*֠��ga�	���� �{_ZvnL����&�E䐪婬;,�;@dG�>���)�d�����r)��U/��c�����|�#���RA�3/�鹡���εN �C�$���QA\DW�{��]�''�f�y�r���*�/�l��W�b��N1�:�� A*�끼��3���y�ē�V��'�_&*�
^u�� �y�[m�@�i3U�녨Lڌ��	�2
=����l�D��)g`A�Hj�<�
�XZZ�W!��H�]��	O.?e��F7��V�w����?������AY�-����ic�C�]�gΦP~���;������f"�l�AD��^ �R׊Z8	��H�^��!JZ%���T�ő�Hq�C�d��������1��9��L?#�R��I��e���Ȟ��׃aFw���*-���(�I';e@�}
�s�3#1���J���M��=���rðX��p�#EZ������1�U��Ϳ�9��������H?��ϱ��
C� ��Ɩq�wWF��#r!o��u����'�g�� 0G�:8����)��>:-}&�o��W��#GVW�n^�_.�sKtX�7�Q�����S����;AF����~�J������a�6��[� lo3��j}b��$uc��	/�ym�:-|����C�uwA%ߔR���=�)�K62c��mv͸���㶵<�j0�^�)5s\����UϽ��:v�,���=�����\�(&&yj~������NFʚ�m(N����;���QI�	B���]_ӠA�:t{��zM-|�:��팸��0))�[fV�c�h��e���=�OF�w�t6j�=�>N櫱M�`+��x Nۤ��򓡬�G�1f
�)8��l�G���U�8$L��0��G����o8�%���k���S�,Y޵�7}����<�,���q�>�S��-�Uj����G��%�Wq�����~�w����efg��q~����^u��`�	1�5j��rE��Y-K)2
R���;�l}y���xX�tM�-2y�{]�g_~�i �f_Hp�����A��(N΄*�T��n*)�7d/
">/�ځ�����1]�f�#������aU�����6�ܞ������M{3�ȞQ���5������ßK��Th���<|̈́|�����o�%���W���%��~n7K\�S�k$��W�yd���3���:�!y`�ΰ��/��)H��f��x.�+ʐ6��F�_����w�h��}��q-R�ߡ+{?I��0�$�n�K\����eh�T�1�H���ޯDDv����\0r��̨8�A�{w��!��>h6�;ϥ� ��0�����Ӡj��	��>��ʘj�(���(�[OD1���g[=�z�"G��g�T^B�nv���"݈(�����2���Po�qƆ�NǇ�;���T'�3vҐPD�!n�Ĝ'��,㩲��Fﲮ©~���/��]���6>���x:�d��8>�T���u37y�Vw��j����i�u �%.��WO��	���
Zn���-�߸�kt�y�C}D�еx���@qJ���VR�ԕ�`���(r�D~Km,�0R�I1Rqg�T1��6���j�r���(�ex�V���W�UIg>1y'�F~�mX}�(?/��� �����פ��V���y��f��/m+hOYfz>-�I�	F�`��Uβ���50�J��5<�ZH��ěׯq�#ɢ
b������A�e�sŁ>7] b��w�T�?����p-��>��Nǻ�����=T��X`��>�J|hM^\.l�&F�묖8km��RdѲ<:�u徣�w��!�҄�z�;�6��R�.J �X0��&W��s�/����䛖n�~XY�Q�d��[n�L�/Sy�D�Wz�;,�FX��}�����O@����B�'m�(L��ߧ�VCy;y�w�֑,�5�&}��6p����E�V���K1���%�����c�Ō]{n�����ة'zV��:�v���������cR����������?��]���C8E�:�`2��"
֞M�lIv�<��b`J��>37&qBP��g��*׭/�8KI��Z(3W��5ȶ��(���&\.�+�e?0{��rw3~�����ZR*I�/��x3wzz��QIQ�8K�"q��젖&+|d�PR6�	-��O����`:X��:���eۃ�j�OJ�SȐc�m�h5E��v��CpT^ܩo�^��K�ʻ�����s�˂J��Q���ijj�qcr��a�Ŵ���A�	�M2b��,�-��=�#���k�c�l�3��x_"S��K\���g�,��;K���������q����Ẏ�5�n�VzҀj[Rш.�ct�.,��Y맶��B(��1�n����0�f�2{��}�Ύ�UD�Q���YGRy�:i�����da�O�|���FWދ�9i �K�H���ɽ����4;݄qc�װǙ�tѺ9�������lh�.��3K@l�JᔣF�Ai�V�?o��]"-��0x()V���ų�2�©<���ŏn�F��G�8>���"���(S_�X��^m[��j)҅YD������}�N��@���o�1��>���!��M�*�B�0��4O׻�v���>T�vn���/(q������	���T��E��̞#bɁ���K���jL .�Ϭͨ$2R@kWkć�m�K�W��ֲU���k!l}��qʹ�׬Vj�i�����\4�Z ��x�y�@inx�d�Dxd�˽8M�U93� �&���k�*@�l5�����B�y�+6J�F�6�o�g���l�GV8���@�zhъ��p�\o�)�eԆA�������«.δ��f�t�㺋�b��ʈ
�z�f�ޒ��k��X_t�5��W霜�����*Qw.P���f�*���H~�ώċ�1��8�(����a$a��E��'y* �`��R��0F�6�Z�8��/Eh�Ō>W�����b �,vM��k��R׽� A[ʊYk3SNnC}�Pc�ݺ5xh�/c~9���"��@�_��]���4�D��`ѳ��R#*]������5J�l˘:K��H�`U"�\�ka��x]b�'n�K��bP�]�
�"��"-�h��	]��%U���ܯ�>���k����W�f\UN;_��v""5�vj+��|.I:��D����i�5>�a�p,����\�����Y�y&��v)�*���K�nJ��6A�Bf�4�ؓ~�-�JJ�T��[��jM�	����a̳b#��[ü~Zk���sb<L�����>+� ��[�ǅ��Ԟ�Lé@_���������BTz'ycݠ[�>clEV��w��n��v��y�.L�D ^�o[�J�]j{�X6��e/�@X��QUbq�i��y�L���"y�p��ī���檚�.U>�����{�1S����d�և������T=$�F}�� ��o0���]>o���T�+���Q�ω53K̚�_h`),��g}������u�')�Te�>����Y�d�����I��٢��f�6��L�x�o�o�K\.N[@�>���G'�IT�B M�����_NПO�gc}�Q>=O �����*�d�g`����(��#{�wM{�_:������o�f,q��_Ŕ�(A��	#��T��K�.�V��d�{�Ma��*�"�ޭ��Q���Lx��X������	�TD��6L��V�-���z� aY�]�2�.�Ϋ�4��3ݩP��Z(Qأ��Î���k��6�-�Mb��o�{hɝ��c�۲�{��1�u����)<��m���&�b,(��l?�B`�1$x&��w�$Up^/o�����3�^~�QVF
���i�5��>��ߗ����ci����y����ُop�A��>�>#�R��9��LT��ۻ�`r�������.=j��'a�5"��x6�Y6/W5Ll���P"Z��TG�!c���-���Y��(^%�Ԕ7�u��+��"!]QM�LH�9�i[9QZ^)���!��m�:>�	�x��d9�ب��2a�D�x��x�	4@���W?^G�-(���Ӷ���_(���1��_��Yg4����G�
���}���h>,-��Ю3���	���r�ʲ�����Scs~�>���tN���J��k�)���
�ӑLН5$:�yu�Q�����M��B�@�	$�؎��Uׅ���se\��a�&~���/ѷƇ�D5הQ�D[�|��[v �_=�|	S-�~3�8J��=�'/��-؜�>Fv ���h��1/�y��>Ģ�h�9�a!t���4=��{|�"<�]����t����v��4�	R�ʋ��l2�V�:0~8�cX\L7:�v`e�D��T�>�b�W���8>�x����1�W�M�3����JZ
{�vl �O>���*o������h�Y�|�2O+�5��ʭzd�K�hf*��q�|(^�K������+cJT�$x������w�\m��qB�I	���#�w���wҸ_a���6_�Weig���U���x�0���8����W������f3�E�I7�K(;�ݜ%>Z>�$�Y�0����Nw��-E@A+����<�2�O�u7�؅�^"/���~m�DZ��nL��9A)���A|.+~�8	L���?�E��S ?��!c����~�rڽ���ù�٭�L�erx�qﵤ�9t�f�����JG�ڇ&��F1�d偕�V	��Q���m�O����i�CL�ՏOއ���8�r�]� m�P�n��4���|=P���	:�������4�R1��#/�n�������p��j۔�c��#y�dE�$B9>yK\����g�C9�v�ѵ���T6�����9�&������+����G�nG+��i��Z�ؙ��K&"o����P��d���f9��n!8=7�u)��8iVğ\�Ue[�U�!JL��/u^�٧*|����($g
Z�#C��~$�a��܄�fMd��S�t�h)�8�5+pY8��SƬ�̱H�ݶC��P���0Z���~�1B�&ћ������̏��q`�2�N5Ѕw��0T�ׅr+tͮF"�<.7�	
O�]fwB1Qϭ q��[6�7��]�����{�'��D:SR�.t�o�_�EMSi�d(w
יS�����/�\���u�ì�sRd��R�|?ӟ����Ϙ,��0CI��/b��B��j�W'%���g6a����-�������)������ᒜ��ъ��t�%�����	J�)��~��v|�|G��� ���2��jI�:�p\�V:X�0&)>��Xy�(	���iN��m��X<E}ٱޅo������Y�F�^GI�D�u��`6��4]
�\�2K�R���V��Ȕ?�O�O����"���� �&��
-i|�+��_ ���cV����T�#� ��7��p�8��ȁ���_:�ً����ȁ��ǻ�k-B�WdH��2\�07ό�м ]��^߭��>"N,��/
���w*>��E�VԈ��� ������ai\
���Z���=P"�Ke*��&[c��cL�
:�u���°{�A��
���y߳,>��W��O����MN�.~ۓV���0�t.R;�"�\T��D�g�a��*��	8S�w\s�@�ND۵�?'�,�İ\q�6b��LBP�fq��~iT�)���ᒷ�)�5<����kvVvT�AdO��Y.oT�lSp�;�� ��r��˖ո{4�>��~n�y��f�G܏w��Sc ������l���oQ����z��8�^�-��'�@�jt�H��o��;;y��B���fEP��/uj:>�f�x�,:�8+���&k�Q�F�7���/���T��O=��V���q��;{./8;�����nN�2�$a�aȜn����pf�)͇�xF�qK��^��6��$X��'_ʄ.�B�U��Y�I��c���k�G�4��^�I��\>F��t����	Qp?��zq�*5��ФO�W�E]B�/�K��>��݃�sŧ��
w]�J#��f�k�/y PʋEZWb��A�X/I�m��&�[i���z�
O�����:D�`���H���Z����I��5�K�yn%Pv?�n�j�?H ���\���	]j� E� AW�wHZZ�����,b'�kB�m����D��: ���`�2qa{"v�APvoR�t�"B�R1�W���㣔[X�ӜK��"?�3�7��΄��P��'-�%�i�V3<��չ�>p��_�;�nq֒���uX����+}���9��;4(A�@M�g+	��5���S/5b4����e����e��"�3�X��>W��"�� �=�"]���p��4� ��_�`���9��9����:k�9^���[J�)���v����� �A@҃u���?�T�ylb��1��?�Q�\l^B��*g�r7���sʱ�y�͟zq�A���Բ�Y@�n����3�2�1c��^w(��z��"Z����H�'� ��{T�Br
�p\�JC�B1?e*�( ����-^�򭜥t��פB�b��)/;WQ��J�t���:��l�o ��ͻ�.͖��r�B������2�%��
P2�T�z���Fm�Nmvq�H��38�he�s~� CQ��d�Z�"�㯮5�T�xI$����cߵ{��'>��@��q�e���[a'y��,u���kOPngz7X��!�O(��D1J�`7����#h�?�$*꛱�y&�F����qv���ߑǶ�������rJ)g������t�1�QmPD�S�V��;ʑ�����eҔp����a��v�	�vp�g����nZd�K�W j�R�Z=E�	�$s��_Ҡ'��D�*�#pu�1��b�^YK�3�b�
e+xG(��N�����/7�G��������WgUN��z�Fn9�m/�=�2�+�節����
7{�[�vN�O�A���L-l{*O��uvN^TL���~��\x;_������mn�I��얇k/�.�^�����:�>,��/]��[��Z��"b��oFC�Ɉ�+��=s�����%�DH0�}7Vܤ���w�@GY�aU�-��.�!D5�Nr������y�gg�p'Ze{��ra���r�p���	�g�g6Ի�#'��D�
��c�R���mJAҴ�
�?����|�H�:1R��h�MBW�uZ\k]��e�����Ck����))�����Z[���J.n���W����`5���ٚ��Mej�.��b��	y�:e���l6_n�g$#��ئbv\�|"��W���e8ZGUB�:rܤb'�@ ���ސ-�?��?*H@ǁƩ�F6�L��L�&35CWlF����|�8Km�ϥ��Č �hX��ك�!�+9����6��!=W� ��Vu,��)#�|��5-��b�;����rWtn[�]�*'1i�"pnߦ��W[q�y�3�O��F+U���jx���ʓ��Q������8Ufl&r]�kn_���;F:����_��"��m*R֯��S�nkװQ4�<œKHy�xX�]t(�(��)\4h���#�ztr�����C.d*d����8Q����T
�`�td9���X�k�^��˕��؉P�V�Ey��ǌ�����<���昫rǆg�b0�\���!�|�h�Y���>E��k@K�� ��Q�^��|��dr,R�66냫���o�\��R���u�<�B�� L҃��g�}-0������z�1�'͘8,VC�D���պ���}�e0�{"l�9��V�X�0�Ա��Z@�æ�5M*܂�l�S��!ᄛ�7�2:�k����� &�z"��.����a+ƳS<�O���/Z��R�uY_�����4X��(���i��(���5��M�=؍��$w��I&͌XO����g3���0.M����M��G4����aQt�9=W�b���3�D��h�O�eq�=l�;T���aތ�٬}��MBM�� ��ꑙ*� j�T
��eɤk��Y���zs �dTL�P���Zn��HN�鰚$Z+:¹e?����5��3��%�d��U��Ԝ-���mr7z���~��$A�J8�'����&~��yw"V�B�)>^B�mL��(C�s��ٞ�%<.��z7���:���7�	?���V2ĸm~
��+��{s=�4�k!�h�(3�C��g
���`k�RtG���&җ������m&����bĆ6�M'у�k���&h�D�B˽��y�F'��l�h�v>�\��n���߶>���3o�S,�
���νT\XP�	u������nzVi!��O��x'��SxMo��̐#͇���xa�A�K�3qٷ{�6��Fg��-qR�s3�bF9��(]f���b��@�8��@ʕ-���c����~�DN��u&��|�?*�s�9A��+U����ti�0O#�L
��y>�EH����vڟ�`q��C#����P�A,R������7�H4���=�c3D���9�O<�5K�|O�3��!���=���VM�ͧ�\�Z�H�(�>l�mv ��j)R�:���tCu���E���~� Tn|\m��$����D܎6������=�:������
�v�2t��M1���;����}�{��hN�XYh��3���!��z�Q����x�G�h�z�H����U����3��Ū=���$J����t[�Ǽ��1�� 5�6q;�pY7�I����5P�jw<RK������g��Jɫúy"r$je�c$0â
y��(��4S��x�k o�p��/�خոz8��?�Ͼ�1�F����5e7`ătN��}���悁�;�BGO'da�/XQV�z�����5g8V�IƱ��c\��Hs��S�@��W�[s6�NL)��G�f!�z�6���\�J o0��*�QH��iJ�	/Y�1/��tR��������b��2�h@��0�ң�cR���6.جG
�Z�H^�7���`�X���n+}5�FKe�{��ہYR�t��߭�/�	�IvtܶxE��fܠ6���#�#�H�O���oD�$�!@RZp �ؘ�^���%�7�/*〱?N��
����k-���I��Y��(ƒB���j��.?����0���U�6���՞��|>���XaT�M�ϱ ����<p+%�b2�䣥2���>A��ז�igS.Ĥ��t���@�T5��Ĺq�������#�r�ʱz,�u�CӠ?Q�^<�퀋S9�1}��ʤ�V���z�@�})k����#��֤?H�t��$?�=��.�cZ����'\��W�Q��P]TS����\N��񁂯�ok�%L�y8��ͳB�����&�D��ĉ�x^S)A�8ׯ�Д�N/�y��m�Ь%1�&5�H�~��Sв+��7�D��J�ڛٺ(���R�'821�rkL���D�D�̠��p��C�6��M��V�wWCbL�-�7���	�|)�mѱ�H��,��$�TH���5�Ncx��Н]47��S���iV���ړ�D�X�b����n&��c,��D�D�mU�'fs�)�75�+-���l�poDf(K�9z8'KǓ{�p��F�Q◵o�6�����_�I�}�'.P��k�[�����V"x�:�2�5���'Jv�yg�[�Z���}r�$�ٯ�ئJtFP��& �$�sc[��_X��f�Yf^m= }�:ږ����$(���.���ˑ�9�`����^n)N�4d�{]�ؚ��������瞸���x��Fiϐ�qmhJW��;����(�;���=N�C��+�X�'06��������ѵ��yYm���M�74�R��%<Q|�a���t���1K�\�&�ؔ�6o0����,u�ڭj��{`f_��C�4��s�΅��\�w(p��5��'W����%a��3D�.Y5%��[k#/b�E`xՅ@+F�ˡ�]��	�u���I�-������]u�n.��dE�4�c�
%![����{�ku��!!�}��;Z�?l	2���G6.V�6�i�,�9�J������]���\�>�l�`�0�i�YRoԸ�L�--��c[UE}0�	�"�/ [�S�}�A�]�C�t�T��}���G����0���R׹���-
S�6t< �uI��q���z�\6Q�"Z� ��j�����g��$�v���&�n	��b;|<����¶uo��\'
��m��>���J*'�7�v����XM@��u��1��`N�I� �v����`ߙ��Y?`֫��c�c�~�Y]�j;f}ԋ�(/������'j��>�_�/*���'AQI�є�W$��,c�N٦qM��� ���;�N���9��:��2g��V�D�\ڬƮ��\�W���!�k�q߹�y���NW���%�1j=XYE~�6�q���6�`�C�F  ��q��K�=����s4�Y� U)y���{^.��*.Vk�r���z���]�c���eٵ�29�Xd;��B?�_�y���{�1��]�c'$W����A��y��^���������&\
�J�e\hr��u�C��,D��v�U��@5����H�]��Cz�7L�O��۞5��H���`"
�<��ؿ��ٖA����HV	���LN����}C�3�Z��o�.�<���l�0��^ؿG
�rF˘��<Ni^%N�#���̽�]\Fp�"��&Jw�ี[�y�X)��S�x���e��5&��=����l-��,�R	�3���<��~o�N�f������̃�o ��r���n�w�E3�TՐ�U�����g.��,nqA��+;;rR�Iy��]�}���U�t
\Q
CC��+�Rz���U�ܧ�'�`M���_?1��̏mR��0���e�_��/�r&���#ǈ����
?h5��\�H�:��6�	��S7�[{4+���=���2(l�!G��Id����"�z�!�!|���$o-���l+C�Xg����d�@�K<���^:K��T���}��"���YiVHX�<�S&��g�_~Q�U�;@"Z㱹�(�ۋ�������L�8�i;����}9�;�4X��2A$y�
I]�[*tt6��e\n�� �fU�(����zVa�� v�!7���~���5�Ih�e�p,Fj�;Κ��^t �quY���E��J�g��b�Ȯ�b��Jw�cp'\*^XWL!��dVٸ��^��[<�x���1l�(���UMV�h=^,?c��t,=���Yi.1%cls"�*�tծ�<��"t@+Q0� �j��{W6�� aYk��-�K�D�wO��2���nU�XP��§������M���}`L1����ay=�P%�J�� �3E��s�!�{��{e�1TmD�9|�G�H�P4�䪣��!	5 0���:�Y�N2�[eH�D�o���~w�I�7������~����9�Hl�0�h��6%%��TQ{�<?��@b����uI�:|�z?>���;R�n)��Dy���v�	-�&s�dp����^�:!Պ��x4�P�.T7\����;w�k8���(����&�,�]+�<��f�8�x&_S<�8�?�A����:��e�}S��#��{��D���n���τ/-�U#ve(e�������: 3[~�*<��c@�l�=:��0�#n��Q�0N���&�Z�j�\d�g9���D�e�E��I��e^{-I�p� ��7{~������Mhp���ѣ��t/�P�Uu��C���
<�o�Un��_�t��Y��;����7W�K0��OR��h��:@��6���P�(	]�n�N���b,J��/�'w�@9D��V�-��Ht��L�( �Z>��%��Id�����2���RdLݤ�!�O �~�`sK�Q�=*Ǻ�q���l݌G?����A&>8f�愓��0z9���/+՘��($O4:�C��/�K���׏~��C����l��|�i���Y���	�(�����l�	�%5�����|s	�R -H�x?�{����>�C��XH�4��4yi�>)&WD��r~C8.�h��\�����^���fpp�uh�&�S��"x�h�����Ek]ߌ��l��2��-2��.Wp����\h�׭'��N�c�}�REi�;b�~�-`����bCdn��jd`����jj�	ҊH��/��y�����t�	D5��O��gA��n���n��t���K=�����n4[[X�B�֣�|Տd����f��Fq��7:։�:��f�$Q�CE`;�VA>��ugG��o*W��5	�I�3iq7��X�Z�0,zIF���.�I�RJ@�2�y~�+�u���I�|lh)+��X�i�. }׵@6��4UL�,y,�ܨL�W�g
�)���o�n�	�h��S��ݒ��"����w���^�3oD���H7�f~�]pP���ѡX��`Z�� �^����#cp+O�	0� ������������X��'}W�D� �lN��AZ�>�ߓ��?�y��K�
Q��/zĭp1vG?��h��4����O�9�n�>��:Kx�����8�+������e�-��vԬ��f�M�?�
u�N�LEXֈ�%�8Z^(��&&��i�?p4T�]��qH{�Aj��?ȳIl��O��<b�8\	=	jp�4)c�������_�Eph�vc>��>�J�N�wB�їI�Jv�z�DB(u{����(� �L�Ĭ���*�4�q4�L,P�����bм�G�B���}~� �1�Q�z\���gz��M�ׁ��|a%ԯh��<b��ZO���eR>k媮�p�E���!#ӟ��o5�F���Z�,{�g�.�ISi� ���X+��Y��{�*���I?(��&6�g�����W, ӫ*'���D3�Ԗ����y/�'-*>��O�K��P�%��l}�{��>s�Ok-�C+I�����h�;C��i���!�b/��;J���q�����_���>}=������jr�X�8��կ�y�&$�'7	�������AI���bu5����Rx�S8����o�R$��bq�.^+ϗ���^F�w3OX��P8�����$K?�ўDԴN�=�"�/�|�>-����K�lD58Mk���I-X0\��eu�\Oc������(`}y7��1 �����q�9�g��@BY���{ЖC�ʽZw����[H.����_��A![�Na/�v�9�e����ւo�/��M8=���>��R�s�.MĬ���)��0!��Hޏ,<���	\���I������_tOp�We�	�FD��>���a������Ĉ�%��8ovPe��bΉ�V^��b�(rY����fw�`)�"����ĸ9-�\��K��U���ȓ��gr�C3ˠ:-�y�N������������AX�&s�����>���Qe�zm[�(4Ƴ�Yժ�0�,4��������$D�a��$l�������B�E�I2��}DSV9��u�������Xu�-��0���:��OC<�w�d�����Eo��&o395��2��K:��p� �~Y�c�F�/x�'���a���)ޒ��������(>�|�4�T��7��"b����|����1�.������]8N�ܥkJ~���';j�z��Tp�������e,��PE;,Ĭ.�>a�������'��)�tAgAs�7���4���}i����P�"S�yr03��6BU�)3���c^uc�����2�>nA��wNA��F)��`ʹ����rl�����mƗns,�X鯔}t~�oY)�v9�$�Z�d��e�����a��+׋}&�����k�p�m�Ov��`9�H��C�:<�f����-��@�U�ܻk'Ax����tuC� D^n	�>.$�C���#�ƕ���rkxe���⤣r��qn@���M"\�qO�7��yB������8�n o�p�\]�G�-�)o(������tds̞��1@�kؔ�Q6s11S��!��D�~���<m�Kr�r�0�X�dl$�.� �|�
x�l՚4AO�1�@i��I]׍pH��(Y����d.���$g�h*��Q�*:ّ,��C�{i�sļ�~��]DN��m䧆�;��
t�85�qE�Nڬ\������l���'��~�	̹��2�*%��'fQ�O�65 �"s���r^C��R�V�W����g�Z`���t%@��@m�Wb�4����,�6��]G�	<��՛�����R���>M��w6���4�~虦-g�aûӂ'���l_�M�&��>[QB�J�c�xz۷-��~ ��`�~%�6�G~��6�մ�P��^�c3O� �>}"�#x��v(�|;%'���^�Yj|(+�k�:oWn�uDdn�h;�z4���]��Q�k1�hdQ�y�;M�O����:��^�Q0}��̿����3@�N�M�ǾR�fFC��l1P�t�{���>�f�#�?��y{=�����L?<Io����4�:.���,N"hwI+*a��;�)r�!����\a��AMnT��L����?��I�+�L���F����$�4�g��a�Q��� �b�2"Fh�횩T�5\�,�9�+���u�I�"��{ן]s�c�m5�2���(�y��ɧ��69ѽQ�=ݯ���<�-��B�4���DO/�
�G�;y��}��F���=e�	�620vsq;�;i��Ǭ9M����I\	k��C �z���.Ū��OV�N������χU9�1����K3�5�����g=�M+l?JJ!�
$(�ye��q�V��Ѡ����!^��v��b�k#B���r�ŢL7\ę�1�J��xY���63���$�S�I*�{�~�Kw|��I�wKv�'��F�Ҁ���P"ۗG&�7�H����֯@ήL�5���=yy�g!a�rS=�� \m`c��lS�V�����$����%G������w�6*$�S�zg _ZL3^�#����E'��.,�-u5fS�?��5����x�]��F`~`�*mj��vd ����B �ٲ�	0���ύɂ�=s� ��x/�����XɌ�~�&
B�(�&�dѨ!pd#��������Ǿ�ifӝ�X�D�{����
,y/�Z~�z��������ћ�&����&Z巟 B�����ZL������Fð�ӎ�"v�	��M7�A#r���h>/�D��exP3��7�Oj�5`�pL�r�����&�
Fu��64bZ�9tSz@��T!��Bc�-Ů1������iK�����)��ed�cNP�V\-4��k�)����sz ��f���
{@�-3��  �x��"�}���\֏�&��gN���li9Y��//��W�sg|]�5'm�;��r��
�Un����Τ��A4����e��8;�d�������Օ�f��Q!�9/�����Ǌ��V�7�����$��Y � �Lw�[�Ip�C7��8�̮8������@Û��bW���{�#���.�6k�_y���(���/t��$�7O���~�k��p=�Zg�����P�aF{`da��� *���C�{E�F̹�,�ԇ)�JW�+��x{I�t�*��D��B��1�vH�{���M�eh)#��vm��?��!ݢ��)"Ș�����Z
�W������FO�d�xG����� �Ұu(�O>0InL�����p�V����>z9���]d�|��v⛍WV$��?\o�p��6[�9 ����ޅmKI+qc�΍TN��jwR��˸PM;ݛ�5=�P��]�I�4b������AY�Q�P��E�s��[Uc �9ps��aajƳ���`���v	�B��0D��p�@2$���p}��=)�Oe;��4�WY�g?|�n�S&ϗ/��w�3���R� ����sRSwHĉR)�d���̔7&@^\6+�\@GQ�_W2K��!�̴e�R�Mb��o��:"KޚQc����Y��o�
w���?�98>M2m��Z�m�B4*�	�W�>�������J3�F.jB�+o�{*.wG
��K��J��������D7���bAo�%/>h��AP�ob���J�W���.76o`^�g(�x�-�?�����V3*E�B#a�ghY�p%�lE	]ή�I�{~�����7��L0�}F7��ƶ��+�vؤ�s�b(��r<����,s�d���?�v��|�q�7������eQ�VmyW"��N���E`����O�E$jV�Ԩ�J�'��a|a�دr�P��e[;q����栍5��Q����8�tB#v��׃v�-7���{�k��Kq�=�ml��r2%�z����<�t�:���f8N��Z�"�B���m������Pz��ʹ��}�:��I����Y*K�(�4.U�WN�LKu �]&+��}eG���,��bU�{�:��S*�+�`���©��5O��I0�׸?�BI��C@����K���>TΜ!�f��v���{�s�'��~V��� �T�!pb�&ѥ�ՠw�����i�G8.��vv�]],ݔj��jtf~��򞱓�:2�FȻD�1�F��7[_㼽�ҡl�����aZd�[&�S�k�~�F�-ꔈ[ݖ�D,�v0!-�6�*�W4�>{�m�	aA[.Z������ː6\[u�L;��}sS*� ��	`9�}G�md<#�7����
��\���w�2Y���(��B9�?so�����g \�Tl��o���w�`�	F�~���cIgoH�����防�i#���t�﮻���ѻE�h"�qA �q��S%\4�2O��y�d������)�m��h�����`�k���dC�z qȖf�Nۭ	pL��?^���� B�Q��{_�&��̢����`�>�M�f��wā��c�PNڷ��:8���2�FZP9t�v���t�?}��1���#,�+8��>�^�J{8*6�����2E��B�/VtC@����#�(~Ҷ���郠����*���t��fT�rY}�|p��{��i* �Y�{��vMs+d�~������M�\�h�����6u,U�v���'�ϭ٫-���"`��f�����ᾚS����,,��d[1�v=���b�p�}g�A:Mh+��V�����SN㑚�e���md#���(�h��|��=����w)�F��UW�ވ��c�߇Z
���s���=�E��G�}O$n꽰��dR�Y���QjҮ:dq<4yD��$Uܼ�s�xiVq�E�cɜA��bo\wa��IAѕ��Q�<<%�#ux6tfh#�&N9"��^v PΊV�t�]9vd��e���Fw��c%�a�)�>�"��	a'�Ckm\� �@B�Zǚ�A�Ri��h��9�D'z�ϛ�m�ۧ�n��O �XX>&�_���P2�*2�Jv����bl)@n�r
%T��'��
��į{!���ltmlC;;�P���(�u��w���f�ע27�ZX��܎�:�����] ���ʽ�X�j���h��2$�p!���Y�ҳ��"a�Ϧzj�{P�Cs�=3���L�7��Z��K�}���=/�`5��%<�=t���'	ڃ��Qzl3��>؉�oIhܫ�(w'�t�?�>>!dG�3~�5�{Ybq���g� L��`}���@�;˼��dd�� ��g�&�9	#�l�˔}=dk��_e�FR����CK����oC`\�����O I�j�KDЭ��՜�2M�!2GnO��/�{�Q�9R����\9&�x�q��������9x�=��4�;5���ZvϞIN�;�L�R��}�fH;�Nl�ߣ�}
:C��OZ�j-�=�7ޢ�D�_�(|.�s�����խ�y�@^q�K>�u���|���_N;rNϓb�fW�R��,z��/-�S�|^��*�P�Ki���Q��T�<,G����u�v�i�xm~�Fꆢ�+m�He�s掔���Z�nٮ���*���u��^
�l|�=����u܊��uKyB%:�G�\O;��kr8&ul(�̱�����Y�}2[� ��#�fĴ�f�W+3]�� +��%��@N����`yB$w�Xu�[��5��K��b�������Lժ�[�~f{�P�i��i��a�j��K3D��m��D����(��7M���J�*F5�6��w/�֝�y�-Y	cL�U�$��3*����~��j��L(����c"Q<~R�8�#2Y�_�^����)�$*�� =B�-[o/�v�"W;|�����a�'�~na�>G�������:�3~���dr�� ���T^�s�2�7	���˚��.f�煮[#��4���������%��8Á`Jpt����bHB����/���Bcn6"��7e��#��Z��/sj��k��Vk�[ʮ�υ������9ҭ&O��f�T2e&�>rڟA�-Tt>��9�Jg�p�6�Ѯ��av<B<�.$����fw���d��3N7�$�e�{c�/-*�zb`1;�e��m1T��2�Bې<U廚���!�8��?3��唚]��;O�fy���R�K�"��"������u~ן�m�崪D��}\�d���%���Վ��J�:��<�loa��>���B��ԽW�
�:K�NUߑ�"ӫt��� ��Y�vL#*`C<���X�����y{ e��K@�Y<���Ɛ��7�>m�B�=pp��{�Xz���+g~�;������'��c��IJG��\SBo����M�b���)��������)�o�f��R���C�x�?��3�4ep��'�������oU���6u�69��Q��ؠR&y1���}��fb��v0H�̂�X�b���y4q��'m�T&|�sݜ�v����o>'�󒛌G���a�΂N��T�򁈝��Ç1�=�-���a�>k�,��t��Išؐ��`%l�v�|][��F�*#}_&�
�x���m�nh�'�kŅY�Yٷ���;'�i	������&�ha[�]>�y�J��.Z�\��u`
��`�2.�]~t$�D[���2���G�r��-w�4Z `^�{�����;o*0��T��;en���r(8��=3c-��Mt�*jpn��Nr�[�ITФ��7cL��^;yB��!��!���spJ�i<>:�5A(/�e���ع��L7
��Y��Tj��Å��*ۚ�}P]� ZQE\/�sS�&���8�r�ů�{��˫enU��q��?I���=pK�4{�f~hf��-�Ԟ��3�V�燎�-��eq���@*D�Ưj����gW��M�t�� � ��K9�Pz���m�#j��n����e&ܞ�|��>��35�J�v~;�SM��i��(E<w'	:;��\�w"���*���dK�G���[;��o�+ȕ�y�����h�uv=���H���&�7��,�1_��Ob�ײ�mɓQJ^�H��ǈ-���)��~�`
�߅`��u��h�}B93�b�F��l���6�����R��IѤ���X�5[<l�Ʌ��~ȡ��w~��tZ�Ob-�G�U���E=J@� K)���\{��bݬ=�{�X;�s]�l�ȅLx~�Ny�`
��K��7U֒E�C?r�qZo�$_9(;��3��cOY����{��8��τ�xdl��]A,����h`3(�Yz�փ�6�{��`�dQg�]�r{�HP��F ����[)(A�65���$�[��5K�1	��xHS�PK�d:�	�Ui�r�9�u�G�8bY���{1x�_���C�6��i�ч˱M�۬��b�f+�+(t�}d����s9\��L��׭���.��6����� >!3���sY�frw`2{2�h��������/��:sMY�S�K�;�l�Y#Qad�3pt���[�	��ǽ	7�ܔ8�!bY�l�a�bv�6��`�%θ��z�<#�c��lv�K�Е�ɵ]�����y�������.+��I`wͅ�ra�Q+�S���/�8��d���&V����U�w ��8揀m� �f"m�=Uv�5Ѫfg�N�Q���,~U?.E����!����]���>-����+慴��m�S�i@b��-Z��WcI�~�3�BП����`T����:��WQE�E�wZ-��ζ���Ў����$ӗ���"���A�rX���An��~��dZ
�n��@Ξf#!�t��1��Z.�ܓ�����+�7��Pω� �Jv��#1k�����ЖnU<캯V��Չ�,��?��X�l���>�'�BS9[�x�\!�oWI*�8������>�|�ЅC���a�ą:����0�	:5k�Cc�p��U��x
�!S��k:�\S�ĚZLih��j�g:��%7O�3��>P���h&���_�u�9�eh20�Qi/�9�n��][!��%ě1gRO2����&��xrG����^�V>�ѯ��1v��C�s�#˯ט�/r[/�TS9�R3��H,�`i�Dܙ���"]�ي ���ԩ�X�/Y0e�D7τ�8GF����ᦺ�����CZNO�f�Ҁ-��i�߮9�4?oC4F�m� {�v�c1}��%fI�|bϠ~F:��fZaN\hs�������o��q>f�֟����8���>7����9�%�?���)A�V�%mg�P(��5�ZX�N�]!�e I��E�����0Cf`T�����QE��k�,��]���|�&ko@��@�oك# �L�����6z�v�Q��v[[��sRm����\N�����������P8��{��i��|�u'�҄��ܽb�s?0!Z�	#�����ܷR��!-�vM|tX<�VR|xe�ј��z����0	��F�R�~�3����Q��;��gɁc�(w�ΖʁO�	 ��ؖ��/��2���M�W�|��	�k��[��A���qݜ��55"����K�G����Xd��|�QV�E�����&�8�H�JF����We�M���9��{�_>�e�����;�O)yV�Z=J(�i�VJ��}G�����ʲ�0��j�����������`�v}Id�ɬB(qث�/�}=3�Lëxe! ��E��Xߴ�@�
o*Tk�����;��5F��W#�����O����lg����w����U>�mQZI�#	�R��t�P��Zf���o��2Z�~wg���4��ƈ����+ɯ��+j��4�?F�@�C���/3*�f��=�H��攅����,Rd�a;"@��/ů��o�A�m�0�)��h�(���%`���c�4��^C��ڀS����|�I(i��^�����j����\��./��Ġ�Q|�4xeÎM��� �����h�����*�,����E�H�i�d OP�5>�G��� ��,��}��m���K�"a�p�HK�;�ĝ���{���V���m7,B��g�9�}�#%��ٯ�}�Q(�nl-�$�A7l��R�{\�p$��N�J���좶)S��F��&"k��f;�j/�͡PH(��+��w��Z���L,L�JJc=�p���y2M�Wܸ3�\����^�k���"#�G�tcE^�;y���B�	�"}䡤�� �c�Q��F:�`a@>�x+�m��.�f����z�+�e-�����w݀�S�-@D�9 ��b�;S��0�m�u[� � ֋����n�/ص��Z�#�/�;���.LFP�x�s)�v���>G��#�� �.c�!�H+��ڬ���+6ً_��m���}:������=�%���QNrX�zoIr��B_�{���|* rۈ�ro�?L"�4��(�#��<;.�ި���Ϭ�l8�EP�;\���JI{��z)x���	ޕ��ܟpL��@��8����Z�7b�*�xf��iZ���Lڲ9|��ND��d3:P%���4�{-�X�Y��W��[)!H�1��Qr��CAYK�q��m���Iw�D.����*�Bn7�@�N)�	�f�u��]���b��]MVΧ(j���%֛M��k`�g�e����D����<��ZF&��ۘ���9��@[	:��HZ���C'_���XD��8,�ζ%��dj
�ʶ��;|W�H9~k pל*�ͭ|�o�|�a*b���r��ʯ����b�Z��LD�Z�\����< ��4���p��T�p�1�����]*9�'���̀{�  g$���:�6k�ldP��`�(��z�H�\�ߛ����l8K1�!�feVß��������/!;��̈́�3T��
˽]���r����o����{{��^��Pآv�wz�3E�Sȵ=�	Ģh�_- ����2>�&�_]�����
;�L�h�u�9ȟ�K1f�`a���?���[52�t�2[�;x���X�쾣m��A�ĝ��j��Q����cl�L��3�q�R�b��X��	?�V�d!VF *�u��̹~�W����s�P�N������߂�/sBa��I-��E-� >�"�KaC{���f%ڳ��nn��;�d� J�f�ʹ�H0���� ��2���ȡ�wٽ������N���������q��H��*���~ذ�#�]����ч8)����Eߖb�)t�>���E{�|��uˤ6,`�����'�,��Ԍo���K�ݧ)EU-G�[H�E x�$���%B��k�	!*�u���Qx�{��")�����>/���P�ևu��o������d�_j����]�>�j�[�d�M�M��D0H��+o��zq0�X�=3�7�C�����li���γ"}�a.ُ���]���c��:9P�+VE,s��9�"N��qL��[���x��ˎ�֣�P���s���ي�X&��R�nւg�:B�ؿ�n�nx<�2����7�$<��-"�p�O1O�3w��{�oߒ�m:��F��c]�-Q����T���:��L�>�E�N4�V�Xg�T��%�>��p��j���:��7�M�L�ƍP��d�D
C2R��ţ<ʔH@�A�����Qi'G�1�<�\jJ��)�:
�uH�?�S�j���S1�({��|�(�^(@��;U�pP�5QΓ��i�+s�2y�8��&Zz*�x?��Fe"eOk`nk/6���Ј�������t��2;V���ԍ{�ɧ�Tt�� �F��T�PN�]@�ͽo3�<[dܨ�<G�<=�4�p�5��YS�xg
���^�f���.�עB_7չ�GSD�:���U�	���84X~t�vǾz�5xg�(�@��&8��=(2m�TS�����m�d{s)��7�v��L�����3����B����ā�;f{�}�r�|LD�� �!D��"O���88ޱ�r�M]F��v���;�630`��:5%ly	ԮS�y�Ț>r��<��Ƈ �^��@�'Ͷ��<Z��i���sm5�.�jո��`������^�J��Į�6���ȐH�֧E,��\��L8��o�ߐ.,��[t&#��{�|�s��qBz_�,SG+��)��d�y���_F�%��C�:�����c3yd�Dv �jN�5�ݓQ�k�}i�?S �җ;����`�#'�nő_�ą>	s�8<gU$��d��
���(K�x� �*ֈt���q�h&2��~�ǝ��,g�s'�F�(>BA3t�a#U�t����t���"�a�̼C��-�
(�� >߆���L�ܰ��y��������h�E_������-44�p'Mɔ:����A�Z��Y��]���Z�gM�������+|̕��I�*\�3D��G�YL�)V��I�L���(C�y�����,SH7�|{!�)�6�E�2j�� ;�<����O��3\E��D�s�[���P�k0&h }�=\r�nS_����N6�i��C�0��YO����#�B�O��ˊ���Lnu+mjdO ����O�T^�_O�2�~�pP�#/0��h^@Һ�Mֹ�@�6`�[��~��μ%~�D��h��E۩Î��k���3���]��`b>+s���~�M���`��*��Py���ǈ�)�ɂ�t�@�1x�|�?�Cӥm���S�l3X�.]+K�6ֵ�����w�V���۔pbw���Q����&�c�4�P;�ګ���`Z{�����s��I�y��f��j>j8Xj���0�<:}kSRE��e� ZC��e�k���G��l-����� z9��D�p� �Z�������ҷ����?�%�'�f8�w�mݪ�G2��MW�*@��b D5[�o�m�_��;��ٔ~ȟ��S�T�`AH�˚$|�-24vR{�N��5�Ѵ)���Ή�^�����B�?�ӧ����5�,+�'��j�,��l"p����)Vf���Pg=4�'�FM��|������ b�k��[�?x0���
WC���h�����;��6ͽ��hs�Im)�F9�>���"����f�J�]����u�α��=�I����Sz9p+{�!}��1@�W/ý��}JU�y�Gf��o�h�iikA��4s�����Lz}(j7^-(�Kɏ�}���W ��֞b9���`��a�(�5u�D�<�Z8�׉N��YU��m@�&����A@�9�u͗8�{W�P���6S�+����{r�=��e�x������_�/�+%���/��0�8{躕9,�O�v&�,�&�����*E�\�Z��8�Ty�gj��"�/�I,;o\�4��O�X �Q������a��|�ҡ��<}�~0���w�W����L!k�YA��c�5=I�F�k=\�Q��چ�]s�� ��;I"�5�O���I�B�	�R�K1���6w���ϑ���ˉA5�U@���i���W��?{��`
sM���?�B�b������No����ݤ&���T�vsר�˼�iP�4%x��T/f |{d�X|�X/�F���@~�e����L��]߀�B.�Ҩ�1�"	�p�o�[9�te@���s�Y���U�>�[������2~��v~פ� �.�ς��2����MID� � s��U�O�.���ĕ�7|���`�Y>���PL�uƢ�m�Қ�&Ӽ,���{qE,�H(��):%�_�ƚ�;vo�
�1S�����	w�nqrGgF�������XI�I����m;��d�m���r�Ԋ���B��S%�4�i���_l��S�+��Z�5T@!Q˽����� �aO��B���jD��`�p];L�1�m/Ok�A����k��0(H���^���.��~�:DR8�0��o޾�H�{�=�e��3�&��2M`^��A�uV�+�H�	�"�4�	O�D;�٪�Z7�D�ῙW*��3�����
�rUN�:��YNsz}i�>�4�|���O`��7�VT�O��D6P��K|����G�D���<b*�� "�����.�)Y;����ɔ��B��D`�5�$[�^�|�Y>QǙw�/��m1X-ٴ�u	��+@Ej����2�d�����=�����1��p�D�0�S2���\�����I��v.am:H'�3���T�� 7|�Ġ�\���Lg:^"������ Z�� ��$T7�]�����Yo�f�'ֆˋ_�k�u⑜_������OqBa�T�2� ?e�h3c����4�gj?C� ���Z���^S4x�_��&b����2��X+7|��x�O�!�ԁ��
��\����cХk��:�-�@?[Y��m�ur�i�7<j�˨�K��5qHzB�8���W��}j!ށ/ ���Cǫ]e�cp�#��Ys0�Ks�Z�~_�2��:S���#�{��eD'2�{�0U$�����>q.�;~�(���9���o"�*�pBچ�_��8Vu.���������5��_�(E9I� `�P=���Gn�+c�E�?�SM����PeD��T�6�{�L&#�0��.�'3�dK�<��0?:zB���u�\�[���h�0�O�=S_�?���~`��`M����<~Fӫ�ur|QՐ��y��������+�N��j��ʀ�p]�7����M�%�����ٮy+f������j���EAK3�d�3&+�؜H�JO8�X����5'�.�<'�O�Э�܋{��I�$�Ć a1G����wՓ��ȫ��������f�$;��N�U�׷D >�!9�I;p`利� #$0�Q���,EY�Zָ�}���Ct���k���5��Gv��_��ӂ���	��Sc񆘖�QL��I�J_i}W�U��	F��f��-?zQy҆5)j��ц`l��G��B@3�y��uL���x�Q'�VZϳ���Aè>]�0.���3YQ��":�tX�ĵ��.]���a����W�;�٩I�m9��2��ȼV)�Ӌh�[��Ƚ�YA��6�E7a�C�T��ի��ek�1q��&Z������Δ��>G8�a��}��o�J*�Qr�y�@x�DE�%]�1&Ԛ�炝cԤ�+k{��3���-;��� Q��ޠn�Y��6!�_���'M9ζ�Y!�w1׾.^t�Nr�:�ՃSU�):&�d_���߰e�u��SA�Jj�{|���1OXg��q(�8�;0��W�e�;q��� r�])_����Q��
Q�9X<WF��++��^�B�0�j��R���YirU��n�/%�89/*%Fu.�":B-�M0�A�5iz�����
i@:��0�v���,H[��y�	���w��7cTl'iuՕ���u6����ʽ�ZA�F����`� J+n��a�>cT| ���8'�8��a�b8)���1X�e�����[5ko'_������-1�9�9Az]}�%�£����z��u�O]�#�,��g+�b��Ë/,T�*̈́��4<Z�g+���ͫ�V%ү�Y� ��*�Y��T�ڽ������S�9�����(�2��4�:6khY'G�
���R���N|�G�)���������e.&�|9�b~Q����T.� �J�d��\B\a4�����Ǭs�*9�^o&C�	����RD����arK%����(	�^k��Ѓ�U�q�n����e�:����U���������"c�p����Ϲ~�f�Zr�X����-~N��(RE���A�p�8����8���zԉ��n����D�<L*�kO����敉��{�\�o��D�2e�&�,�ǂfs(��Ĭf����;��g��Ou|GK�~����S��G�H�L�|�EA�$� �on1� �LP[5蹓� G�Z_%�����0\I����\F��ߣ��3O�L�pG�j6ў~����Z�� �6���q`�8�U�������@�Qh�Hǚ$\v>�H3��)�y'����d�moy$ӌu��8��vb�"�n�|Ƒq<8��*�X�Gc�) ��"�SW����5@\_�z~R3��a�]"�o����� ��y�\\��)R͑͔�w�6{30@����MQ�g:)l�R��<�-�?Н�M
��HT�T��o>6x�����7!�V�:����"��^K!�xב�@�:<�PGIdl���k������Wrsn� "�U��꛷�F����Y6�*����ncu}#���;�Fd%M�ȶ]�ީ�J���-��Eo��׾G���m��� ����J�{w�W���>Y˾u�lT1x��4C�=�vT�*곎�Y��HOC��-����{1(��F�OY�KC#Z�>?#$Z8eEΎȫ��E3$59���!�Ou�	�ْT*�Q܀Y�|3�,�įyw��LgT����\E����m�U@%Z�.�(�j�7����x����<g~��`1��-�A�����n?��h������=)*k��U���0�O��/(��zu>)�>��.�/���*��e휁z���ݥ�&ѥw�C�sD̈j|u�kR�5}Ō?�yG��,������U_���/fe�����>��D�[��T	�=s���cg/���q+���G���p|��v��7��w�ɴG�zĀ.F^ʢ�*��a��0w���j��L� c����J��7�Yx>U�<`��f���䯈)%�*���Rs�Z��d����MI�l��@_�-za��"��o�	T@
C]O)|'�O��9�h_�RGs/�ݡ�8��Z�5*���3yꆻK���9y�u��޼�zo��w�3H�fMr��L~K)pb��0����%(���kq�l���t�����y��䱹J����f:�Sl�۶3�y�����|���	%��.c�ΌN�0ӷ�C�`,���X(�V�1��Nx�����P�AW�e,:h1;�2[�L� �놔�vҘ B����c΍�J�E�`c��&��� ]U�vl��>�jn�p��a-Ds̰�0�pH7����=pO0�7N,���ß���wL�Ɇs��r*$u��R�	Oݛn��7�I����6���{۠���OQ,j3��CrH�[P4a�i�ʩ���'��w���
|HYם��И"��97{��Ե�fľո������G�d��1���q�k֡�h@e���k�˚�{(ĉR86�f��Q]��j���ط`�&��x�sZ��U���9���`WIs�ڃ��!,��|b�B{��D��W+-�P���s�K�Et��Ѷ"ǔ������L?�Q;O��I�>V$F��X�^|�V֞�=aW]�8M5�����lѓ�a�r҅\��t��el�ch&?k9��	�p��F6���9��\k��u%�����ZT�΍R�����>%�Gxߪr,�~�lV�,gg�he�Uzvc��U4�R(^$M]���lz����?Q��U��^L� �B���O���%�g%ԛ�Y��q��tR����mV(��@��D�L"��;T���ʖ9ix�pt(�w�`l1��\mZ���dνSg�$?� �.	(F^E���X�H�`��u�Ջ7�c���G X������cg�Wm�c��,�6>-N?�h���H҃^�F��*���xRW6��9Ԝe(e��m���m��,�.-p<��$H��5VS��\�N��ȵ���
SuY�^n���b�AF�`�L;�GS	�M`�Q�>d��w�t
[l�W�V��;��6ZS{�Õ�u"�+Lʍ0���0kL������Ղ� ��1����ZS��y�N,kEA,挛�P�6oj��p�R?��b��;�)���o�k�`����ٽG4�P��hi���'pJ���3��!�j&$2�=N��2K��},��ڸ+vim՗2Eה��u�d�$-�e�tP�C���h�du����c�h����0S�G�;]�Q0�ct4
�2�Pi�Vxmę�B�|�YX�����9љAw�$黚�,�B��&.Ȉ2���I}�0���'�'�k\��6^��wTƎm�Jc|���=�l@�9Oc$z�`��_���]�^∂�J#%�P��C��8�w�����T��Ń}A��E�qZ�->u"����`�����in=l����s;�+jތCl��hѓ/|������hͿ�����X)*�X`���IV���9��O%����R�q�OK�zx*�,���U.ธ���l����Ť���z�'��V���29 �bUş���2?]p��� �7o�a��J\��g�F�����u1^g���@x_n���WB��U%�z�޶J� ��R�F0����+Qek�����D�~,�rЙD�d��z���Dغ���F���=���^5>���R	Bƕ �T����D��Ҿ�j�]���"�鬩��y�A��-xht���k^��үG*R�����/�7u�I-4�**/�"I�
Pf�c1&�6�=LT���	�Ն�H���3�˞�]�=����-b>�B&����2u!���-���E}K��3j3e9��tM���j�O�9iR�a����=�A߬��5ė��\ }�ͱSu{��HeVy�DT��"����;>c^�_�D��ԧ����w{�^�L�ᮗ����rz#�1x��-���a*��Ot�R�W������\���<�����3[�jn�~�q�cUs�S�����e|�}���b�p�C� UF �>�}V��g�,��L�����ڌt�b6x��_��&��g|g���hx)��@�<�"�5��ek��3���H���?���U"�x�wњ+S��k�4�Л��Ie�-���{�ᄘK�qc�d⣰��u�x�Gy��-5�<�a5"	yE4���|��H��J��>	��m�q߻R���Cĕ����5��"�ž�O��,Z�d�WQc>۟�K�Pju�m�$�Ρ�U���l��u�{֨GT���?w�+��aŔV�HNk��;�k����|��+җ���x*�Qr/ҽ�&ٖ�VeN�?�\ z�*������٭5���"ُ"D�����ųY�'��[�֥�[c<,	�8O�,�5�n�U�zg��a���z�C9'�C�m��'W���c:�/�}S�ȅ�4x 	�N��B .��$���wB>IJg���{�?C����l~�s��8,�.K=\�I0�����Y8��\� �v�j����Z�R��ģ���ځM��&n&b�`5P	I��9-����_�b����k����g���>�Z�مgu��yROXL�?BS0#�[_��?ڌ�� �<�\Jܦ�!=�b�F�r���g7�_@��n�ԛ��t�ES�A${��PKB��c�8�8NT���;ט�)�f��I�8] �s��.�Ђ��@���3�����k�����\#i��[���\��T�$�=^8��B�4��\k�"��UC�U�J� �.��!
6�Q#"f���f�ݳ��pC��8��|� �Q
��m�"�?Ddm��DځO<'Ā�G��[0nT3Lp�Ei�~cq��Gg��y�4ay�HL�\�?NH�R���^��zN�UP��zG�
�Ŝݱ|M� �}`�֨]�b.e&z�M��������4��6��c�L�\�JȪS�,xE�X�AOf0�}B�T�y�N'v�J�4�&�ڙ$�zw���H<W�ꮅ�c�D�@$T�Pz�%rH�4k&�%�|���$�½�^�p��]���ך��E�R��µ����i	��AP�� ��	�q)U�[7�c�b�VaLQj���zW
X�r��_�/���5J�kWw ���$�}>M�%��>c+�	8�a��*`�M[_�}tTi�kk��Ma��.�EwXH�q!msV��W4XVe%�
I�pt	bQ8�Q�.���N
C�"
����n��k�9[� L��}�ͺQQs�p�#}�5%)dŮt�<�"��^Ka�b]a����+연�C�%i�n�K�{�w�$��2Ng����b��|��\5U�}�O1���#3b���D�k����ǔ�,|� �Q�B"����1u�������o6�d,��ZG:L�kN>F2�j��~�D}���/Z�l���ZHGR��G��pŹ���J��4�)��V=G�ދ�'g�.NO"U�RN��̨T
A<�� ���g h���sZ��� [4��I-�mi�$�A�L�Ga���,]�~�*!��+y���=��*�T������|["�CĹ? M�F������̡�X������G�q�;� �S�8�f/��je��5%��_�ڪy��]��Ȑq헪)�����E
�.�a:M^z�����n��Ha��p.�t��P�6G�5w�51��}J�0=u���4���P�A�F�*/�я
N�>I�5'����m�}o���5dd�U��!}�3n�^�M��-���:� ^.^_`��c��#�RXU~���¾<n�A,��#�`�>�o���ސdA����e��i�M���[4ˍ��������`M�Uu;��?W��☶M�L����Ȉ�@m�o�}���5��Wl5�/��4�a�
�Q���"�=G<��-�,<X� e��|>rN���`���>`��;N��Ac�40�$�R����ª	~����/E�Ѐ*V6h��G�ñ��%{*��?�d^���K�u)&��S4b4e��
�qQ_�a���z�<���Y����� �9�T�j������ҟ�u�ʫ��RR�v��$��_5��ѡ�'�b}�	};Bj[���ѭ^ ������M м�	�cLl-[r�\�o�'��Ķ��C��B��.���.�{�P�I�����**
�&ۑ�4(@®.��<�`�W�Y�s<�$�hO�I�b���\����<o���ҋ��{�����'�	����-#��j70���U(�IH�	m��YH���[h�գ����/�2�ܣ�Igh+V\�M��&S��h2����o�^<iEI�ӥH�Pa�'GEK�fP
���`-��9ɊP&W�T���0eH�G�Ɠ���Ā+�`MA
O�u�n�8��o#���D�4���ۯ��~Cm��=v8|��m[����ީZ1�仴P`S��F(�* B��s����� �����~�ٽ\$����l��T}�gt���kbHzR� , �p��<Ϣh�d��wʄ��EY�mS����ՙ^�O������%�8��+ �{��1��	��_.U�|n/a:鷵ʛe�&�3I$�w���Xb��Ah�PQO`տ
M�9T��K��9;�Mu��c��� f�\�-�Q4F��l����(��2���WǍl�i�l���(�m��������f�K�+G*���\jЮ)� ��4"9��`���.h�dK��A�Y���HJ��&�_�����k���������yG���b?	���������i�U�o��:��ѯ�㗌����3�Q5qr�����: ɡΠ�e��*�Tq*�C����������<����.�sf~�;sb[�.���@�9�w�g����1eTȤ���,��|[zٖ0ȎO4_n{�������m�#o�2'�Ճ���y��;M©<���;��-��@}�%�CW����OZR�3�����;�E�z�A`w�j��P�I��sW�E�x���{7�7��R?<�u�8.�UHc��S��<�q�s#�#Š7�2�y�d2+_k�( �����O�\|���~�o�ni������n���-���]����bL�V�7�����v]������n�k�nl���Q ���k$<t?�|K}[�u��N���2��`��th������ً�2�Ht� �-���R��7#s��ExY#�m��zÚr�q���ޖ�^Z }���d��D�FDQ"l�|�yf�A�i���eң���0 ���勐�s�Ko�O�1�K�]�d����W���a�A��Z��;��$:����&�+��G%�1��LK��i�$dhHb�#��M�!��{札p�m�ѣ���~Pɮ42��ܸ���R`�B&�V��*�)�ȧ�(Lr$S6�n��j�D�kQt3�]���v�f��P�!�X�� �(�:��/�?T�r���Y�cS�Ȩ�8L�@�jЉ�d�7�����s4�\�#���{���fP��%�;�*��t�{��^/�7׎Ч_�ճ�]r�=+�ԋ�����ث�����<�L��n�~Y{m�Vϑ4,m:=L6G�%�~�s�Վ�v��Ӂr`MR�@w�(��d^>�ѕ�w`�����
i�����
#r��j�`�����Z�Tc�\[6���1��,�*s��eDI��7�p��ܦQ�lQ�$Ǿ�cgAc�w���4Tׁ��H"azV���>��%Qt�0_���A�؜q��.x��/X �!ycjV��rj��0&�����̪��f��\�8쿴��zɸ>@,�%�Ӽ���2��O�m98�%�����*F���m�f���-&�DQ����P�j1���Q��2�	�݄���C@ǈ�����ٷ��0�C���3E�Dg�D>A�Iо2nr�kz�k���3�]r��i�GC���ǥ�V'��k�/��U
�c7y��:kWZ�c��
]�$�̃���%fZS|��VU���r�!ƈ7��_�2I��9�����+��p�F9޸�ʜ���Jʻq]�6Q���E����Gh^s�����CG!�l�UJ�g��
�A`�8W5!m��{���g�v�x��5zi ���<��ɣ�J E"4�8'�4o ��へW)I�����~~���v��iO�+���Ua��ܮ���z��yu��.�^�U?��;f�%�, m�NƗ���@e�i���`�2*��&4�ǟv�W�)����8ͭ�'o�����U!�j���X�"�
p~m���9��T�7U�ڊa%�l"b?�GTP=W��ī�M��=@�G?k���H�y�$��^�NæT�~����y���W�B&��_�uN��<=O?� X�j$�� �Z2qP��MW~���?3KY�m������Դ� @L%�_�e�}|\g�:P ��6�t��՘C��� �K�9#4ΐ�j�`$�]��5ҨDi���Gl�Ź���*t�#Cٯժ�;�N��T���qm��v�H{����߱�I�j��;c�ot�H����@g��;;�C%���6�ש�=�1����4���>vړT��)ג3�q����-n�N�J��w?s������L�E��>�դNz͞P]���va��������Cࢥ�2h}�O]����=�h���)|�\Ѯ`c�m�D��F�ВE�T���~�K�╿�WF���(~���A�{ �ꤘ�USHR�s����8$�7dj�;�s$ߥ>ϭ��W��y��ޕ��(�:�l���g��+���hg�;l�.Àl��ǈ���NRa�F[Y8�oCT
�׍�e������A|wl��v���r����3�Qʨ�K���F�v���#�Resݯ�@�wE����ϐ�~{A��Z��,jK/a(���j�4��Dǒ*M�Z�+U���뎡Ð�ܙES��4��@����e�ɵqJ�­�Jh#��<]�H�z�o/B�ذ��;�ݡD�α�M��ʦ��8Tj'���NЂ��i�ʏ�C5'��-����c��U�=���m/�{�1�d^{��T��&�����]mW��mWc�YiLJ9
�j`�:Т7���UyR0S���7y�#�Y��9�5&n�@�~��C�����TۍH�+��c��%�d)�"؞]�U�g��LOH��4�BB�W:vI�p��,W����P-X����K��Һ��#�q��( ��m��T��ŭ��F�2����f6XDez�����Ow>����Mh���.�~�U�L�vΒ��H��� <RpUK���/Lcaρ���.���P(#΢��FJ�K����9��M+G�b����'Vfs�^iXI����!v.��ȱo�w�&쯉8�Sx�R��tM��Dz��j6QEkg/cDb�m����u���v$ɨ�=�JhЇM�����N�t�H��Tb�2��Z�� =>������j�x�"������麧�P���S<�@
Y�~��χ�2F?������;� �2p調:X���9�I�}��'�P"�N�<ɞ�虡�4�R���Kv�V�sf4i �XM#�pO9z�R5�&������ΟQGD�'�vn��tU�,2�M<N�����+�=��p�BHC�wgI�'�f�sZ�l�ۼ^�*�L�m���糺�j�G镧o+)v�C����d��Y�$�cGTv�A�k!n�9���L?�Մ��n�����Wt�[��M�$7	��_��A�)�3	J���FQ�>��Uu��O������p�W���(l7�_���$U����Hd�)��̺@Ą[̭���;��n�d+�sY_�et����]ѫ6��E��ꍅ�9���x�����|.������O���8��ܝ��������m�[fDz��=ř�I%�5l.����,:n�;$��G�r�3� �C�U�Ͻ����Z�
@�o@�:��Y.}|�ۦ�׎�o�4{��+�/OD��p�b�R�W�є���h&kH���n��h�'�_�7�S��NJ)�I�]�2c��Y�<�PSB Y���ؚt[fKB���z`���rbZL���ĕC�����kk�F��UN�I/��<c _�gx�f��./cW��f�.�6�2�?;YA�܁�����L,[f5	O�y&�+C���c�U�?�CBo9�B6���})�0�S��L��>��G�bt6�z�֐�mH���Y����cձS�I��y��y����wO��b���@hcF �e)94e�XV�����/��.�׾����>�coAZk��ÿ��s�> ��l�j��@�qq���V?�P+��=��eA�(v��rG���cz��%�"m�'��	b�^O�T���> �L�� !J1.��r3ʳj*�&aF\� ��](���㑗e�	��n�Qa����,"j�m͋�z3Vf����oF<�����ꄁx��}CrÝ����>	�k�K�z�K(L�9�T�>o�/PN<a|�"HBC�Pҋ���;r�ʿ�����G��F2��{��v��>�}&:�zp��6 ��������QOI2�V<g�s�#<�g 2���ds#1v\���7S�7r��p�p����T
0nVj���gڳ<�	ĕ�R0/�y,��X���U�����-�#�{�ӷ����U�aߛ��gx�-U0���m4�f�L��8�$���$V��I k��p����e���zv���R���N�o���O\��O��%-��p��)w9�?�r�{����Vu*u��%�64�|L�u��'�Լ&�1�8��<h��[�vC��MI�2Zt�XϷ���� ��	�do!�O���!��V���=v�d�C��)
�x�*&�)�s�|�A/Ӵ`��QB;�$a�,��
�����7>�b�K'��s�nY?ǽ��K�Ǣ�{�3���#�+��W���<���F��A��?TcݲK�4������3Y��[B�
�]��t �`!����6c�:�V�[R`
u�"��͕#'�G�S�44�T�3��x�yQ�,I:��]q���ÜU���2ð2  HCry���y�ԍi����On9�� ź �L����H���������@\��a�-�{A&�D��7�x묭&G+��i���Q/b��Z&��"���ک< #-ƥZ�{Dvx������6�a5�F>���K�͐%�H�,տ���0���]��x��pg��E��#��W}rq-R[*�T<gSu[�V�H�ˆpe���]VH�yD#�Pd�uB���Î(���K��Y{�roWL�0��c��J����A���Y�=��{��jh����Zus�3�34y���E�(!�l�
d@A�)"Q��	�ي����ũ�Nsel'[�hFle�����������;�0���ߘ܆�U�_��n�{�0�&�����^C��ᶐ�z�%_�L���v۬���gRC	���֡� �1�9$r�q�x`}OKK���t���1>���p���Q��Q�ߡ�F@o.	e+�����M����1Y��f�=�������l62t����,�P�j);e�7{�%��]	,2��+���9���=�W���|(��,@��Z�4������p�
�l
�X
OV;��7_�{\��<�B��O�Z�Сt��z��:a=늸z=H ��Y��.b?oݹ A�0��B���ݪ�,u�+b.��^��ƍ�V8v`͹���q"�)�>w�������'\�gq�
]���]��Mh�R1(�LU��`��L��pG��*�5���d<���~N��R/���-�XUb�ep�a�}J�@4�~�zk�4��bV�/�$.� �����'I;0f7��mT!���m�[#��w���K�9�|I/����ݥKt�
o�<~����`��t�xʕWz1as9}^c3#�8Q:
�A:���I�-0sYpo�n��f�cIMe�7���]8ʫN��'4A����#Jk����ӣ���~��pG�lRt�`i|��1�mY��A��	ħsV��/$.���6n������7}�����&oyr�t����:z@������94mtH�M�����,�Ċ�V��� �����
>&U�F��!�~�V)�e��0���5��Ҍ�>� w����֢nd����H-��f3���x�0��ͲQ�ZY��O&[��{.�\B絴'/���|<ߎ�h�0j�GF��A���t��8;@�A5 ����3�p��뛰
4OE}�	v!sC8��AT�H��+�xؼ�������"F�� ��^a��j�	�L^���6��$���(E\b��]b/O�p�^
�2S��/�nmfz<~K4n9�'���/���C-� /%ރ�i�Z��%�a���Zy=�^f\���x�D'��[��iӛTn� �K~�x�D�kB�P��`����D��)w�!$�yp�A����
Q�W��6�H�t�۪Z�mLKgꧏ�訸Mk(9V{�����+獳��'ҒP1@#ۥ���Ǆ�X���p����T���Y�>(,p]�k]��%�9n^��z1����J�B�V�~%M�$�E��2�Ĵ�~R���#�N<�up���[�>L�S�&U������$�ɱ�Ῐ���B�:�Ճ����,�-�֗Y���츷�ܻފ���t#�n2@z�}4���~(]�r&��� �QD���*o?���tPHp:�߽�#:���"���,م���F[w.�/C7��oZ�cT������5��p�
�=1�U���N <񲯖H%��>�8��9�2����O�矼;�i�R= �o�y.(d��|��1|$I�E�fW}"��)�J�R�ŢO�����+ᥘ�ظE���"Z����V=�N�����e{�M���]������
&�?�>��N�d|�V�8�y(��tu�X���;�F�L<��M�w�T���2 ,�m�@��w	�E��KV����������&�}���0Kw�<���f%����BT��咴�f:"cf>ߜM��s��ߞx>����~�^]锼���|���
y�E����kڳ���2��}`��=@@:)����yd@{�ݚ�c=�i�Qm��q�5U��4Y������R�4��6�	���m&��7�J��b�2|$��m{yft�XwN"��OA��0(��i���%���Po����p㉈<J4v���Sf��D��kD,���|>� _�l|.��-�����p��3���g����%0�|p�?��t�9�d(�t@��B�{#�����^�	�M�O�90��NI����Wk�H����H�v�2Uׇ\�R�L���1D��+�����Iq8���N���@HU�z��`��(�c_��-cê�W9����4� IBN7`��f!ڀ�ɣ�֥��K%9�Px\��,��J�#���	��?�9ܶ���C�S,�L(5ˏ�b��+��9Q��u��$qi//�-CL_���*̤O6�g.�$EOJO�#��.`�&>�E0����ِ�Џ"^�O�XZn����{dw�,�w����{�n/R�p�P���A����ͯ��5C *vj����$H����t�������80~M��ڧ'��Iq���t;
{�5����.[@�/�i(�:���n6��̓��l+5	�c�h�;I��a;�d�g'h�XȎ
������'���u��$Z��S�ɼ�ny稛?�b���~��hg�s��r턖�8�]��Y�"Z$�i�q�
���.��� ����1����T��&�$ܜ��Ǧ��Ŭ�*��Ġ=�J��$�%�鉞�G��C������Eb�H��+���`D�?�D��yR�������I� ��{�fi>Cҭ�ǌ1��D]'qړM�s.4��O�6��_�jq�x`���fӈ��2y8Z=w�W�n>�F�G�ҷ5dF^B/�@Y��ږE��Q�d�-���ͪ�^�՛8z�l`�f�f��u��
����-���T��
�8�khl��PW����$�n#�+5��:i�^����ǡ���_O]�=��d�A8i�e��5��-D^n"�3�6h�݆3H3eͅ���{�'!:UY�x�V$K�i>�̉�_>�������[��Z<�E����:�ȳ�H/;��T.y��W��k?��ФǦ�}�YI�lŉ��K�w�FE#N��爐���qm�5���J����KP��2j/������=�__<��� Hf�1��@�{ᣏTŞ'��@h�d
�!u�a�:̺�tL,�� ii��?���q?Ҁ����PE�A�Ďn�̪m�@P�]DC��A;�� ����#�P^-ty� ;���A�c]���Y�`,���g���V�+H4��=�;-����,�֍�����#�[��j�>�}{��� ����{����Q��
p�EJ�����!Mdm
%���z^K�s��jb�y��s��z�S`��\�8��8���AW�Rx�;���N�H]\͚���~!��jP�Yu���Բr����5�Ox-n����0>��FI��)���}�k�xr�[�l1js����3�E����щ��N}�b�c�N���N��oK&u���.	�=���!��=�.�.)��R/<kt�Ǚ��d��.�4�A,��!�JT�I�j?��c[ʨR�a�������~��)�-�M��i�FGK��c���,怎��يk8�f��d���]Zo@H�!�@�+�_ǣҩ����+��zoy7���1�'{m}fJ��5_�明]~��|G9�z��z�����D�n�),�o<Q���=����)<l��Fz��uh���Cr�Y�'*C�¹G3H?$y,d��X����8ƹ!Ȉ�P�ҪTh��J�ĪQ�����XQ8�Ez�c:w���=�UF!C�]��t^G ]�V���w��y3�Bb���XC0"c��lk�T�]�
$��cD���ǛS�,e�O�ϒKՋp���oQ��[���Ѱ\��;1��J%~��4�J�or�]�Z[�|�gqf�v���R�5�e����Y:�Bix2�Zp}om������K�r�1`��V������?�ߒ���+�.�WO.V���D�Ym �0Q{�*��ԿQ�%�78������N����  �^g�ߓ�rD � ���ّo�~Vk����l&B0Ъ�{v��JZ̃:@�c	\��N'2XBAy��+�H�!���bC1k���hF��&
�7�O^�=w�j�I���������U���4�a~�<�U��]p��3�B�FCζ<F��}�f�PԹ�Z"I>��!��9E�z���^8٨�ȯ����Ԉ�go=J�X:����uG!)�i���.��.Hyf-Y~��G�gJUz'*����QѼc̺ �̜߯C&��ݷ?M�I�� �{'�4��ߺ�ۡX��k@�#���]����Ө�f�
�(��bA�jݖ�K��h?��Wh�q������ Vᭉ�� k"�9�a�� ]3���Mz��!(
K�}�>C�F,�I��`<,�n�Z¦�e��l�y�
Ci5��ݓ�eg�ό7 �m�V�(U���d����9{�2%K�{�M<,ޕk��E;�jPhz����3F2"�fj6C������x�z��g�jF�O�:1x���_f"�D͆��o��Y�n��m��́��+���i	�:e
Щ+]������ٮ��fԁƝ��$����pv�$��m� �[]H��g$1����jt`)C%��Q�}�í��֨�O�$j����v��t#��lU�d��,��AD�#������Q$CN���K��\j��|�����˻'��JA
��."!ԑ�L�U�P;��r缔Aˏ�.��L4�-�9N��U���F���`���~d8�o��1K����&�eЋSf��v5պ?Ľ�Cj�	u(�?*�����Ho�4 �d��Q�2���g�x���8:}d�Na���^��3c�q	�<zHg�>�Q8�ygi�g �"�i�¨9Ij�	��4���5��ç�0� O\V����~9��e���Ħ�0]Z��R�1�D�)��ų;���>#f��n/�=/�]�f;���O��ߒO�+��W+}����!L�2�v���ٜ[��� �Q���@�wi�L@Y�#ۗ1���|��=N.U��d4�4HM��^o\��ɫ8>��GW�|xSeNyx)����A�]��	�mQOHR���@D$��
aI�j{��6"�iҙ�퓦<���I��(���f\��>�27�7�a�o}�jH��Ư/����j)Gsr̯��<<��I��M�~�]�d��,;��/d�\��qj�5�+���>�
?A��Ր/[[��X�8��i) \F�HڐK4�n���6���]��}�)?G�g�l2*W�FA8J[/�?E����UtR�N\�7�F��q%��������Ţ����;7}{_E���f�2[���>!�pYM��1�MYd����Nk�N����`�4�'e!�t
�)&�
K���*�p8m��#������sn��Q���������:?b�B�h��.g���� �G"u4{rK@Y]N��{'�g���̱k�=������r����c3ҕr��p� �*����i�쏸�����G=pDIZ�,�o�Z�yN�L��B�� z�/��0�eZ�)�1���L�����k_!�%�V`#I~3�Q�=�Sn��� �](��9_49ʤ���t�xߋ�b�E]�se�R�j�24Q��y~��{P\�*��8�CC�3�;W�_����;F"�7�/8�~����Yo/�4ř�'�-�X.�0?��f$�K���Ʋ�����=ֱ��d�bo�/�'�w4�LM���9�^a��v���+-F��`p[�m��ѫz�u����s��[�$�8�Z���p���Mc6��5�T���2�p%F��H����r�`��	��!+�+�#��U�.�~�AW�
��&���+QUz�L�
��׺��JV�b�}R�J!d.Nu����L*�uJ1���:O;����q�f8:f�+v��5u����8�և�0 ]�%qp _������C�X5�q����i�<���'� �dv����.W-}!��'��٪<&_E�u3s[+'��G���Ʀ]�S$��G��f*�B2��3��Z�%����&`�/�����u�U"��};��Dr(U�cUtY0_�ԋ-i_�-�ņ4ӂ�1������m$�D=���{ߴ��'��_(\ٜ=mG��S�قrG��b/q~�I��<I)"������!Nq��~�D�(������^��#F.4:���\���k�X&{_����J��"v�xL��n��qv镠�@�sS��Dt3��Y��.�Bb�xs,�.�V�R#��&�9Z�'�yr��� ˼t���H?� ��"������ B۶�'}��e��I9�AS��BIc
5~N��6�fG�X;p�Q�W���1�N6]ą�\i��\u�$�u�!^mvI��=��o�l��S	Rk��{�%��~Q�������[(E냿��2j���Sk}1�ܗ�N�� ��QI�����
+��~e��*c��J����FHs@����M��)��,�G�5�k"��tr#�&g{�s	i{��uLX'c�F���,�.����x5Ԅ��޺�o-$��ՇM�~۩a�r!֡�,�e#�H<}l��-�O)�f��^�@�b_�/B�`t���8�A*�	�����n
6|���Ք�xO�l�����W�	���3��X?������.;��x;�E�8:"@��̊vp_�c��*��e	7���{{��jm���.��O���[�N��G֖�u���n�?��P�?*d��y��|Co�pw�T�h�O��I�X���C8���\)��E	�<IJ��Am�t6��iB�W�>A-N�����ь�i"��Z��wE9�F&��	p�=�'�%�̆�@�=�dX(��*�GP�p�?�' ����4>*�~��fY7�`׾�/�Sy�`8\���
�1MwŃ����uS��*�"���b@��b@ԋ��,��@^☟�����"����<J@3��b,	��y6'j��0��th�P������:�p�U�$@w�����ǭr��N�W2x�"�>3gU�ki*�j��6��$hoމeL��y#Doo�<��Y��o�n�ÀC}�1'P�kX���e����O�"l�4Pe�m\xd�U�_�Y�.K��@Ȅ�^�{AT�C�Ȧ�a^.��cjo43���"+��I���:�6J�Rz��o7�iKL8�B)�����3����*zS�~��Ч����n��4�;��LI6���";�Į�_3dk��X��j��j&^�4Χ��������b��\5�����>�"�G�[b�����a��I{�d�}��Y���Lq.�Y�'@���Ͷ�5,,!`�3L3|A��y��]��1(x�t|�s��Yw�چ�\�`�M;4��υ�㨇[m��ވl�ErLB9. �{?�jwY��F"}�N�>G�� X�ɥ��\��Z���,����*�G��e��22k�����qN��%����r/��1d,�5����/��BR:�!�:l0:�{���t5.)��0j��˧C@08����\�׆����_��a�"�
l�e2��)�r�ݻ�ٙ��*���5�z����q������g@,QFϣ����L�K���4/d����8��p���L
�dvrN�~(� �
*�(��d�@7�zr�0�M5�f��>P>��"��)�����ѽ��Ylx>�?�w!V���K)Z�/�S**�1xE�/c���`}����h:��_`<<U+�! G �Ȫ"�ۡ��H�������l��V6�J}��,%�v"���;Eh�Ac�:�d A�j"w�j
IZXVa�,��45}�π]ţ����7½~K��ԑ����t�$b"����� ��Y��qt3�5U�5����rG3��}NO�Dtm؋��ˢ�gԅml���/˟��ɋ	�7�Q�U��ID�������/v�_��Wv��Ǹ��T}�QË����ؒv��&ِ�ΒB��C�d�<��%Tfa���(��3��(t2�Q;����c�#��w�����)'��gg�
�/����V�oǀ۶��?ܖ�J��Y�U�0�'��Ca��*g#�5�؞�ne)�4�g�R��l����g�4d�h�C�����	bXӥ�'/b�`5�,�4�9���ˌ2���ۋ(���u�\e��D�V$7��l����ޫ�(h:����*�z<c�T�]�/�+o%��JN�>t�1�^hb4A�/B��g}��e���}��u�ߚ�ԗL9�E��&���p���[�� �c�_N�p]�/��^�q#�+�ﺗ�!*�H�mxb�-x�l�U�~������vIhK`��?Ӈ�b���w�-�"O2��?,(M�a�D�/TWڀ0��V|��qW�RW��TO��71�,�4�5Fb��)�ޑ{A�9���#��HeO� #a��^����)�!!徶N�*���X^����qgk��EY��@�7?�	Ln[�ԫ2b��e�y><0�K��b�3'�k6���YE����怣�b��|�N7��;��%5�ľHң������rCsU�SO�+r/@/�K������O�=�/���������ɪ�k�U�_��/��!�	���b��H����(<��I����(í��|����eV��:T��'%-9��A��p��+W�׋2�پ�`B�� G�-����0K�)fǻR �:�D�e���/�ifV�۫��9K鉍���Ga���'�<o�}H��D�:�p�-(��������,�2UG���NKƼEq����ղՔTI��t$=�zWB�m���|�܃hr�^ ��Y�)6�HИ0�4�4��su�/�ZQ��b-�� UMO��&��ؓ��\(��D�����>��x�g؋�:[��6j���C~>�y�G/���Q�c��,i��i͵��wwƶk��p�����Y]�q	���m���&[�����PS�D�Ԕ�D�@�?2׉
w!��$ nxM�'�_Kj��B0@�	G�f�t�ק���{�ٓ)K��$>�#\$Dy����K���~�����ޒ���@����Vټ�����@=X�M%��1��A5^�ׄ��{�C�e�}}�B<��Åhݖ2�D�f�]�κ�§��;�`7 R)���DR<��Fr`�[���8;$��$�p��T¿��Ǭ�ߟ�,���6Yψ�D�����HQ����Ȏ����?�Xp* h7��l'w0��� ��OB}=�_|��9ss��}�|/�\��9��xN��fD�|I�k�Ew��ƒ��>wb���0J��/���݆�'���������&�kC\i������2i)Ъ� �K}	��PvOz��؞�Oƈ:�^]2�ob`�t@���M@%��=0nk}���K雭<^˾î?+�d	��A�JH�d���h��0�6H������������D	o������ǉT"̦w?�'y�8sľ����Ej���;f3(=���x��}�'�zRt��d����˜L!m;�)Y��j��J�,bᤤ<�/T_�gG"Hׯ������z�)FM��U��7�F*p��$���@P��ld!�F�!G���
�P����!?�85�9�-��R���=���N^Fq Y�-���S R�)m�����+qG��6as�1�},�oj�i�1����k�e�\���M�� �o�S�����-�%�q$V��2ؔ)����_�nʹ��I���5T�l���L��iC�Η�ݘv��b=�<0�+��ս���r���c�)�5��ы}g��z��R�%Pg��u8��>���j0!D�á2����~�@X��̍1F���(C�2 (d�C�S��,R�������ƜS@���.�d��J�7�C1���i�͛����A̿�>bm��pw�抅J�PV6�6�Yqx%��_W2�҉2̃q���2#â�th��y�����?�vR��'��(M@�����6T[�D$\�O��6Uv�x��YK
��Q���a0�� �E�6��I��a3��f�2���w�k�;r[&<fo�m�q�3�Հ/�$`!q�{��̇^
�I}@n[�\��V�c��+��J8����C>_ �J�Ǌ��l_Q:�w�?�⋴�6��3��~p؜T����m�N�;�U�t@(�%���h�8��A�֍��I٘��٨@300=��;��\&��>������Z?b4� �9r9Z+4g�})Zu�&�q��W�e4.�1[���z��-�(M'i�?��X�%o��^�����	Z}{~+����Cz�&�G�Cm�bu�tǯ
<B��"�G lC1Y�W�_���5�\)kuMw���5o��̘����s�/��f{f-�i���ϴ�[Qy�"&�t�i��ׄӐ�%�Ů�A�9T�!/n�,�;�[T���ř�����,L5�> �lc('�J�6'�H��Z�S��
�E>���P�G��#I�����ch��	��ғ~9��<�|���A%�}�&��D���s܇�qQ��%�g�?�'�؝����X7��DSGg�Zi��}�bK*K��Q;`�%��[*�ё��uo����O�~M�M��E&��{l�u%m
W����@u���r��K�)�^�0(����G�:_h����)��9��O>#�S�7(�`��FL�����wM��C2%9����ʩ�E����Ŏ6�M�1�}���"���o�S��jDj�>����RSSk�F��2a��}�TV�ʌJ���D^@A������Ѿ�EÜ��:�PUG0�Č;c���d]uE͌�g��5��!n!_	v�� s���	 `�/jRv��F�N �U� ���]��nv���/g�PkR�>��&�Q:��}��\�P����w���
��L�o8�s~��v�Y�Sb��W��:�?����k���:Ƙtv���4!��g�G�Mɚ{8}񾛢�9��L*ɡX�k�������|lE�b=0w�8�)͛_��W�j��x�C��p����G��N���,q{��3��;6Z�|n���]Y������.ޕc�3X{�7��b�J����Eu�h���v�Jx����sxr+ ��q\��s�����`o�܆M��-$�ȯL��/mo\M���/4�/���e�4�:aNg;�-�~�:��"�m2�i����y�^/4lK�6~	�*�L.33�>�d��%,�c���Չ+i�ix�1�Q�
(:�� !\0�K�e	���y$`8��f�zV���b{k�;3t��{�{�
�^�mz6�lPV��� 8��g���񙴜�#q7��i�l�
L��l�@�U�1Q.��∿6߉��,W��?�@a�� ۷�q�q�[;�QZ�x���oꗔ ����hpYg�*(|b�u��}�Kܛk� 6���q���NqN��ʑ�X�'0��y���r��@w'��;:���gp�Ð��=NR��rͨ�f�j@� y*����icyN薜g�*Sg�Ì��Y�g��@�3<'�o �jf��=$
Q���~�>NC� H�Gs.�s�:S��Eut�	��5w�u��V�I�ځ>[��UV�F�>��x!�dXO����"Dk"��]���j��_�����8���+���D��c�������w��}Da���"3F���P�,�����{ϯ�Ww?*O��p��w�مmu���r�Hء+Vy��N��jʉ�D�'�}���ֈ�ǴS5�� .g�Iw������A�щ�Dǎ�aOKV	�͉F�?bNd��q�7z!~7���ZCJZ�;;lņ��&�θ��BSv�ω̹/�bA ���gEaw�mĮ�A%P$z~\1��I	z�1��>���p�*B��y���X�h�7�/ri�/�/!�6��	T��4�#6'ker:��ia�gsB��WZ�H��I:�ؖ�F1�_��������[n���y��+F��?h��q��w�M��ADTi+��b�+Uv5��{s�Y6r�)���9/2D7�^��3�|�����V���S~�:u�b::��%/�r����3(��^��a`ov/<��C����wK�a`V�<���ޅ�r�\J�m �Ѽ���<)dz���<w�	���9�N�G*y��<9h;0e�vSb���/x����(���H��d ���>�3�W���NQ5��VEz��� �K��ۛ��i�ȿ��5L�i8D1���Ú4m�
3
q�C��
�C�,E6��T��C�W_v��y��"2wN�+K�Ư�1�Å��v`m31�7�\�>2r���s��{�n�wۇA2��(o�`��V��?�/�X��)hv�C1����/ ��|ƻ�c8�ء���gU�m�R����M����i��FZv%��"��2����ܜC�ڶ�k���x�8G����*މdII]����h��W��A% Հ��!�M�����a�I�����\�{?����<M�$������&�?��J�;�vP7NT���n�i��Z��E.�o��q(�ug[�!(���Ci�fP&��1��IGM�0�G�k��9ZL�~G'P���(�{�0$���g�!Ks����<���2 �§~�K^ڔl(Pr:?=���
,�6�V��t�L�h����hԻ�܊�Y�<a�����b�U �ϝ���i:��Y�����-��6���ż�e���/5���u��8
w��I����BTM�`zh#�P�~c�v*r�-5_e�d��Mqi�boXU�/"��kg#���U	4�I���PA���0`�sZv�ÖCeP*c�?��m9�E�AT�cC�L+�
5v�ڊ��2��1%��.�lT��Vn"v,�8Y���"ԡ�"��T�j�S�R��9�b�>�MLM"�`~$��˿=���t����]@�j�}XtV4���%\y�
���S$�\X��J'm���Y��y�7;�C_a��S�hc��_�dr{��>H�ţ˱�:�5D�%����՘D���"f��U&��͛FӞ>çť��m�Ұ�c=�)�ڥHE�߇ިk�t� S�y}�@�L��pc3/����g�^��l^�ψ�/;Ws}~��`��U� ����ɚ���	��"'�Z���o�� L��,�u|�ŧ��F|��kn��#�n����.��V�zŒ�DGo~������Ƿ��O�<��Hgk�B��n���rwcb��& �!K���v�����Z������I�V/����J٬����4iҞB<7!VV��@�7Q���C��Ї��[�'F��w��NDe/��..�;�d_U�5Q��WV��k ?>�x�B� "m�gL](�!���)lg6C�����J!q�4�����euڜS0�X7nr!��
Z�/E��ө��ɭ�Q!:"���e�0Ɇ�_����.ǫ+�����Urj��e6IBGqo�2�;�� P��7��^V�HY���.c��U�f�nv�u��B�l����8�AXZQjN/�$c(!�ً&��"���G��(i���m3���w��U���P�ؤ��u����h�K�*b*�+��ܒ&����˯����/L=Wd�M��;��b���b&�,0��Fq�a��-�ԙ��L��z�C1�o�3�xIQ*,Q�RUv�O��MG�H���A�˘��)�G����S/���>�V"Ɋ��������`�����b���]��]u��r��B�l_��5�t�d�}��8~޿�T���C�!7��U������1��`����'3ɵ��~e�t`LAn-ݣ2�d�e\n!��J��5F�
,��`�ׁ��{Eat!�<ب�y0y<��1�2,8��J�z"�8�p>��]�S�U��5� �����d�<(�o�=[����2|�b��:��w���)J�>;'A��߬=
)�����hr��u���+��/�k(o���-��j�7����	�YNn+i�&�S.U�ɺ{T�vњ�8w����������yXS����4�6û�0��{-pc��3z�u�E�e��߯.1����ZJ�K�:�����uDyH���$)	:ufi0�Y㧻n`^�Z�[H�J{>�w���{���6��E|=J���Ů�B�Hln�R3��PP�����+^�ZXn�T��w�s>-�2"��]� ����	<|�����9�R1�+�st������3�uGV�y�ح�N1U�����ӎ	�d�U�`?! ��� �Ք�\.�2���s-��wj�y`�߀��
�6�x��D�X�l:��Exɒ�8I/|��w��M�:� k�Z�t���@��=sV��}��E��T�����&ځ�+��5m~�̼-��D���Ê�Ova�ȹ�B,�5r��C��IE�y&���<�l���,�~��Pf�>;-a����"��!��I����/�D�"�k�Lj�2��5�d����7�*�&�n�9��eX�g~B䄕�������V/F��ujg=�����A��H������暍<�5:��v�i�O��-'.Y��N�W�#����TJ{��wzWb
ot96�������͈��ь��&$�)�6�h�W��R���
�a���6V�೛^~��Ȱ )D�����7_�	N��G�xF�x�g�1�D�a-�C-D=]�:���_�$��JэB1�#�ȇ�����	�1Z�R��`�حnt��x�`�4'���+�ރ�k@�n���Zܕ���sۚ������4i�oz������7�~
5��~�=������q�Q���SO�,��3'9Ѭb�5.G���G�m�\SΣɝg���t� �uM8�%
^���u>sn��[8���r_��=�	+
�#Հ��'�Cp�@+�C̛T��� ;͟AlY� !����!'?�&c���~���D�\��g�T��������IԄ�i�Q�8<���n��8���$��3�09�;W�2q��k��}�f6q0GS���*"��tgQ��]��	/��r���~�o@l��T'CMWn�˰Q鬵�٦�ԙM��IX��͠��B��?��[��dv�c����#�]�9�<�قO��t"$9G��uH��RI����wS?��l���E+����˶����<��H[q�y�ͦ���X���>~��0m���[��D�#����T��,DcZAk��Ym}��C�8禿_�U\��
��҉{��$@�dm��ƶc�F��ϐ�)���?��=��QNl5y�+u�x��]��ݹ[Ғ��.fC���V�z�?�}MkK���0��-���2���ah�Փ������]W(��&`զ�ۙ��
�Rsw��a�N"-�R(1��O��(�C"�U؀�������4���]���Y��_��t�r�4b���٤�ai��	�5�K�`sxF�DwG	���k�}�-���.�ǥ�咀m�
e"ڇ�D�K�S0�DP���:�� 9���)zy\�2H-��� ܅I�#"@��
0���Ja���l�u�#A���k1�?�m?̜�*{$]�ѳ^�Z>������h�w{�U���`��p�.�+�LǦ�	�b�AK�����+t�e�6穽�'��c�6aQw�j�2ӯ[�F��1 *FU�I�Ѭ���ّ�V}R���ta��RD����p+H/ö���p��uz�q�����7[�K�UGic�X�D�\;��B�K�y
�����p	q3},�t�,��(Ey�FS�����i�W���踳��.�'3�8΢��"C���X�H���R�`��8,�Rd>HW	�]�@��N��r�!%M���@�o�B��v���o �rtv~{��?;��k,(�9Lw��3���{>��i��(�{�~4_D��~�>7N��}��K)�t�:� �Crz�}W��9B���B=���&�'}�R=���,{a��Dc�H�����5@�j1�&��7 ���|`��@#�n({�L���nBj�g L�xew)��+�xCڲNG$�Qn؉��2!����p�ßK�`$�Kp��OY��;��?��]�<,���UMM���zk���~�J�U�VI��1-�˻��@��%�*J��m<��6��j��P4zy�' �	xJj� �h-C�ɕ��Ur&3�o��&L��ą@��[�5F�e�a����&���E�)��y �J�3��u�H��A�W�ׯ4�F�Y�w��	0K'����˭��u�$o��zy�s�#�S؇��$���բ8K�"�	�Ve����;��UL����q�� )3u|�Z��UY�Z�����]?������`*��P�z`�d��#�2���}�8[��ӋH@�~�7�F���I��2�;V"����Y����7�C�d��2�sj��?�v)�����s��2�Í`���+<M_Bփ�-�P.������~-�\t��3Ҡu��Xqnz���1����ře%���nz��ly�h�8�����SorJh��Q��M��G��N�4,��K��%�Mt��컄�D�v^mw�!|�O8G���mO�ON!�	���ۅ\����򛆉��9�xD�����m���IU{Z�SC�.���Ic�.T���q�vE�V�` ���6 �]�f��	k_!2�HMÝ�/U�r���(W�q��v�4��]�g9}i��v������6��h�eA���ko��0n�Х���%� ��.j-7�$@#?�43.v�b��ӬS���J{+��C���߼
5��jw-���l59�-��`�kϺN�L�E��hb���g@]wE)?��W�
e��n٦�;VP�RV?9���W�����9�߫���ą���"S�����7_1��Mz�6;�2]~:�Op��y��J*��CX�w�ި�ezT�]t�$U�iN�;[��a9�����?�W*�����q�x��l�A���>��]�t*��@G忻1�i����� �AX�Md0+�$�W��A�"\�{�,^�Z�t��#��hy��нK~�����Y�wO��ܡ��
:p�,�q3jW���7j�!pv���N�O��r8��Qr��p��<�z��?��cXM��-��Ѓų����k�bt��t{1k}�OZ����R	��� �N�F+q��(O��cy�wU1T�Xk��Ƶ	�æ⃶��$ O7�L�D����
�o��N���E�0�Q�-�4��*���ЇqG�U��A���2J�=Ļ���&wZH��f��A`�Et�� G���{p�b��Pl�����1qg<��@�^n�}Sp�s�Qg��S��&��7u>�9��Y���Q��/=ic�������x��}A�9�r6�?�����,|v
�bG�F�R�O��`.I�r�V���a�A��7e!w��"夻��z�����f����\Q!i�h(��k᰸�Z��#�I�պ�~�i�l�b�F�%0��Xǳ ��h����빗���L����1]l"ҙH��o"���FX�9�.�m�R\��_Jށ�b^0G ��	6���9�}G���c /t��V���੨���p�gʡ3
�3����� �����=�g�4@�!>��N��3t�/�;P� ���x!���z����N}�1�P��"ٿL(�`tD���{o��Vj�*�����%}1=�>E"����T��%^��Y�.���;���'_���X�M����I��s�ؤ�BAq�T�+|ª�h� ,P�+׭���8�d�����\oBo�����ΐ�]w�P��� ܡ�
+-]��f�,ӐV�Z��H���,�G�5h;��CqW���N�J�]� ��0�V��I��9jOiJ�,w����'�/����=K�8F�QO0ڨ�C�KqX�ŊR���1�hs�-k�R�����Նq�18F��e+F���4㪨>�����uF�oF�+�w��_WW1���`�`���B��F�izZ��k������ѯH�9@�ڭ�����|�\���W�B!-C�iw��\ƝQ����Ë|2�A�qѕ]ϒ��k�I>�>M��^�s�-���J+��(�g�\J�������
4b���ä�|�0�l�����f韭wI��~8P��x�Y��� ^��e�?�b:�N���g���x1��p����iI-s�3���ω������C6�=�bϻF�'��{��}v	h������0����B!�9�ʈҵ�����y�	�2�ڷ�I��"��3�8��@G2�����Pj�������V	]��F#�*CT�}�nd�eģ�צ�tYB�=�����Ms��Y�m��@qa�y���j�V�i���05�����3�!�5�l��*��~�����i"a	�J����p�X�i���rC,�i�����w���`{m=��u�� �y_'���ENE��Z�NAm����Śt�k~�`��v?K�ZY�Ks7�(�O�&rF|�f����A� �T8ej��F<�VHOp|S������KŔ�e�4���̺��fh�΋IOR3[b`����\NQ�Sz�xY��u�{���?�}4�6=���j!��Ӊ�0�<*�c��"4 ��%�~˚M+�������0vF�� ���ڡe�ڔ<�;�e������tZ͌eL5��2��]-���>�������|��l�7�,���8����}��%6g���`Ќ"m�j�ۂӐ&�����)qf4��0#[��ǧ<��:�5�D&���k`K���SPjl�-?f�,���qR���Y����PY��&� ��?��֦U-��IsoZ&!?�q�-e���{>���t뗉��K~U$v�i0��&�'%��&_{�u�c�㈞�����?J]�9�KD1�9�o)���KF� �t��uv����V%�t��;�^t]��+L%	sr�<����i*?e�4�:/L���R�����X�r?�ww#� �"~�F�+7\74�Iؿ mo�L���v���1�"_z-7F�4+��hd�Y��M���r?p/�a��1������t(���b���v��P,�����] ��\kJ����[FK�ڶ�b���X�N�E mR���&b��*y����d�����n"��X��G� �h��\��7~��\6��Q~}6����{)��h0�ஸ(�|+aJ�@&���r _ȶ�qپ/��ʖi6a4���e ���>�^K�k�B��#�R$:�����������Q��)a��s��-�4!8�@�;��)��Vdy�őԫ�
2,�#���qlq(^q(�吝���DA�"5E�2C�
�"�R�־DTH���cԩR��b�r��Q�:C
v�x�K2sA�Wg��Bp���� 1���>ys�+��~�W]%���g l+p`�A���l��\���)Sʹ�(T��������� �b�F�B�[�ε�+hSkw~�N�%\���ؾP���D��Q8���*�teކQm���`�wp�_�(�_� B�F Y>n�+Sbz�s�N��d54(�nĘ}?x�#&���I���±S�s0���`켬�Jk�+	P�Jz���c�4�[m�c�i�rK��ʝ.�^b/��R�@���І�ci���&f�.Ʃ;ˍ�d>9@B`����|�m{��-a?x�:�wVi�$�[�D�������<�?؉����W�o����������Zn�s�@u\�ƴ jhX!`���`�Z��պ���2K3[���Z�bC:�4K��>�a��L�F�=:��ʮ�qJ��V*}�nXU*�6E�ͤ�0|UY�ם<H���[[+/�k恴e���,J\�����6�6�`�>p�I��Uhr�\8�;tnΧKN.Q���թz,z��K��&h8JU�e{�{Y�qX^z�H4U�}N*�k�Re�)�I�	�=�I�w�T�*y�t���҉DQc��$����3����5jr��w.�C�g4��ȋ~��*f�_��ٚ[ԳN����Z�G�0�����[+n���y�T3ǣ-��ko�GcAIx����&�3(�F9u�r/W������I�s���$Y�7Mɧ��;�h_m�#�6��5�*۸�րק�q�l}#��[�N�#���i�'�k���r�s�ܗ?��IT�5B	��3�v^�z�ª��y��T����l�w}��R��Ńs�����ի�Y���,�L�(��&ri%B.�O����fy��k��"$-��^'�qGU��2���9�֩�|�y�j�����Z�S:�t ��l�?9���z�;V��U� �y���2n�P[���R=�^�\Ҍ���d��E�3��/�����`���z���l}$���Q��LO��Ԇ�aiY;��ݽԮ�Y��FI8߫m*Tx� 7��?����r%8��W)��Ǝ��Z��|0^��̱��})!�f��.��Q�`M'Wj��@*�l�-䮁���?��i��+��Ő��1�θ���$r2����6�-�혩��Ş��9��%�ВBŐ�Wxv��&k^T�3#@J�yءE��!l1���me<^.�_�ы��Ы��)��g��b�����4Uo��n��z����)��	�r)w���_A�p`w5a�h�MS�]O���|w� ]�-�՟8�T�Y2�i�����Xc�_<�*�����-�W�����r�5&�$4@'b$��\;%�_�?;>�������k�_��?�kڈ�+U3�3��k0]�+d���AV�:��jq&6�#�r=:�do�a�%�-ٮ���Q��4v���٠� xwm8I4:rϲ�ӱ~�%F�0^j��&�W`�+:SNpɹ&a:#î��Уk�û�L���;�J����+��'-�Ţ��M*�H�z���>���7��/њ�
sn�5�	����zB��}.�x%~��~^��昒�(Wc���J��ݲA=�����c�S#��U�3�fN�����������#ԧ����(�8���[�EW���r���L8<���l ������e����xB\c6p��i����vyP���o��X҂E���/	���!�VQ�;�m��q��~�\14��By�X^��|!�dw��̂�\K8�L��o^�WD�f�
~������j֙�f�P.����n��i<�� ��'���iJKF{��� ۹ ��*��͟DY�6�4!]tVk������]�']{"�X&��,,-=JcK��Y���7�a��{&3���y՘��;y8A�J��@��x�^���Qr��=f��������O4����@���<%N�>̚�_s�f~D���.���'q[��ʛUP�9{g	j�o��f_�\�ܛ��l�i��
�N��z��/��+�ћ�%C�̄�o���?�"�~3�@l�o�XE�-5��&V�I�&��!焵������%(Fk+5�ȯ8�:3�KG�,*Y�*K�{�f�.ʢj'���N��@l�d�py(�D੪�aPNA���)�s�9+R��:�/	���7��I�?ڽ��a6^�Fb�i�wf/�:�&~��:{������jߔc���;˒�W�'����v��Jt�Wǚ���!����,�W\��.̕��A%�`:,����zOT$R>3�T�c-�	Y�SO��V�����u g�J0�p�=���2��G����B�`z�����[���4��B��z
;� ���h��8�>n�?!U�)��������{��s����ϛ�z#�����Nm��VW��e�LP�B���>��&ƌ�+�B�"��aIs�E�� #0xw?vnKm��p�������Iq ��O_�u����l6{x�AU�
=����˘�d�[UX$�1�ڬ����e:����|�2"T�����(�n*�L<m�1׶tj�pa�J�#�.VsP�r_�W8E���I�TzPx��%���,q��Z�޺��AL������oâO~�Jyn��8ˇe�'ձIl|*����3���h`���k|81m"���9qP����^{����f�|s��I��v��rD�z�S���,���΋���c�5H��4���L�P{x�kIW�%����K�י?�p�W�rIx!����p�6K�>�ZK�F������^���R�Y�)4�^>���9����a�rԇ��W���.��FDs�
��{+P9�hy����{ܕ�y���[�_!���м�)Q��^����kz'�k�I�&�+e����ž�(�� ƥ�Es�AR�g��Ԓ��x�F��dM�C\�-d<�n�7!�Ι�pjpE|� [�z\L��Z�t�Ti%��54�A���_Z�ً�� ��7��/u��q�j�z;��O�<���.�re�T�g��F�.N�Y�r��ȧp�ӱ|9S/#��w�\������ip̨�wl=��G�Yz4���ȫ�V73_Kŏ���g6�X�[�Zv�?b���VfܮxI�߫%Y��it=U����r�l�}���5Jpކ��|�� K r�W����F���ð�Ÿ����_�75�| ��r�H歨깭���H��V|�� ��s��}�#�+���6��՜w���"�E�/xH!�)�>�����#Heg�
�&�U	b��;a�)˗_��IT�����N�E�L�&e#\=_^~Z*^�х�˒��O�R��]
Z*d���c�)eP����E��_���-�垯�HГH����x�C���ij��褄?m�\��69�	hH��R	B��nl=w�vQ�=�C��������㚡�c�NvZ9ݗ�W&�����+yY;�xiA�q�����d�C�6��~a7�i9�y��A0����m|b�_߿e��+�)��F���t���2H�ۃ�ifPX�)7΅B
5 �#���� ���G+��{J�24����'�@ۀTr��a�L�;�a9�<	Y��|��
ٽ����ҼP:-�W\Hr�Z��9��fs*��P��Xq�.��D�c��yx�H�!�[I��ꯅ����SDL��pf���H �͉�_<��0	��F��Y�7�뇱���ݿ�$�]�zG��ϼv�3��_�u�W^���f���~�3)�~�6S l�g؁����<�y���Q^S�nRh�f����9�]���&��Q��q�w��v��/+�?뜒����ʣV{�垪�V�'��%���¼�Z�܋����������hZ�����C�g;���l��}~gi�Vqc5H!������j�'��b����P���Z���zg}�A���#V���R�>�Td�E��Uߜ֥��\����4�T��b�q�
_Q��FX�ܛ�����ʌ�O�N������\�8��'�_�.�H�m�|�8i^�ۣ�B8�3���g��կ+�:��P����P#"�/a���E�l����齧E�+a��2O8f�)CB���Xll��IlJN��Z�'!{&��a��rg�Y�+�l}��-Z3�4�%���^�v�^���{��̱6��x*�],o�xH,p���h�/-�D��	�#�M��Ѕ��s����D�Hm$�+��J�Ph�1��h,�5�<���ă4V[xG��`�7Tk�ԓz�������,a�
ze�2�\	�G�Li�����2r�[EL��7�B��3d��m<��9��Hp"��עyD\��r���ş�K����=ԇus��nDa-�l��G��Ƕ�_d|C�Ɵ]U}R_�ɄA/�IV9����NSo���M�)�)��焭v�C�6R�vO�u�@�IT�bW����2��8�V:h��i'��0���.xn�\'���сRbw��M����hEB�ݬ��-�ޢ߈0�4��4��)��G��~���k�����)�6�?�A��Lo����8m��Fj����#IR�1d���⾫� �(��(I���%�;�Y4�RY�`���(��ۤ��@��q�<�M@��zn�F������`G��� l���\���ko�z�~Xy��q�.��2
 [��L4A����y�A�?�C���9�ex�|�����ϋ�z�}j�ͻ��7���2�G�[��B���:� �98W�#��}�)�uA���s����0�v��o�Z�<:�|ɧ 9�P��t��w3H_\l�]�G<$ҧo^�(n�IJ3�2��BTa�kܵh�Kl���NN�8σ^R���~�:w�s�p�Y8���D��w冮�9�aۢ��t�0��ū�kY�E�s"��}��l� ��?$U��RoQk�"�n*�O�����tA��H�6���o��\��>�`�H�U�3�u�L[FI��%e�lS�2�9�U�~�F�'���9���:+�\̐��Aq�o��Ր���!�o/�i93�6F���ic�V�x��f�q> �PC�|�6V�@R���_��{i�n��|&:�Y�h��i௛�.�qk�V���g�����ff5�MyDnY��߲�Ӡ���݅�­���3*'���LEKv��3��+@eCN���'A��$���zwCxgH��M���t�?:��u�C�Ŏ�� �[��Fl
�W.���'EaX�PU�S�!�"��\zA�J��YաP�I킚���_$r�L�+������=�ㅀ$��FO��U��W×���Ϸ�2ؗ�pn�J	=&��0��x�Ey�T�T��\�s���'��mӀ�A�>��s�j��J����{��6�H@X-�ʺKxN�r�T�",�U9-��Uc�Wu�j�(U�@_���_q�b}o�X�(�/����x�^�)�Rc��`DUѪC��;�1��1��s��Mf�~�3��	I��߆i�[᳇җ�B���^9sX�#I!������[���b ����Bo�u�SATRqfEs��7@+.�E�⽞�_�ic|p|�����P�d�d&.�d�M�����־S�������X����3�2�-^�5&Sȝ�Gި�G7�@�_��"|�i�w7@��.n�Ed���*�%T�՘>�v�u�8K�m�3f#R,�*k�B1�_�����l#�|�V��k�悢'�\��4�j�ğ��fǗ�ڰ�	�S�X4#�A�>H�P���e�TPZ�օvJ�^��l���Z,���F�ٛ���y��TS�4)˼)��'FwS�tS��Fe��곖�g��Rma��vFt��{K���h�E�Y�<��Q������ֆ��E}��r�:cѮ�Tt�U�EN���]�o��Tǅ���'Q(��W�k�<}�i�}P˷��'�I�� k�%�����z�6`�`LY��Mz�LС�!�KY?Ӝ5i�*�jV�+i��7?W��$������mÂ�O*�7�i�D�>'�\em��_6G��}�-9����y��	����K���X#���Z��\�f΁w�A�^�!�f(�o���O������D.���7�)�-��#2N�p�Bʦ6����v�Mq���S.]⬌L��2�@-,���n�`![��.~B�FF��~�R��@ʷ��,r��3�͙�S�E�S����|�w��1�� op�?��;u���	��� ]<���C�n�*ok�A���j@S�A�-��`�A#�qa�L�Ι�"�5�Q�^� XN�;T{���a�k��2�U��E��Gy\��;�r��@+��4Y`�iv�c��ޫ���Q��u��@+bq��J����ީK���X4�\�DC٭� 3�Ժ���SA����j
�8��v�	n8��O�Y�(\��$) X���N˂J��gW�q�.SO��c�s'��u�6��|�.�S�SQq
���F�S}֫7���lzA�QM���t��)����O+�鎊4D �(�p����W�|�w�~Gr� �WC����C�hDE����m&�#�tǧ����҆�������N������X�������Ł�@wX�5W�҉%���ż,�4Ն	��.��9�$��7���w?��kq��Q/�b���,������ˊ��_��X叁iר����{������'�\���8�.�m�q�A�8��	)�C����G'��TZ��s}�d�͝V39����� �8$���e��m�=�w��:*���� 8@C��'|>N} �S=�m���X�a���;w�4�c)%k�`��#a�2�4���lZ�v�>�\��2��Ex�rj��f]�t����TM��-s����c�;\6A��w�+̦HT�b���0�X�y)N������J�>�����td,��7��G�j������<�V��*3�1Eg[I�H_32����=G5�-�,]膹zR��wp�K��n�t�痈�މgu'.���Fx+h�K�R���>�B(w�����=�eʨ��bK�P��፲I�p���Ua>J#���=�1������n lY�e�'���/Ά�l�F'�̜�F�kt�&����G�Iư��՛�:�7���?>�g�FN\m�_G^��1goaM������iE}�L �Z���N��G�3��Y��5z��H3d��� �Q1��vdJ�ۡ*�o�U�B��l	�P�>_�9=�x��1^�D��-�9Bw����`>��f��U�^�:�Y�U;�̝�Qk��w�)��&�[#U���G��F��)��m6LAH.Mmp�e���v� �c]�)m�.aG��G��̩��|�`44�p��]�?�A��6��_3�h;o'sx��C>���)��s�XƼb\}ߏ�Y���*6��)V��r��2`k�`�k������7�.��'|q0Xj��������&P'����2�3t�b>�ɸ�Ӱ��QF��mE�s �w/f¸Q��]-��Cj -����a6� D02�[Q�b|����ɍ�İYK6hxp!�yr�l��~�a�-u��^���5p������9LHu����-w���d����;H�(�BN=H��TBbkk�`Iذi��@U((�������ϊ,[�{�ӴM��ޥv5x�'�t����f���ش{��@��Z-f�4��������ժ7���皎=諽YI��ςբ�jgri��<C:���;R4� #�@M�BA	o��ߍ��ִ��Y�75�n\Z?�S���S�+���� [��1�������B�Y�ٵT�bq�_	�}�ٸ�'�����,)NZ�.���l
�wI��w؇���ږ���Q�LqR��:xWm��ɗ�K~�u#@��������L�Z����ˑbg�������M�]=;�ui�56�Y��C�r#V)¹Lld�Tŵm���/�3
D��j����$/Rdk��Rl�|]�/�)ݮ�1'X�@O�$�5lߤ��c`�0���f��Hi��,�2Hd� ��r�F6|�f����E�N�Z���&5b�B�5oQR֤᭽?r=�N�;��"��lJׄ(	��h�@nA~}XɎZ���l�Hw8֭n��#��#�����ra2�
Ɔ}H�t?AN�� Ɖ���IߜZ6�5���_�\ pG[(� �>U
K�W���CT'�
��ku8��0�hW"�JbRU8^�_+`��$��An�GA|�.*z?a����N�K(^�RC�ZF�ѣ�;,�t{�JT��:���6��1P�� V�Lj)ț����2��o��XG[űޛu��;�$�m5B�g���_L��v~.ž�_�m�d\Y�����\Z���@nu�ϻ4��|>�78;;����2_�@t�T&c��s�Y[�G!$v�9��xG�@[�1?�h,�4	C������B5xwJ��|��h��YB�c��)V�w��TI�R��R*m:�j,qi�r*V3�vd�9p�<��C��������""��ܲ@M�V��*j�wq}m�$W)�.Y͏���v��������$4��HÊ���18��Y�g%'�7�,'G��=e��+3��Jת�Q��a����Z�| J���I�,�(
H,��wǰ�PT���Q$���D�.���۹�����#>��h`U��e�;-�#ab�P�&eae�d���e������&�����o��,�U�,[SstSC���MM�A�XTV�j�����<�ub����O��1���e+B�S��ة�zSR>��l�a-}���˪�<��	(���g�< 5j,o�-~�m��f`��}ݠ>1/iP���e��8��׉@3�o����"�Y3uP��%��3Ԁ�J�5@������~z��|	]�{G��V���qD�r���XB_�B*i�)�hf���YM��ƙ�Ü�0�P�PFQ���f�Zor��?�O��:��R���� )�}x��xŵl����j�&�'_H%Ǘ�] �*��Y�ں�������H&�>���_$Rs��ǆ��Z�6{v4�*��<u���w��KK��M��ńe���Q�ԯ�&�%�K��蘾�S;�2�c� ���#O�����.2�/��P���V�٪s�f�I�$S	�#�XZ��aB�iѻ_�F��a����J��հp���19��t�r��k5}&�y\�o߻�a��Hsv��|��!o�3D�*��ߥk�?���H0�S+�C�m�1�2.� ��$�+j�k�FY�L[ӈ+���M1[sb��ںg�X�)A��,�J7��<��R�e�f�`���/��}�/�O�T��'[y�bT�{�n����Zr:�y��}�_V(u%�N�s{]%�� 
���D; B{e���3����x��Vq��w�a�ƙ4�l�/u�2��h��_�+7�aTGY�=�\ J����y���{��Ѿ��=�W���pO��7#�����"����&(H�Ϙ�/x�י^�;%]э�EI���Ф�儘$�����%��nGl�<�ҳ�4s�1G�[qS<B�:G����*$�>����@MgE��c� ^b�W���QK���pI�Z�n�K�n�������̺��k�	t�ؼ\�&^v�6#���8 2t��?Wl*�j(7DP+��9�t	���(=��"�	NS���Q�^���?�`2��Qz\���f"B�6�&n{i�K��_�,��m�7z3@k��CKc�y>�}�wc����Ǧ��l�񇎄A>'F�ܻ��EA"#�ʟ7��l�er�+-&W���J)����vG��}�IՒi� U�*�>�ZB.*�����	N�������f΀� �I�}���Uɭ�%����B��]u�4�2i=r&+�?�~�!ǲ���V�#<Yx�vX�@�1U�@,�"�� }��Z�d`$u6��R?�X}����"��+�����5�ҵ����V�J�6��Uy�#MV?o��%�ӣ�dP�<��K�^����	 ��/�5p�1�-E)tK�}��<��#�N�O�VY�������b�B�����w���G���C�U=���X��t#'(yh�<��﹦Fhr�q̌Џ�zaE߀;��I�t���E�NVwM���럝X��W����^�a���
pm��[�|'���i� �2pW뛼�פ~���VO����쒤�1i��Ȍ�X�C�5��}���?��n�����OݗX�6�s�7�I�v��W�]_�Z�S(���>vE�E�an�x�(t���J�\V�L}��I���P�����|��,�LO
�(#�Mwj�(�V��!��=%�J��B���e���R�д!J;�+���8~��<�7�B�El޿�8�R�� t|�(x<#Li �����CH�@jD��Ai�ug�'(��~�ʻ΁:*����y��Ejہ�=t�{�(�՟�Ĭ�X0+�񒆐W�y�����.d�E�t���f�]���4e[�ơE�ٯ�)a>���4�j6�x����fB z,��;�L�����p\�IA�ʊFO����*S�OסA����E}ힾ
�9��5�߱����?,ѵhV��YD�Ʋ��Y�rK���q���=�@��cDH^]A�xYu��֯(R��3�(�{hNx|!_�X�Ń����1�����0D���$�������(�C .ӭ�'�p9,�ӫ�n���
/P)�Lj��􏍅�<�ѷPC���z���HsX�u`ЃJ�����o��� ,_��o������1�L�&M@�����1G���6]c�aL乿�3�f�3a���E�8���~~������		�7��
�/�x��6�E�����M��o���U��mT����2=���/�9')�K���ޖy�'���ڻ�e�|�X*��O����?@�q.���.�=�Ĺ��C�������F�F����A4y�H�q-F����o{~����
6���<
�3Ө��Qff�7�S��,�F���q!��4FH�"T�ƫ�i����z���_І~j7R����8\���G��,�(l.��T�e��n4Q0�2��c���z�ɠ���l]��K����~��MJS5��f�)��7��|�?��ZO�`{����0����Et���Q�w�]�X�P�,����(F���(tL�T��{����L�`��w�2�n�0?�B�`%Nv���Nw�!h�|\F��|Xd8���[z�a'��黍^��A��j�o��*f�r�!�� ^g�eZ��/��F�L�7��LMW��6���3�Q;�B<�9Z ��3��6�6?HX��ϴ��#~p�+�S�V�mdH��m2*�@ۨ���|v��,����J��硝�� -s��Z�x�"��ٞ�����@"����BO��2Q��gZ���֞X1���ᐮ3���ds� n�(����9��������~.JV����N^Qޓj%��qV�3?���jG~�DռȲa�!s0���=iT��ލE�P��R�K����J�lC ��G]���L��) ������yd��N�3N��u�:ϧ�s���jzй7
ι����i��Am��=�υ/d��ze�uG0�w�c�,�a�#	�1�lgE{_�6&�2��~n�Ęt�w>̦��k�[�֧�阘���V����5�<�yg1/�̔Lxg�.Mn�dzH8bo�@�6��8~ԓ��a3�L��R=��s8�<�{t�F7"�QQ1h��n��9�)N��J]o��A�Ŗ������w��#Ϭ�#ȳ���:�;���6@��r�*S"2q]#��g��-�/=�X�WG^�&���*�
��R�����n�}ڞ�\g�,{�,����Z_I��	��Q�s���R�ȫJ=2QV�*C�@����6���m����v���5�����u6���o���xd�;��K�eIL[�1�wݛ�Ͳ��U��O^�涷Oc��*���y�R	1����0#�c��r����
1�� ���|S���b��m��o=G<��H�}���gI��7�[t�%�	��h�QBe�J+�{����~^���2�7��'~ߔ�7[^�L�$�K���J�Q��F���k4�n*�$+��
W�������@/îs��8ݶ�I�T5v{7�߁Ϗ��Ou�/�@ύ)�6Es�?��Z�XM�,�#���3#�=�46�gU�j%��5W������ц�sG����W��Q���J��((���6��x3��D�/*��I̴oO3nѠ���Zu
<�o���g1n�^ݐc��9�pN���~jy8�D�:�"�?��%��ģ7� a�+��̂4�s��g���M{dg�0��o�[Z]Ig2T$�i��̎ ��b�*���j�/W��a��'����S]�����	n�N�,��۷�gj���_���(o� �������l4��Fl�gȽP����]$��XXV��:�s�йfe�C��7�o|�D���Y�oB��K2��j�����l�����C|��:��`�9MJ�f���c�lI�"P�
�r�"9![]�z,u��N�կϡ7X�/ׄ��|�2.$��E�*�S�L4���Q_�U_c�gI�A�����/�o�cGn;-T��Y*Ps�^kK�����X�| �`���S�s3P��囼Գhe�Z3��O"��-ʷ/
��}�At
V��P�r���z�ʳk�e0�����������π� ���ĸsd��VW��o��ڸm��Mw�(Ŵ��[��¹ �X���|��5�˄Z�1���j˂7�vL.)+ʼ�##��<g���m��f��hŕ�֋�
/�URY�}����1,gz(� �ΊN�6����'S�$[;��׭R�+���Zl@����
H݇ȼ`v�l�s�]c���-Fl�Wls�DE�����M��7�Cv_K-c0>^M�2=�z.�v�wy����aY�B�/b�'ZP��k �u�"�Jio�~�FC���Q 2'�7�FK�`�CL�Ş$]7w�oH�ۥ��-Cn�9v�7�}�����0����s�q����l���Q�8����v�F٥U��t�F�W��q|b���n�ŭoC9��*߿?A�7�s�W��,��ү�m�ᗛ@}y���$����-�k�N�T���ׄJk�/`RX@Xַ�D+�r���"Rv ~�`�R�����o�^�L�a���\���z����7$��>�0�V�m�tP+���h�nf�j>��dE�#|��ֈ�y��	m�w~a�E�:k����(�GE m�s4GuQQnI�S�аR�4��4^�_m���d�z�c|m^�$��R�6��'Jހ���R� 0��8�O���nYw��Y.�����%@J�^�|�mT���qPh2q�	�ǁ��_WڰT"�u+$N�cw�ٍ"Y0���R�Yo#�V2X����rlK�0pp!F��:��|��j8E.Y��Į^�-{Z:K�J]�;��Ys�{.������V/峋��w���b"��e�i^:����-Z�S�<����;�છ�|b侕Sa?��!$dAN�
��(c*W��ߊ�ՍV"�	�@Y�Ф~E�-��u�L�������fG��moX���CYE�I��V����v���I���n�q|N��7� Ev�?J��f����S,BzR��lDm|��B]��W7�W É�v/c��T�r[p�5 	�֜S'8���XA)�3n�����K�{�R��`�^�k;�J遹�}�y���Fk�j��� �+���qQR+����~�v�,l��U�=}���7����O�I3LJ(�:5���f������#`�,��eZ�g]��nӮ;#�%���-�>�bOI�pY�$�x�7���jV�2iX���Z�:�AFJ�O���J�b���/������E�7����3���ʣ�^1���qńkr�����T���[�B�h�՜j�۾o�-�AQ�3���,����[hm�O�
Wxw�C����U�t� �����KN>��!D$�:&�?aGeqFs1����(@_�jEn��ǣ���#�R��~ۂy���Mo/�0��Ju��ʪ��m�Ԗ�H,^�	���!�?&}@���c>@;�R�� �[y��':�w�6�د�c�� ��v�6O�ܒzf{T=� �m�>Wh�~^�H<^��w2�$N�y:�a�xa�I5�`��yB��xgTA;�+3>:�����.e��ͣ&��e��k,7@��b�,�ݷF��mʱq���g��Q\��Ñ�9b2ja��N���gU$��˧;�k-3�%3��P�Z��w��s�L���)���O���J�`�ޏfv��|����Q��3�__��ކ�w�r�!U�+{�YQ��L9t��R�S�s�����S��9k�ʓ�������!~�a}�.�oz�'s�2�p�Z6L���
e�j.
��?Y����#O?��cXn̗s�Dݷ?_��P���+oʊXd��M_��U�De�5J�V*=u�m�L�d�(Dܢ&��
8R����[���>��[��ܗ�[KՒ�݁���O�C����>׵����ә�����B���q�T	Հ��/�MT50=i��
�8s�C{��!��Y8��p�T|w�fzG��iwq�HQم��:�����*�Գ�����V��	�#R���wCp�%vRp�H0W�U�d�){�O�2��'�4;�a'~t��/�e�)]bVl1a�Rӣt+�fp%˗`�ޯ���v�x1aS�׆�+��.�i' @V�ӱ�A.���O8�H��F�0��#�0<�a�*:J̠��T8�J��N���]O~���o�ad��R�o 0<C��HH82d�|ǉ�4�
�U����u�[�v
�nc��1�����o3L�X����M�ҁЊ�xB�n-z����.�"N�6�^(�����~��#�6ςt�iT(V@�j!g^H�.=mJ�v�H΀��5E��}����S���r\��]����nAV��o?�zW�Nח��f�E1�,S�!�c�p�d2qor����`z��+?t;0�U���SK��	J�!�:�dO.� ���r�MZW�bt$���������
�6fי]�4��8Ȼb��U�%�a1*۴�����U��.>�[e��,C�@m�������_h���e,1z��5��"�sm\�:�-AФ���zs�H�+A|�q�"9�������8&y�Xo��m��qw����AKt��k��',Zj�#��^h�#:�Ϩ����;f�Q����q1�+��D��ʱ-��O4u`�@*��s5�e�p�lE�)�\8'VɏJE&���1�x��'č�U	:DA��3��%����ֽ��Z�H�{f�+�����eYWg��njOZ���е�ŭx��	�\ë�!I� �/���=�݇U����^����M�|ɽ�)��dn�=|rT���v���	�a��27�0����js+�^��ͻ>�d�R�F�r�aqV�F�#�P���Ԃ�	�4w�5]�!�<
wf��Χ]��eR����RL����0Q�Z�6����y-+n�X�����?�u���/�z�;P��ۅ�Z�Λ1o6��Gܮ���_n��k��LQ����9�����J���"M ��G�"m=���*��򺩰02f��h5]̻g�Yx��7Ԟv� (WcS]��a�J�$�H|=B��x|P�Az3!g����Y��g��;�D��s��8���u[��*!B�0xUקDDp�LN}�&�/Q��s�6Ͷ�a�c���a�Eo��W�C��F�/{�o���K��fh.	�חl�F�ئV�a���S�f�����ׁ��P��3fа��y%�E+����;nzm�ڱa��z�~A�? :c�؊�����v4J8��NA�mW�:���5��}��K����Ϸ����Ij}�򗴽�̺�ҏ��oq�:���}:Y��d�o��	"�ȉѨ⑖��Unv� ��5����x�<��Rj���%�f.�A����uT֒[#�Ze�kۅ-����
�EoC�T$KWK�
R�z�h�e��q���>���{�n)(��)id7k'��	�s�v��ҁ�ߏHT��������tP]"!�J54of���,���("u�.XƪT`��<�Wџ�e:Xr�sTAy���V+<jNNw��Sx��,��.&Y�fǻer�������Į������e�m<�&W7�+�
X�ٙ���9R���F��
z��K�JR���'R	�P���B�@����ǲΖ�SU�C�K)���
Qnc��3I��
���:&#a��8v�2tt%/�f���M�����f�p_�	���w1�j�Z�
�b��}B_��c&��3]�������g�#|}����S�;��vG��q4���ڞ$^��Fo~>��E���#A��r�Q1������I��C�;6�q�����r�	\P�z}?x���x�D�:�sv�\�8Xr�&6Ϗ���K8]j.x�B�E3⑸���ef-R�w��63e�8.��*ï�mJ�XM4�+��yq�"�
��U�mы4y����h��,�#.����fc�
+E�e�0YD�V�[�l.��ۧt@����I���$g<u��|�>c�\]���E�{�얛���CnY�K~"��l�	>����iy��(���]8 =�ײZ��ݬ���d0gI�	��8�P�8W�q�Q�S���+�F>h���I*X��Ss������:s�߈�Y]�@'�K�Κ�y�ntL�6d{��]��e�]�E���͵�Ֆ��Fc�++n[dW��6ɱ/�N$X!��#���r����S֚�����ӧ˞𨝲y��uO�*q?rk?�J9[��~f��yb��! �ݯ�+� (����B�4�bՠ?��=��?g�\FU1�˔zC.��*�*c�C��F�9��W6"\�sF%�����{��\��n�Q�V�P��g*������Wb���u\ǳ��^��R��7��B�&2����"c\㋒؆��d���`�sЀD:�Ɍ������}�SQ��"�ŏċ��R�q�[�08�Z��L�|��u!z�����w�q�s:6ؖ��F�T��bbS�6�W8z[��\�H�h��t��!q]Y��=j���s-_e� "�l�;�e!���7wι>E�vܕD7Ҥ��@j�fH��eP�𡦷��Gs�NȆj`8#])n�g���$�&�x����+��l���Jw(�V��3�)h�_�4�A���K�(o�'zm�0�� !��>*:������}��(��A4%��{���g�2z�Zs�qb]ߣ���J��"�<��gW`�J��*n3�+�u}�$?��|�F�2t�i6�G�j����c�/�P��Z����}X��}��O��=�X��v'���4�ݺ��.�w=)P��zWo!&�Qju�Jg�*�h`Ї�x���!s ��ӣ�'
��n�_�c����Z�� Q5hnb�}� ��'5b��7�L�6F��*��`AJ7�:�z��U���w*��/�����˜Y�rz�6��T�� ��w���CBt_��?�w<��� �)��I�8�`(�vPy�AaK���x�}4v�#��G�N�! *5����@�������d�����`�^�O����U�2��1~�'��@�A����_�ܯ{��S�>���	�?D�-�~hRh�+hܙ/o��Q��6k"�Ŷ1{F��VC#���{,O7�Ih���g���e�B�~ϸ�(�nt�z�}O�-�͔�)ʛfTW�������C2	~
�#9~�[K@\8rN�IMr�Ry-|?�� �~`�	���bs���Ч��Ny��-Y��^ɕzz���$0-��U��rR��Y�;җű_�'~��s�0��`�t�a��n�����k\5�n9ϔ%��l��gԸ�ۚ*���=Iu����J������qse�`�Ob���.�캘9��}���s`����y$�������,}�yjLR�V,��}����2�����^Չ(���e�9wi�3�[+j���:���ɠ��E�V8��u�'�QW�ɨC)@`���Ew���|^k��>�AR�3ˬk#hf�k��x�ؖp6���0���W�]�G�n����|�zdc61��I#t��Ո�f��(E�c�j�j�3a�3�I!C���F{�m��T	���^ɕ��mz���ZKٝ�^��$UW�w�3��7y'2Uڱ$�ұ���W��UE���n��0D}+j�`
;���'Iv��@��U�� �@MZ6���8,�۲�x���q2��1�&])�U��ܸd��ppސQK��5#Gd���n�J�Wy���R��P��POH�3C���gB�>X����>��c��~��:�.&ʷ�(�07d)HDeS��|��������&� �������T�S��\d�k ��b)�|��]4�/n��c�P�]9�:��9��e�F�,z�z-��ʎ�!V�qT_o�a��̸�4S�]� Ivi(U"nw�ް�ZŴ�@��28�bOf{\N}Ų(B��x�qѽ��w�����#`���7��A�$I7��I�wH��Zj�h�Ă���Qޢ{���7����O=��篷8�� ��]B� ��[�s���-�^YU�7�Y=����Z���c��ଖȤԮEy��B��K��B[�7J.L/����ۅ�.+����_��ͫ��}:���&,�.a3�ڕ5N9�D��!oS7Qu�G�����B�	�<ʊT�� \vI�t�+$�0q��s��a%"Z������N���342�xl7<�.I�q��\Cm� �i9ۍ5z���˴�A��_�%��h�f�����s�2Ӊ�ˬ2z��;�FQ����Pa�mG��u�5�n�� �J��;C����_�+�G�ᝢc���y�CD�=�"�%���O�P����*������٬�n!o@
�9��UR�K���u2f��x�z_�$����	"(�:���v_@���� n���m(�JPs��u�1�����7�^��?��Ԝ�s�|n�G-Bp���8oy}!_�@	���M�K�'�&����	�F 70��^�4f�J����&�eF�b��#��G0S$\�n�x�'��"5z�ۺ:=�/5Պ�X��mZ�뫾x,�|�eEUK$����(�7 �㼛_`��%�<^�=:m'5? ď� 9�GY`�wO�SP��,���.�mhC�=�ww;����a��ͤ�]U"/��w��$�ҸY�j˫��US�(	�4�b'Qg��������N'.�#�Ṕ�e��`d��+���r;��+�,�z�,�*h���G�O�V������ju�9.�PƁ* ���HB1�C�AR�+����8B8���b|��M���(��������,F��]D��;�x{,�p��ߤ��f�3MǍ�dU��,��W}hi�7�ZI�������,����3�Ҵ��b�v�m�������f합C2��Ǝη��h�G��(�$��VA3<2�i�1J�#��0����0��M�:Pv�:�=xac��#k�=��&�s�s�7 ��S�7	q�%l��^�w��jJ�W��ʌ���S&���Y��]����t���cJ	O�7>:_�Q�9R�?OyЗkH?A������ܗ�t�<�v@d};@ѓ�ev9Α�Jl}�/�H9�����ޖ%�Vp.��sxn1!�ZYbF9���۾k�֎F���O�.v�s��&u0= Я[Rp9�Xa�D ��[(�|}@dRq���Ix�C�F�y���*���N���
���DF{����g
�[O�)�}�K�%�ջľ�oo�=�p=+f���%V�;v	 `�����nQ`l[:�V();}���V(G�d�m��[&����2�"������d�KnB/Af��j�G>�K�M�+�����	�Ls^l��nή�ٖ%y0Y�S��Գ���]�_k$��O���ֳx6V-���"?�4dA9��ߠ*_�ȵ�H�ϒ��~p/��v�ft��#�ra7g� � ����tg��x�^�b-��!� i��8�#�j�6�RN^�Mdb+kkm���ŁV;)4Ea#���ӑ��E�)��:p^�L�h���~�{8 �#:��%V��եd
Mp������*�6�jD�l���U���e/~�F�h[��3�_�5�X����N������������2��D(Rc�K7[��E6��
�?��g�@�A�P0��eT�Oh;�D���)+�6�z:E�h�N���	��w�t���m��%-_SnQE������W�!��N񖅭��}�9�8�9"���`�_���Zӊ'��p�(�F������i2��?�'5�V��R6��7���'t���S5~�=s���@$$y��829�e��yZ�(��nD�fM�MiZ
���V/�ݸ[��;\�W���T�R��t��-��ǴzT�̏�����B�N1�?�u{��S+J��6
����A�D��ȣRtZ]{���e��-P�fr�:�i0~�o����q�I���3��_��8My��=D�E���H�W���f��}���flT־
�/����2�����C���o�7�+Ӡ���������̵��Ҹ.?n6ԧI�F��<e��Mu>q=�~�>GIYek��\�9�/D�K7���^,�Dj��Uj:�Eܿ����������*
�q ��S�`.�O���Kbea�1�(Y:�唨\5{�i�q�����,mR�n�+�b��q�5��T�J�}/� ��PɘF�@`c".�=��Z.�\� ���iБ{T#��ta��-	�l��-B(�8%x�r0��v�ʥ���u(�����$��Q7�����.�P�.\QS b�y�����������-�p����%�6��Aʊ+y��nVU���n��~y�W��#�+Ng�
&Oo8�������cZ��B�?r���.�Lk����_Q;?��jP�՗յ�7V]�� �4G��q���jp���/�nҬ��{Ȋ�6"�:ڪaz�U����.�q܏S���3)�fp�s��l*�h�GhzHh,GC`,S��lJ�*C�M�Vǆ-�h%�M�=���,���7zgf��O��!ih��r3�
j��jm{�
��w���v]J���u$Mr!���ѿ�'��fMZ�R��$�:FmQ�@󍠶�eb/��2fP
YR�����<��ڈ�6ʹ�U|�O���X��Y �KG���*����Կ�b�/�A�i�_8,���� ُ�u8�P3��;���>DyD�w�mG��� ���"�5h�O2X�u"Gj��E���W��Aú���G�9j���=Kk�%'v� �mH-4EWƻ֦���-ӣ �S�Nҟ¿��p ��M���h���jV��,��-�ꁞ�i,P9b���%":�g�6���$�b5�b���l�l��dQzB�M3��&��@��
F��\�xt>y[H��!��ζ�n����ή����hA� A�J&�`
�{�16�Kݿ� B�[hL-�:Iq��aBjv�#�=p�8�ً�HeҠ:���?��&��xQ����𪞸�`Ǯ�^�@G�w[�.="x �ઠX5��h�o��f���rR��+VUl�.2ηv�b ~U�����
Wڝb��Ӄ��:�R����i���,?����X�@� ^{�c�8@	�,��͚�ËXOA&o1%�v��Ӎ��nr_�LG������om�V��c'\;��]:�̗��	`�9pSs�f?����e�#;��#����c%@2�9u&ڱ��:�[CQ��d�r^��vW�=Ӽ{�'X�������܃���z�������o9:�i��@�-��d�f�5�GQr�2�e���Q���R"!�Hb��j��f'OQ�^��z1�o��:h����%���3=����ۂ�W*u��AeMh�&A�C����3SP���9C���,�f��X�jS�ByQ�>/)�9qWF��\���L�d`�9���;Y�AF������3'B_ۭ�C3W�������E�e!�{�k66��?�A�A����.�y��G�u��株g^�ǰ�n�Η��=��:u���}4�҄�&=�Hs��q</k}B��T���-T�m��h	s��i�j�b�ҏ�������M��NR��kM��5/ql�bFj�!������/�����+�aǥ?�b�=�i�p�=��5s��9H�95�90��P�'�����Xi�N�nK��R6�����wV@���A{�R���A�Y ��&��(Y�)v!�r�83 ��:�������bq@h����V�;1��'��T�n�<�$3��,��������+�{�D�����m@P��d㬣rK�q�n������r*B� �^<�N��zj�+L�0��#�X�*Ŵ����!K�a�nT[�0��F<�w��fB�(����?I
����@�2X�ᯂ�I�V��L�RǒE�
��Ӗy�;�
���qł���bYߩ�X�i�e��'������kt�`P��/^�'ۚ��O:�� ���]`wW�{���&��T�J����,���5�Yk�v|[;+�Tv���bO,�J�1Tv]O~$nFJv﫝�����a�WS�wM�Z��t�@'��8��v��Iǭ�]���T$��U���4֜x���X����nk
�R-�}2����pؕhʃ7��oHu�P_. ��S��� �G�
�&ԩbxx�1שj�`�4n|j�ˑ�Mq)���LM��:�d���&~1w4��{/����zpU؏5F?���/r��.0�ڿ���Ɣ�P p 都��G���QyDŧ��r�oʵ/u;b��,g��Ax���{�<Św)B�����*sO�6#����k{n#���j9@I��	q/��Fb�W�����I�d��������
�"��]*�� �k�f������r�<O��-�3�).���#���MC2����>���>����
/}��?%�n�c�O�nya�TQ��$ҷP�qeA)�8'�J��A  ���a�_�7�eW��.��'�ujͶU�S]������RP0뺽ћ�և���,�Z��-(�q6��9�[���3���U��Ԃ�j�r�)�4��k��Vg��^u��f^z�R���]��nшm�+��a4`Ul�Էdҝ��y7�r(��,��E[#�@���4�/h��i��{���7��?��:��.9��tMKt�8���x@K����o��+Mwg�h����#4��tf���]�l?��5�G��;K4Ɂ��)c9��H^�*��K���6񫵰��I�(o��l��OPq2"A�Df��enJE/�_����h��&��6 �6Os�%r9�V>Ü�+Qm�B�(��`{[���A�Ә`c�D�n{�].�{+���6A	o�-��i�(�8��&u�����Fϔ�QlʚD�J>>	M��Rq�YSp�y���zf!�l�g�ۇ�L��בY������KuJl�P����w��J��|��>4ׇ�u4B�H�k:*���AA0$M�i��'�W��8J�.Z<<OKn�t��_���!fd��7�9�.��UW��/�à�V��uc�R;w��@$��L���a$$�w���é�Y�+��ݘ�x ;ShxU�z��
5���&�Ϲ��O#�8!� �{�?�]V�I0��YX������ē��>[��%������!M��~�I]��{�������/�1���Z��6ǵ�F,��d�����^��3�e���z�P��\�"Fv��벲x���j�42ZD2� !�:eY��+���?��E�{���L\%��@˼18��W��&�4�oЁw�[5�1��Z� ¾���B�R�M����JJ���J�X�I���n�qZ��#_�als
�Gw�L��{{�S��Q�w���;�}��N�U_��iz��ή�K�(.%�'�		�X�C	E�kn��Y��'An�|���Ο�v��	�����t�,|�N3y�P�\����*q	1�o�}���ц@�iy���b̔dT*K\���r�wv��u����e�<�����)H�%�< s.���BY	�s$���)3�WW���Lb�0i|��j��s��O�}A�13�Iv
�Na���-���ڢ�S�!�Ez��V�Yi��~<;ȆԐ��!�{��W�o��`(q�U�p?�hL�VYl�:������K�f��E˴���s(H�9+��k�������3�� �7t��`qjh�q�38܎��ÿ��f*H���3�[�sE#�&�|���M�R\�bW�P��z �4���j�Q}��
����rg��`����~��Z�JH/��\k�����!��ԓj�{g�3l�b����v��a��q�!K�Na�������_����DUɮ�IX��o�j��o�0u��e��v?�M��4��3��E�@�=3vH.�!���]���&&�q��Po��!��4�
v\v��A>���<ƎG�J�2]��2��5����j�
T4���Y�j��}�.�MH���������X��#���9@}ũ4pu�=~���b��\y�rty�H�	�o,��㳙i��$,�Ys�����s�9�w*��\��p�12��5+/�M�2QfqW���0<���b}T�Z��;�5��ˊB�"~r\��`�mv�]'�˩�6^�`#D����.}��w)��Yf��ݍ���w���ܺgknMZ%�&��T*���A��8�|L~�Q�w�g_��"��Q�6Se�\0��Gˍ&�� {e+A�I�.�p�n����s��<��г&�1�~(Ղ�&���G�Ч��W�vk�B�V��|��}�i* ���ߨ�����Юqz�I�ƨqj��}I)ix1W����!j}���C�L����C���)wk�%�L���H���h��M:fƒ���ޟ��A��'�m�}D�'1Kp�O����(&sDN��b͟�H�.nތSM�C���k�5�E��1�M+���NWff�F�1:��6 %ɝ�6ZK��z��}Y(CJ�����XQ��v}d$c_��>�F����?~&]*6&�;u�Гoǫ�w������!�OT��O.�:� ������,ԝ�Dw���p��f<,㇈.�7� �ÆG���R�QPfp~)�'>���?Xoη��2/�䔛''';�k��ΆDO�` ёD�iol��	��bOM��>�uP������}\��I+H��j?D�[�	U((7iZME�L'�z��GȽKgu��!�eo��Ț��ڷ��	��\K�S�kCh�<hOr��O''����Do�늩ӕ�$��V�La�a��H��E͎G�oƻ�����o�T�
F�U�5֜ڟNI�j,@���V�L���qi�@�������Y�P\K~~^6gf���FěҸ]�W�]`��u4���B�G��ch�JJ?�WT]n�?��(���3�������&rz}�r�=��uh�pI[`QN(�22�OߜK�, ���7��-�Aج-�
}�&i,e���]����yD�7�:=�MA��~�^D$��Xs�_�^�ºt�>��!ڌ�5�פ˱i8Σv���m��8_�{�{��/�8�]�M�E�^w Q�D ��W�����[�u��te?��'��hU�v1VQ4���,A����m4��w�1�;��?[���C�\ �~D ��8hY?�wL�'F:A(2 ,�?�LG≠����[�Α;0Ǡ�g����V�p��� �bYa�ws��i�,�nܙ@`-ҧw�{�b����<�Y!��qPMB��{�	;�i�.̎v��'������ `l5P1p�UA�*��B�<}��a�IX̐h#�GLFCF���7���qK��l$+����'��#,�ȩ�qr?�4�ە� ��T6d=���eqsd�T�;S�n����\��J�%S���E�n�9-'~��eMSg�>��ϿV���s�њ.�Qѧ�d��
%����KW�_�ZD��?R9����"���ʴ�:�2��vr�����5fx�t�l��mv nrs(L��"�\���3��D��^}��#>���6���t�^i|��Y��z��2I�~�d1Կx�wy1���[���3�����tT��3@�[�	�)�3�a�\d���,����2
�/�if���\��-�7BE���Mf\���'���]A����pXZ׍��i��:��k�n��8�E���'���]�^^+*}���ß�N-�*�:���	�W)L��e��4�oekY>AM<�+?k�,�D�!X���NУ�Q�X�$��c^ޛ�t��������fЯI��P{r���Z:%U^E�l�ǔ �7t��]�	¦Լz*Ǒ��!��K�l���t����ȭ?�c�N0��l��<���A�=��[^'Qk��"d�i��t��!f͝u�*��ͧ�`�̡�㸺�N.�+����X�����[hF�?Y���bO��ܓ�%WH�'p�KM��V����ŜۉK�Ȣ�"fSN�x[H���uڞ`lx��0`�ۿ���#$D�Ӡ3�4���W�lo���6{��f�,!	����rv���	��lTԍ� �l�S�H���V�S�eFjv7/��Q�襁n]>t⢋޲*��m�6�	5=T��^F�ޘ[��X����G�o9�۾��L�Kؓ6�0��Wo�A�jYP��
��{oQE7�t�g������b�|�����,z)�?��H:�_��#f��I=^bb����3{�3�U1�b��׫�t()��!?D2'۶�h$g��VȳOce�T�T7��`-V H�T}^K����@e��l�kߪS�￫8�
y��?G��qW�ӻ_BDP;6�3�~Br��5�v.12����̌@����sB7�:P-�#���E�Q:�"�gXK��O,m&S��_��.��M�ݣ~��u���!A�J�*�5�:���Ҥ�1r���	�	���]�h��5,¹���b�g����~�]��e�L��)�`��%Kw�J�w���EI���p�g���6��4���R�%�Г;2�OWI�F\�T�U����yZ�����Ԝ�u7KE��@��k���W�4+�(?P�OzF.���1cC���c,�Wm=S��I���Gz������>��5�`s����G]����@���<��� ��e�J�a2�ہi���*:{BL<,�M;4����9���k��)]��d��tp,/��B<��Uɺ�Fdڃ���ϋ]���<��_!�$08y�llf�n�]���u,u���Vy�%���ő��~
u��g���� @M607&���@����o�j���y`�*+���ޯ�y|��O�e��^���}WqCs?�I��P7�uk��6��p�1C�ɽ\D���Ϙ�a�[��0��"+�bEswO+F�)�ק9��wU=?`
��A�[�2qG��AD���nT�6˯�.��ԍ��&@P�Z�!�L5w\5G-��Pn���w*�����|q�7I�nH8�Iu��q֮O�}�Y1���D�[vb��4k�^��$a(���ЋֆWS�ŏ���o�/*�b}���=��Wav�V|��VR����i�=|�b=_:�v,�,�g��q�ÜXx�wȬ��_���Dj' V� �=��$s����a�0�:Sj���f�rKyJ|�8�P�Ә��H���O]��dF�SE2�U���_�O��K_L�-
�+��U���I\O�K�)@�<�)̙��C�V�����c�����La�o#���x���"����zCm��]�<��(�UW��k{�ނ 3�%/]?����/+f�Y8:����p� �_��
������+���;��)�|]�C�9�n(�*N�����^��}��K/�̶�b�(�3 �����������<.Q���8<l
&�jeA�+�x|Ӣ}#���ٗ��.M
L��ePY��ϱʩv��1����f�r c����w:�7�H�J9��0���e�7Dp��_J�+r�{ȌG{<;������5�t��vX�������~շg_����ݖ���J��j���l
+btuR�lQ5�ޖ��a�3��������8IR���O
�ʏc�X��]~�����=F�]
(?�g�g��f���g|�E��9%��zn�:�s�����ȅ�/~g`Y�n����	�b�_��8�@_(��X�ɰR�զͥh�W��:�g�RW���ۢ�Up�L#6��E6A�K*o7%�χ��1J�Wt������:�9��`���s� p�ɪc
�p �,R��m��ֲ-<� ���>\B�����ϑY��Y�Q �!Ϣ�l�A^ݛ���;��~}G*X5��$b��󢵔�s�d�'����Ck���B6C�E�=��V�$ӏ����t������.r��I�[E�\�wu��"]�_7�4Rro
w��WL�N���?��)�?�P&���	��泦�pV;�B{l��r�Q�������͢�eU=/:k������:�=�p��}=۳~���E���=�"3��{�cu�����
�5绰����՚ʁ��whӒܴ+�)؏�o��`M�	8	ZB�;�il�`�ІD�[JU/%J~��������u��mh��r�!|$c:ٷ�m����L����9��0O}��Kb���9
t�|`H��"�bmQn���������-:vvV�D�ہOT��oOR��յ�F��ĩ;̎�jq T��հ�.w����籓<ɼآ5��d�eӏ�G��X�M`���sL�5#��-z�L�饃��2.:/��Z���� ӂ�Ɋ�S=�������b�������xя2[L�kHaHpTG�)�W*������M}���"���Q)a��;hǟ�{B9{�j��WЍ9��M]=)Aͣ��	�,�]��m�.v�so)�?u�N�RfU3���� /jF���(��kѡ�u\A�ֵ�6)��R>_�	�!$B$r�&+"|��99(
6��w����ɧ��]<�Kc��|o?�C���#��m��H�*HUP]=��P�L�0���)�f�����򒉜�͑�Ⱥ�A_U#-���ȹ~{X�� ˉkR���<͢��o,�:��aͤ�%x���'cA�kg�v9�f�' q�Q3:�Z��P�+��[���U���R���7�,�g�5q3\jX�.�0|����]~�Fq�1�vd{�8is�(	eX֨cK�(�����1㼞�rS�"�3�	�/���~y�i�r���z���3��1y��(�Ezd|Ū���Mp�y��Jrq�K)��� �$P����	\�Dd9caivĬx���WJM��`�}���[1O�M�!$�#j��]��٢�֣�i�C��V+���2��\�l��ħ�2\4�˲ق����9G`4�iXa�(�n�U�>ș~#�ٽa��㫎�Xe?�$>`	a�Z�*�F+��_=9e&�ːe�����S�#m���5!	ƈ���]o��,2�DN:D`-:������c.W�;�5"�����=��l�>�<ۡ>c.���{f�����+[��"4�p0����(b�����I�q���ov�6.vO��sj�:�
�%��Zٹ�hyS�#��I`y2�B����O��K��~ �ҡ�c����H����5�>��(���z� &���Z.{Ď�d�\�=�@
�y���e���\�����/
�W�ι��n qZ��85ݻ4*"��(�<��R�弟���_!�v��%�SN%<��ng<{�݋u ��I�"���y��Y/ܧ���X�/^�oj�'iZ�K���=�ja���?�)��S�M*�MrLx���^�cR�Q
,��cyWv���6���� Q�6�|G�2�D_��mF"�AK������5}��6!e0q���<�A�ǖڏ>���3��G%���,^��JN�[~v��HYfnzAy�
�Ӱա�aH9���e\��S�[��W93}Z�P5���R ����n��*;a"�D?`@2l��L8q�#�A�?�0h�JS�M�ՖsD�P
��N+w�OD)J�[g����Ƈ��9��� �Րق�vW��:S�v9|TR�ոR���&�4��5T�>Q�Dp>��=�~:�$����n����.0�� ���K����B	����u�P�+|C^;}���LV!���ZX�Ĝ����k�S�?h+K/%LyI��.� ��x��TD4!�Qˀ�%|�_����#�����XG�Ҥ��d�U��e�x&+���v8sw�Хwn'�W98�K[3&�����O�Y�9Y?�%.?�R�0�\K��T�w�Ɩ�-}Z~�T� �(�YT���7Bl�ޢ��I��	t�W;�d�G���o����a�o�/���f(IC��.�ù���7_A%4'�[t��&�進�F-ڽ9\>|A��
w�������$�O���E_�gV	�쉮I0 %f��E��̲(c���))�Űܕ��&�����)-&�ɭ����S����9y����I\���~K{
���t�2{�-�|0u$^Cv�,?�hk=���;��T��������3��Feɱ��B�3o��l��@x���a�7�o0f�h��A��T4Ý���E�\��R����R㹷IR�K�9R�1:��.j��䊧1���>j	�e��VIi�kHp1��*���
��`��nH�dhO���"�Hl5����c�u0�d����6�c�Wq�P��N��P�g�>���)�Xt^:ճ�CE������Y$����41��Icy��Z�)�*x��7o�Z��vՔ���=}��4��_Usы�W�d����|y��clȲ���֊��q1����E�1�D�P�;\=s��74�&ʣP�&xs�9�'��&e*�YG)q���a�5	=՛�%�7�6�9h�,n���wa�7��P��8�o��#�xW}&�3�nDf�gllF]��.��C�����"���=��{��-��KX���$�Wt�l�°ų!����N���gW��q٠��r��HM�-���׊i��{y���΅�A7�Ȅ+'���t��@���!Ƥ�`C��d"mK�e��/V9��<�k�����F�~tS��,�S�2�HЎB�Ӗw��F��6��B��9V�=ΰ���2"Y���LR}oߐ�(,N׽N���UB���l�F"@}2���*P���D�+T�"�'�����9��m��4G��l�U>��/��{��g�We��m�_�^�߇X��bPjS��vb;K���&QOI����p.��߻�������&Xh�0ӳ�aw����+%��縧�'���d�OY�h�u4
���Tٕ�gb��<ia��fMa ���';?�����M++��Z�r��ț?t̝������"�둪0���-�rבY <��BLh�h�C�&���A�ZC�z`�ǿʞ0[����6[ɚ~2�J��Fd(�ZS���Tr,T���8�󩁱D�'*%��!染�nM�p�p�^Q�5��?�Na�bj�rl��yU��>�i;
� K�C�=x	��(��N��r���It���n��c��Y�5Ԗ�Y�� ]���V��Fۦh�Ȩ��]������$SP#�}u� ���1�����|�W�b����#��ݎ!���y�r�)*���2Q�҇_$rN��/m�?���Qa�x{GJ�/R�_���ǒ938_"n�jQ�C�^��vӱØ��RrgUs2mT<�i���Dc�u��}�N��$�<���W��2���f���lx���{��&�
!�|��dp���B@�d�&�0���j�n��"@��K���q=4�i$�3U��6d 3ƽ���C�iH�.,u�M����\2�,SQ��:&Xd����zC�הDe�U�fJ�t�m�xu��C>���"��'�Z4����~=>Wc���r���_F�X`S�b9�NK��;[����{�I�W�S�Ԍ�4�|��������^#Tu���$9G��{�縂��5f;0��#�_�^�6���y�8hTf%;�`$:՚Ȩ,���A}�&���ˣ�O�Dht����O���z�Ic��'i%ۜv��0�z��n��`�C:��',�.�W��^!�`�۳W�[pu`ۮE��;� �o���Yn����Ӆt?���]!��=��4��}Іd�����j����K�6��a�^u�]{-����K}����eH�Z?�߰-)=�nF֟M�I��u���6�׸�����7�W����P�����1���qq���"����t��4�r��̐��eRV(����p�����\�c%�?�1���R~�����(�7gi�V�7��Ї=`�j� F`��oSF��;N�a�7JI��HDV;h��1�����8S���o��7��؛'�e��ͼd̸{ѣ�,�9iBߩDBTt���d��喼�C�5Pϖ�xǢ�j%X��.p��X`�
Ny��ݟ�E���OT$��3f��uggߙaq4�J.��(N� �i�Vݺ�^��c3"�8ք�������MmN'(�>%�xk�u�k0 �T�I
y�#��Nݐ�y����J�Z���SR.�EW����0��{;����߿R�N��K�z�)=��*.�^��	\�}��gCs��wF����ȁ';�h���e�p'Q����G�'`J�_��E,��^�=�G��!+�>��d�	r$-D�JElU����������x��_X��!�8]1F��AhQD��3��0�$�%4��͒���M�[��u#�fa�	Y���P���d^���������ECZz~�	}W �� r2D�|W� �bs������^� P��`��n�/أ�cʈ��=_7�-�&?���ٞ�v/������x8�$R*̌���m�y�bY�O>8���}~����u�E͆����y�A���j��}EX�L��W��QL��v?���;�ʠO���9 ����}�]��j�T���1�.<�o/f ڀtp��e�K৫�x* �]�ֽ&���궥����\]�W�lh���=�Ml��)��a ^��ԇ�&M<�D��%#k:��Y������\��2>O�vؓ�<�8�3d֓Y5 ��z�u���t'�eMH�x+��ǰ'��i��c7�W;��w�L�������k�~��Ɂ�p�Nn= ��(cI5:��-of�q�@-�u�x�F�ɯՏI��U��u�Kk!e�P$D�� X��X��[_/�bN�*v 8�H ���~�A0���b���~��;N�s ����T)��,A�vyR�����~}"ؘ�=�1��+w�xƜl��H�U�N$�}��;o1q��^��t����Jt�Lh��d�w��#.�ݹG0e��.]E��a�J��o�0R���`��9�G!�ⷷCN0�
9^�U/6�$���07�Q���f`�~\�r~,|����9EŤc�df��$��6�z�p�4�������I�_�7Xʪ#l�i�k����y�Բ-e���)���Z�v�\ �X�/�#8�(t��_h��{.}�t�bIr�R�Ԋޓ��*�G�Ֆ�Zn��M?�p�p�|��"M�J��XʌX��Y"_��^�7��E��%�������>�oh�d����\� K3��fw������wΝ���Gb[����=X�tMry��	Z&[!~o_���#ZKTm�����w���3�n��Uź�ݧ[����b9GOqK#�}��s�B�Y���$i�i�����F�w�7�_Q�w]�uQ�~�N���U��0j��-K�ԝ�Vd����X/�JN�i�n�|�O�A��h�I��7o��ZM�hm�[�qJ���D�.|װ�>�����ګt��<?�	F*j��Ԗ��O���yJ̸��61�y�5b��n�OB_o�Z6C^̯�����^�w�qd@����u�9u������)��E��)@/���L(zEF-�^��
�"
�-P����p��T�?����[��^狏^A���r����BJ��l��
T���צ�����v\ʜ�9eJ�űb�/V#��/������֧`@�Xo"�@~4{��	�x>�!��x�qCI���8��O�y팒lɎTʼ�`�p��s����ˊR,�e�:�2S�D��ᡑ���?CY�t�;��Xq�<�A���y�If�	�N���KC�5h��ql6GbB��\�u�2�\}�~������lu٤<$R|���7�4� ��`���C#�N���SI���|k�O4�F<���~WVm������T%�ȗ�Iî�۵f\~��&�N�n�9T���Wǋ?��������~Q��=�>u
D&{pt.wV<�B��b�P���_��~PMj�ޛv�k3w��1�XN#��X�s���m��F�`uȢ�l��ou�ǁ��ީ�1�=��W$1.����?W��O�ራ*vfjۨ6�k��]��*��ya!E�w��dpbZ>{6�h�s�.�1�v��{Z���SEq��N#=,�x�@�%]bH�%i&�@A6C'x��K��61�@�@�4��Z��<XǠ?!@O�mF�{��:a�TӢ��~T�-�<��r�-�jU�Ħ@]�i��UN�h���.(XO�� J�r�3�}�|�V 7��#����Q�()���n�c�ˡq��;ؿ��q���0�b�'�y����b�sA�ǟ�D/1 %�Э�\0�hw@�:��gO:��x~z�1�χ��s�[����0�����	�?��H6��&�o��l\T@��Ԇ���8�N��˧*���q��6 k�o`�W�[�D�^2&)t^����^Z��ӿ�1�/oh U*���f\s������L��R	�Ɲ4�[D͓9]��70J��Ad���CX䆼�5��>��Ѡ��Q��sdC}m�X`�u��YAZ���?�n]kӯ̚Ǌ���A�v�ÆR!H���ůe�����<����2$��G�~K�R�M��Ӯ~>�gs>�C���wg-�&�TlR|��^~���<���=���89�s췱v	�݉蒆Ub��Pv�-�}�S�/��~�,���2�<��?r��+����J��
��H���xAE�����I�qBE�B�ߵ��X�'�d�#A��@��v���on�ҟ%��g�������ԧ�Bۛ@4�T6�2V��u��FILD����y��,�Pᓬ\���bx���>�.B�l_��rf��d�ٟ�����߳E� �����eqwC4X��6_]��f�"�����Z�J3HS~�@v��-*��7�c��!"k��%�X���s�"j��?��?�`!o��?h�<|P��P�A3ڇ�YDf8	
��"�[�겜�>��X�'��>��Zt��ܥ	&�I%tцPW�=�7?
>w�,�᡻*�Ą�F��Gfxz�&�)��$�ʝo��ȫ��:���*����Iq��d��|�.��XS�S�9��THkN����ܣ�_A@줩�d�>��	:��'��� #XxPLf��V H�#�Nd$�X}>rCU��,�xY@qy���[_���i]}f�o�$J�Ì��e,�2��8C��[�H�8pP�9}�R��B*5��n��ʏ}ѻH���+A��T����ÝJ'i��������z%͟N��eZZѻ�\	W�3e�ۅ�;*!,��S/`E�ɘ���(�S@�OZ�K��mlK�uH)h�|��cgd�]Ϡ�S:5$�i*��O����ؼD����o�(Q��զ������q�$ݵ�|�Gl�3�9�ќBC���h���I%���k���!v)��2¿�*e��Q��<��!Acǃ�NxiX4'��DM- ���{=��(I�~��"d6����b������`:r�gG�����������.���UiM����A���������5�K�W�`��:�W����o�w�J����*=�T09��Ye�_o�y�d=��!(=i�7��kRE��#�)�j [ͮ9dbb��}Q_�g0��-D����/۬z���N�ב���x�K��_�n]�=C9�ƫ���+��q�ɚUP,��e��}����eND�r�����W�V��2PJ���M�3.�=��[3[��!�������
�I�хq|>��	ЃE@hv'�PԷ�����u�|����b|�E��n�6
�F�(f#_;�=7�0�a
7x���si#��À�kRJl�s����K�h�J�mXBeVL�/�����EL���&�� ����|�T�6����SƴvS\(O=n�K-�x�r��\p�z��g�-3QO�����6BLWj�h�Ϟ0�µg��`Ň�Zn�@ػ�&��軆��n\t(��k:�s�OX1����W|YG�� ��vk��;��򇈫&u5���X���p�8V��Đ� L�X�9�}>;��OƗ��O���y�㏞��_������۰ɢ"����OL��n�0���!�:s��Vo���Aϕ8K������s��Z��K�����#�2�g�@^�Y�π����=�?a.�a|��a��&�Cf���h�f=*5H-��0c���/K\գ�����ԥ
��^���WQW904)����0|�c�'[�7Zs�f;d���[��j�F�n���9ؗ�A^#�]@�RDt�����
̫����<��S���~�|/�j�9����k�O�$����@F�v�{��z���ֽ	�#WU/�5TK���bd����W�Ƃ��FI�!�M��) *1���뎁&�i��ճ�x�x-H%��c�x�;��O����@���@l@������]��@/p�r,���unI�"�����;����m�K���؉�/�U ��D�M%+�ON�#nK�z��u��x��1����.c�����Y��5����n|&��T'��,����O�
�kw�׫�U�8^K�ʨ\p_�~��ԤŞ�U��4��	�S1�3A��#m����e?���p�� 0g��b��&VD�e���d�_�M�c�1F>R�����-9�
�KZ�s�0<��i.Tq�1ܒ�������Q�}_��࿕��t���5��B�r�#ø�ˢ�U���J��b�/._2I�g��<�}���w�j6��@�m��w，�։�?v�����2O�jt�F�{v�!>��wc{�p{�6a2[j���]?\b�c�r�K7��\|���lC��]K��g�U �>�E���$�s�PX��m<:�\"���b%n����k�`V��nt��Le!
9�7��� �6�߶��>�o��X�t��lh���B�o�y4��.��?����	j����q�wϖ2�_ eB�~��{�잎��z(^I�#Q�J�~��;����U�8>`n����P脏��Y������aGZ���\_��h��ònbW�}z��! ��Z#��Nz�vv��/@h���
�$ct��<�F��A2>h(��iܑܪ"B��:�Ӷ��u4�B�������Ľz|�dĖ�C�u��N;�(��0�0��Qx"Ke����V꽎��F�E��^6�s�
79�Q2�G�ʢy�Y��1�[���HY^�#�G|����b/x�28'y���7�@�h(�������pϧd2t��L��u���I�U~��������&�
���۴&`���;�BC;�@����'f[U�g����l)���9�F�-x�r/8~��N!䲓$B5n��0�3�SX1��ŝJ,rX����QD����������,�F;�C���a�7	ݱ�&9V�;��Os�q�o�`��~�Qln�JЛY.��!3ʔ��KO�����1��b��8єB͚񐪌}!;���#�ü��|��p�U�h9��$�������5ϯ���~~D��JtF�$�����I��`+D/Ȩ��(����J�U]?=ҏ�+��`�q;B2
L@��>����ak��^������ם\$ �6cO��"�qBI^�����E��B���AM�n��21�=f�Xsg�1\׮W�[n���J�����@ӕ��5�[��۰2�0~s@]4���Ie,�$%�>G��jH�LEr�
	@8@N`,�^��Q��Va yh+8�{�� $�0�eM��H���[S�,��P�Aޓ��{���b�9�����S9ྭ����O�=>6���e���]j9��e�bcL+ςYM$Y��q��{+b:���0����X����f���)�=G�����d�I�RK��0;3m����.��g�"��6=p��=��SU^�/�[f;+;`y#�$�P���S<՝_���r�c�"��9VzC�.��K˵�W���+0�|MĂ���h�hD\�"�q�(��d|���2�4�	�A��}E;-,��)�ajK���h
IB~r�ٵ���k5� k˳��6��݆-7ȇ����&6MC�H�U��C�w�έ��Tr}�\�O���ZJa9ldt�/�f���q��3��6�.SPY�U'�����G`M��k�[���!�j�;~�} ��?��=^��+i��	M�\y%����=xC�K�<���ж	%}�8O��^J4�ɵ�\�(R�(K�!$�S-�ĨbKi{½��b����p^��މ��>z�󊶓�oK~����w�9�+����Ʃ枑��LpY��W���<�9�����~Ӵ�5p��$�WѹCXa�:���F
���wLIʌ�5��П+v
Aqۇ��V֕t(����I�	Rx� W�2���,�}WZD�)�<�,�'�yT�]12�RH�)҂�v���WY5�6"���Ȗ���E}v鱂��ڋm���`���,���=z2)�t⋫��F�:RE�����s�{�֌J�8�;�%ΎNW�|�x���b2���[��2�*����5h��:D�����+�;M��[b8x.�,T$%�z^��"-O�vn*���b��������N���j��k�<e����
L���߃Yc�D��x	�
?��@� ��rm�HJZ8q�T{��*|s�E������[:RZ%[���Y�
Q�����:���� +�i�*`��V]�~T���-�(�*$�(R�����[�;p�޼�:��Vl�k⚦(�u�"��'%0H���XN�O�Z�TRu��v���{��G��z+N��8d���p��Q#h\�������񙈳�&��p�x�'�v�
4��:�שׂ��0�B��ȓHwKcH�F���є�-x�m���O���B���K�&dBBf�\b��B&W)2�J���b1��F@��Ym���0��q����D�+�G��ٕA� �}�T�Q"=�y&�'l�6�ױ�(=�E�y"&�8�2�:��W޹5����� ͑����j� ~3�` �s��í���Ate���#L� �Ć���l��z�7?菪�<�O���DA�T�l03H��BF�R���&��m�-�Է� n��'��S<���e�ہ�|&���,=|UTgS�!�F's��j$��`nZUC�������^�+�,��8:��K��9���Q��κVxe�*���K��j "�WJ�M���7�}6�5n�Pqw���Y�� �hu�M��*W?U��z�!v�<z�g��Ӽf�Ee�\Fꮢ�~[�R�R��mx�g��cs�������OT�j{Uu���W�#Cc>�����N��h���x����a$!����Aa��lZ�kd�. �r1��<���j�Q�nǗk���.֘,e��n۝��E9�
W4�Sz#	hOi��w�vP;���_0bY��3����@�*���E��Q�ɺ�̛�w׳�kvv3��wϳ�;�4��^�_��I�>,��4��(@F���9�>��]�u�$�Z_�,�:a�?�ߢ��Ɨ��&f�F��6�p琈'�J؁]�M3��9�>>RzB��w@��MA�`/�������f�x�y:����"U��z�^޿(��vD�=iE�=I^Q�`Ph����wV�*Nɺ�iw��-w�Cy�V���F�H��F�R
�qp�&��|�d<�eĈ�o��Uη�&�V��%6-�[g�f	�D8���L#lVR*�'�e{_R�z�摨���Q%��&T����������
���V�d�V(�"��U��H��Pԩy�jV�l���ZIf��c�,>I�4S�Zy�ڲ�����X;�(g`;�1]\�@��Bd�[�p�T1x��_���GXo�O:_�	��|Μ���ií��2��T�Azs���@���2)���5�C���6��u�1��$��ƻ;;�H/&�d��L��<��t	;���a�Չ�;�V�Gn̋���rl-�GW*G����z�B�o6�D��V�vUX���rǍ�sZ�D�
@d��trs��p��LU*� ���?�;v	�Z��Zb^�V���O}ޛ�H�AVÖ�A%�m��X�)뤝�~��&�_|c���fF3�׭���7����{O�aB	c�𸰟зs��	fNT�8��J!���<��{2]�&O�A��`Xw��9�Ӓ��b�Xw�[X��
&��4a7�� u�p���;�ܗ��C�r�UL9�7-&�!e��t���Kv�q���`�/u�hW�3�N���R���Z���X\^aS)�KG�qM"��aV�7����N.�|/�	%i�#�F�$�|^�b̐z��ڠ')�*��}�k>z��F��u��5�e`#�y��J���s_����KSl�*S�}u8�D�t3uS�`� (0�@���Wv�C՗�r�՞g�0��i�驔�;⚇�9���d��*��fw̡�l�N�B���U�?Y-�qǳm��j�@V��(�O��i�+�{�9וS���*��*ǡk}+W������g�MLe�����ԯ55;P��ȅ���UЊ99��,����Ҳ��K��圱����J�XL��+�J���K�<xY���"Do�q�V��U3I�Kq|�nK�ίG�ZV)k�؅�0�Z�w��]pcq�����oc]U�mg����+,��h���^�"|d��tD5�N��i�rH0῅x 8�#38	��VKSw-��U��V>3|8�c����4���1�����k�BQ^g@&�;�"x�P��(�_�tl�S��1�(x�+vf��:��V�,~�Nc{�M�[J�S��\m��P��4M���5���kS�?MdFHc�?����l,���3�?�>�b�U�E�ļ@ȓO�q�C+{��AJ��,*�P@rU��VJ��Ty���U�ܖ�H-�U�e�1���Hb���V�䢰�i�jVF[t֟�{L��$��ʂ̰U���>�%$�x		z��^ؑ��(')�������D�o����4W�=�e�L�/.�i�b�FM����p6� � ���367����l��=�#��M4��Nƥ�����GP�x5�:!�NU�1����]A5#�Dx��S�F����{o����h`�n�c5#r�V�]U��Ю�W��j��Cו���I|*	��Xkti}��������yo뙒������h��������u�?����j]*,��] ��Ϛbڸ���)���e��Xｲ�^�ğ��? ��q��Z>8���J����99x�*�BZqLw/���H�]�sJ�e��}Y��n>�� ���Kn������rϾ-�A/�d�޵�7�1�Pu��w��3�P2�Y;���v�=�t�l�e2�8>3t�|m��v�e۩T >d�=���)�9W�Ws��_�Qn��qy�4�.�rq���{2��SG�f��Bpp�vL���X) �����ob�/�t߷T�����������b���tM><�T���Ó��E�)����� ����?i��-k�e�P���Q�b�T�$dP�_�B�_]���C� �I�h*�w�K|Ip���c-SX�EH��<��P�?;UAs�Eݠ�<��YqM1)75�Gϒ��j6�b�I�2�z�:RS ��'��_�<4+�������7M�鳩v=�!�Ӻ3Խ�H&�=׉��
R-�Z��KL�q�X8z��t[����e��b��QU�"��44�r%�ܓ��]��)H��q��o�nY���^��6��LU!����ڽyam�g�uT�*^�w~$�m�7W.�7�ibbٮ��r��	���A�J�~;�AY4�C��B���8Ы5�3���!d����%w.���%Wb��<i�X������ǍOπ��4�VT�;uf��.Ȃegˀǉ���j`�ǻ� ��
�LY�D8���A�8�M������^���I�� ��-c�0�#MlC͒��x�;�Dsr4ٳ�,��ԇ�_�|`
lY⮳$*m!O�_��6"-H��F�E��{���b���(j��it�1�����Ę��1�K$�23�Y�5���2��t���'
C��dƚ\YW�|��#����E��:�=8�Uͪ9�7��&�M��o��n�z�x�Ĩ�C� �P�� GJ�����[� vG{�A��?��)K��𓩙/��xz�!2<8�K1~�IJ�����1������ob�C��G��q�
^�k^���R�%Ä���<9���<f��~e�4Z�I�hBB�&)l��:��\��\ƳϪ�����cF+n�,Mqh*�J �i�ð�'��)��@H���?�!���8��^C�����`y�)��;�qZlj @W��O�KH��5��d��l �+^���M���G/�k��zv�p���!6�<��[�wR	�%5^��?�w�������\_SO�����moI�>�w�7X?����T��X������k��M��И>*�=5\z����]���,(Zs�ՠ�z`ٍ�Z�ד�Jw�,��Q>�3�9�%Q�D���0W�ꅐD�]��b6�}�5�l��F�Q��&��lߋ�l���f�mlΔ�צ����4�754�%��g�{��=���{���|2_S��Q����c&����d���@0I��Щǽ^q��2�Pl�?kX�Y����h@&rS)����j�6-�l����=�#DO7��H�D�;�6���M^�A�f���ہ]vï#�'4x���.�J�h�{���M�3Q�䊀7�*�;��U&Lu�_�G�($���@M���V5�o�|��^a>�<�'�W��Bgi�]vw�Y�h@oYU� �Ր%�3��m��I�2Ԅ���|n���oO"�0}��D�e'�L�+�spjܜ������g�p���4n������w��O�L�ٕ�I�^����\i��� ��v���س6�_ˠpW��9,���3�.�	I���Z Ŭo7��4�a��]��Z/�8wj3�fe�䁥y�UF���z8������i/�MW8��x�?윱��s��>��F�r�S)�|�?\��n��۠J��T� ���� V�dSآ�>�4��c0orB��/�?m|7�Т�9h��6��n�g�摱��:��ezKǵ���r�7mډ��T�P���I�ӎ�֏S�#��m�1Am���߷��տ@9��'���x����ܝB&�D�L���m��/4�>̖a��[�+��A?�O��D��l��$�s��2�:g������^����Pj��3`ܫ8^AxLIH��C2�Ơ�drW��ƪ�>j�	����r���&iG��a�ٕ0�c�і�' U�#s�g]�;x+��lrzo��,�rǑ�D��L+ZG�����0��G5`>�E���T�T»��;K����=�_%��0@�� B+z�������<����b�x��Q~�1)�9I��F�`������cv$U�8�h�`y��ZF�ҿN����̞����/�4I��p ��.�/�����q�T���]��k�P	�y+�v�Ğt5��фTÜaͽ���CԏJ ��w�\�<^%a�-~/2��R�`��?A�K.t�nS���c��]h�G>*��H�L87�����#��.�&�󂴴�n�䶞�5Xi�^�s�L��h��^7��}h�u�ʂ�~�����j7���ڒ\�. 'ʖ�:9�R�-��FA�<�?g�f
D��[4��NG^����j��}�^��m��R��p�M[.�Ѧ�Z5��c�/�^`.�7���Thd�i���!j�.�!��#��d*��r���
�}{��(��sKb��ao��f�c�-Xa��/;y�o[�#_��x���P`O�Iw�8�*6����E�@�V��}�B��w�h���e�}�㚓fk��-�[g ��}�n�zk������P�=�s}6k���e���R"��zm�i�v�-�7��w�|��޺&�v��γϬn���N�ӂֈ"���b�wW�P�yBD�}g�rj�;@M�Z�}q���-���D���ق-�t�V���b�ji ����F0���AS+���Ps�\�ܙ���sB!G���hX�6(�nJ_��m�����2���\��rl���|�g��F���&�P_�*}�aqH�A�x��8Mx|�C��B����kf����
$��y>5Y�6�_�4���Jd��s�.5���I����˽�Ӧ��1P�Z��)}2��+�6�e�N6��2
@�틼�US8m�=z�j��g�Ȅ�g�
�܄���}��T��{�=M�}�s�PZ$z'a�].�+;Ġ�8f�t�h�Ĳ<P��P�B���-d��q�HČE����[�/Bʟ4����RI��������"�ϱ����ʆh��k�~ď���8{�;t�?���`����ݗ�hn�޺�B	?��^3Fj�Δ��^2�Y�Č�Ƭ#W����PX�P�Vf�O��:�cC��5��F3��m̞�F|^����̉K�}N�5�3���hΛ���0�Jqą�:i
:�9Jk�^�v�BQM�K�21.�(C�UX��û`(�{�h�v�u��ک�.�^5���D�I��Žl�AmE���aa��D��{��kY�T�SnpN�����7?�X���)ҝuH��h��f	R���)2�l����l�qp8�E��Y���_� g&�F9�j���|��P�vX���+z�k��N� �ֆ5�}|�\��`��'�����pby��8��Ďݎ�]�������r�o��.�|Xz�SٛP8�H+5����	Hl�= ��,���0P����n<��=L��n? @�h@��3�h 3�t��b�FAZ�Ӗ�����R�JO���=q�5����.�/5}#F}�W�
����O�%�e��4��T��%9��Dr%n��e/�zC����`����hwz�Ӣ���"!:ɺw�����'�{�y�/��-�/�4-vW#�,�4`�������~z�x|XD�zj�Z�v����H�Ǟ �q7�~�$G\�"(�M��:DR�|e��6�9i�o�ŗ.�i�3+'�a���󞌞o�7ߦ0$���wq���W>÷ƏU)m'p�\�ʬ:�J�/��J�P���Э�����p3f	��"���rO�'�G��\�=�V[���P	���������<��$F}�ӏ%T�V�@@���ũb�>_�{�^~�>s�Z���?e�_�Дtt	0S�) =��YEd$�B���3���$��]�o�
j={b��P7�k��V�!J'⃱�s���H|�����3hhT��b7t��p׮l�2�6>U��gr[������3$ݮ�"�iC���Ie(�ALj�:!.���VX�"3G1*�;l|�{,,�UΙ`~��۷#�; 0�K>�KN�S�l�L���r�XO*U�6�(2,o%���sk*��T�n�K�3���+��^����۫r˾�?م;@Ĝ�BK2|e('��P�s,ۭ<5�,tl(!��ߵNWr��ԕ��UL6jA"+����	y�?�80�w��ߑ����^mb��S�쩇L9^��0����=!�?�fk�������=��מ7z�ѐ���er�2��sI	{��G�Y����Ϩ���[G �� ��`�l2�ƈL`�b\��.8�r/�:Ъ~Ή_rC.C���c֦N��ڋj�$Y�(�:��৲�X���F�`�W����}۸U���8�@92TZ�7���Eɍ�o"*� �i��=N��jv�˲>];X��}Ӱݏ�ք[�/RrΠz����c%��uh�O��j�~�mL���/� ��9�����Y�S�7�&\l��h�ɟf���pSkKհӌ�Ky&ܓ�>�LZS6�u�Y��5�W,��l��n4��}���i�x~'ITԍѸ�0[z#�"XS�59��RȘ���-2U��
�+�k������a��	˭���s31���<P��[N�lp2!�a^�	즀S���_��MND/�3� ^fl;�%=u�&
y�@�ڔ�/�
��A�TB/��[ΡB�
�s4��K��,� �l]僑�ߺg[5�"͵��*l����O���7����GRd��C���J/�섂]�0��BW-K�NU'16��d���oˑ�����Fs��i�F}�` ��ɽ��h_��֍e=-�F����RnF �]{�1�5�[C�G:P��3�H�[`�8���t��b���J��B7�+�T/���ǁ��"~��:�����In�fFA߯S\/`2m��j�c���0�D���3�^��D�*6����x�x֝��-F-bh�o�+�~GKDM �;������v�d�
�Jzi0�ky�g�:{�	���4�#Sk���f�0c���
�FI����n��&ϏQ�72�����N�މ�(��j��9e	qE���ϒ�9�ϱ>O���Xq�o�8��*޵���Xɣ�[$2`:GͿ��&�^,6��V��x��Y��*ȍ_ϔ��?�OC��p�<�8�[�Sl��a�
�[Qvu�d\��r\ҷ+���عd��g! �C}+�0��(>�qfE�ITa�H��W��~�P+�����Wt���<�5g��uE��~�d���i��p����0���I�����h(vҮ��������2�/iC�J9��ee��+8OJ��w��T��E˚n�E���AO+4bk�V2_����Z�Ё�F�4������i�
�i� �X}ޛ{&�h�6�xBs�S:��+<��Q>��	�L�nXݦъ��˺"�e�')=�X@����7����)�$�|�uo���J�����f��Z�7��8�ʼ��n%�Q�47��} �8M�,nPlA��u�׋�`�\��Υ��Ya5G�ZI@e#�w��0��v,A��@e��J��+��*�֭-�Ú+=�`4� [�P�����Wa=�|�>��ێ���gh_v�~���o�B�.(�������.5���\�-��=*GqD��)Dx��`�z�;:�T�-��3<n6`���*`�ڭD�c���� �=�����(\�ʻ��a7�2�^ i�x�K�e/k���b�+����=7�}^��`���N��k/�{~x%%	�J>�H7�����3���K�:�2� =t揊�ɾ�Q�+и:��d�q2+��{j�f���Т��*���?��{-��a�fkH��VlDs�����PP�b���.N�,P��ê��q�P����R*�S!*�wē�)(�Q��?-荇ޠ~��8�4�;�X���	#��3B�l�H��5�)�q����֖l������7��*�������g�>	���D6MDZ��N-��D4˩��U�\
	��(A�Y�~A�7L���Q���}����c��\E{�S7�����������T�N03Ϭ�B�y4�Mӛ��Z͐�j����B�9t�8|�F����k)7)(]���l]�����"`&jDl��R�C��
�h(����V}�R�$�����[�3;/�yf�j�&2���A��
��M��L+���
����� $��	�d��W)v�gë��&�-J�Y-��SR���ֱb�f�W��o��6 �s�Pe�i��=��h��b������ZWi�%�o����穂�&�`�σ�8f݃RS�K�$Z9؝����_K�v	W�����GB�:�ux<�����tĵ���[����4'���^�w?ԕ�"@"�r��	�k�]���e�M��Ux����';C�̘�!��u�3���kK��ncy�"��g�2*��-�s~fK��
z��~"�Q)�EK��P�����njh�ٿ'��P6"��J�P�@�"	��|=��\��d\x2����R�KӹU�X�ɻo7�.:Q�\E��4��%������6�t����L�@l� �"+Nq��k�M�Hf��JI�z�CM�(KY��"��!��o��g�(q����ҋ����y��n�&bH$�HM/�O�{<��w��R�6�d=9f�@���r'��t�%����%%m�y)>?P1Md�O���:��Swo��xD�uvԓo���7�wl��4 ��N�"֜�!�GҮ�U�/�4�@v�����!��A�	����iF�nS9aʙ��)�����-�S�����G�Xlͻƴ���7� m %'}W;��Xv����pUu���(���5ׇ�?��Q��m�����e��W~ͼ�g��	}��7M\����½O}��e%=Q�� =%�:�NN:=g���)�Oȱ3�C֞D3�f�T�{�ħ�)0�GpRt
G{~.v�[8E@���[D�#���qD&�u�L�r���tI�4�����i��,>M���e{�t��W��I(����I%�#`)�[1T*4��fk5�TW2^o�����C��\�ҝ7�@W�b uk0ߺ7B^i���VM
�ȑv�Rl�x[��"�����b�ȴ��Ғ������Lâ��W9�q�j�S��x ^��^ϴ���7�w����l����eE:ndT�P�Q>S�^'�^ZE����������z7�U3�����
��[�,4��`�ToPRU�T6[��Q�5_�G���i��;Ұ�>�қ��襏R��X8HxP}Sb0�W�>$�Of���/`(*�e�O�� �W���R*I'K�"��+n"S��;�:b��80pjV�~���S�j)f���Z�K�l��s��h���A
rp^���k�i�۟A]r>0�()�J��=��d}:����6�(N������݋�u�\�(v�O��8����H�Z`���R n�3&b�Tw�سH��\1�j�!�G�й��������h9�nӽ�n%d�����RI6+IN��^�A剧�*�Wʎo.d��?F|�8sҋwE㓟o��q^���mrk�s� �h&q<@]l�ۚ{�`��Jk8 �C2uO���T.��_���I/=���-�W`$1���'���1N��D��B-UZ�EY��.�.�{��N��nb��Ϡ�k��������g��Z~B
� AX�ʶ�QI���w4����h�VbE~��u�+�~�8�%#��Ȫ,�~ z�)��?x薖�i{c��\ �~y�#[��¤{hP�O<��#ЌI���0�p��'�tWM�[����t�'q ����O��������xM!=�#���Q�wY@�X݀��l�<?�Դq����4���l��D�(qh�2��ރ��Y��vJF���Y+k�3f�+@
8���o���1a4��GVA���<�0�	�g4��J�[���nۄ���s=`+��1���dn���0�F��}���a���>�RC��0{���ۋ�/*_��tY_�"�� o�ӽ�~'�}��G�s�y1{��-�ò�>m��u�ɐ}2���yL�y\8�ڷ;H��i�tM|+2E�U���9)���RO�9��@��e����<��Z�Fa���C���Q���|�p��~�;�t��f�q��3���˒��
N@����3͵�7��3$�]N*Zhk<vl"~%�/s$;�\�r	j�f����I	[�����K=����yh��ϵr���H�Oŀ�lM�e�Ax�����6NW���5�(hgֹ5=�;�fjR�e��rRT�ǡ�����4�/�(���0,nl[i�?�2���(�G����w����i�u.6fF������cKw{K�V�ٯ&I�G�}�2�RB�,�Ud�Z�-s�p2�N�X��r�����@��y*g5�*����e9�,�K�ۅ�o�q!x��d�5<�M�g"�VN��uZ�������IorpKj�P�<Y���j��n��8Gc�s-���-n@l���O���R�4��9R������KQ�8f��tB��@([��;QBMz�o��x���/U���� �L��U�e����E2�N�0�S�_2�&��:_뫤n�;O��]&D�7�c�ozvR1� �j	9s✃��)Q�Bv��qr6]�;` !�4��y��N�c{�?-SGI��WV���E-�8R�v����T����/��8͕���\�(�JkV�FE�b~�-���X�V�oϜ\O������&z��,�̾#�S�!����g6E�&OI��ms�E�.G��no �� �ܟ������Ɲ�ہ0 8>����r*�{����b�4�D��de�@<��x�GQ|2�s�LK�+ ��)Ê�	��6��$�>02V�#��[z�:ntr]y�|
L �����a�x~�"
AP"��]Rj�MNC�.Z_���ќʏT%�4Sp~�G��:����+�-!\#�%�1���Vg��?����-��Q�b��Q}�$�zux��׸���}jW�!�����c�L����FJ������y1�c?&��w��S�>�.�����h�=KePE6�OfL��W$��f"g2�K9��+�m�[ކR�V�`����$YG	�-��2�Ҍ����T�7�����M�(%��S�����}mѠ���Qe�����o8K˰}7�#�lN����X��rF�$��4+�@orZ�l��5�ӷ4���赣ۯV:l+�]���o[WL�)�5oK�uPMp�����=6)L.�&h�xM��X�`��s٘~�N8��[�b*sF2���֎i�ۭ�0�g���zپ�LVE��s7�Y>�tg;22�p�A�L'���@iE;���<R��5��cj�<�Wy�6+�y���#RE��c�#���{��M_��K$So���;l��E��}�{���La�'ƌW�����
��U�ˑ�wT�@��2m�͖��Lp�g6�.��h*�����z���r	z���#�;�������_`��ZE�x?ЋR��D�s�������a��]U\������.�V�:P'*x�]�;��R�2i?S4َ��-r�5��*��ͻ�qHN�7�;��A�v{�o�� ��&O�D�Ż���o��EŝtPNfQT����R�6@��&	���	�ث�d�u���ԭa�a7g�~�h~��}YQ����(Z�[SJ���/�����N�SH#�
��=���i�jT���4��KlG��m�#��A�GaxYi�ж�N��A=ſsa��p��y]���dVA�V�b�A��_���9�NAK2���QI�1��$y�D6&�E��<,���AP����8��������r�$�	}�6�q�lN�=-�f�����I|�cz��Î��M���`wP<�)��Sh+c�;�.l �A!{Nd ���]�ɀfr��]�*��ގ�G}B=�p���_�����Xq�����Sj�#9J�|��r�ǮpUM�qw�[�!E����:{5�����N
1�jt&nT��E�Q`�`�@��a�z"���_���2�]�3�z����t�k�r��mSB*&��!%]� �6sPT ���7��v�P�Z[S�y�*��]{^.�x+I��K�ʁ��D�+b�Ñ�7l~�q�aK%C��%Yr�4m
�Z ��/���ίOC_˵5
=��6��L٩:�_���>��\2�wrHxW��L2fJ�H��+�u�3���L�f��6P�]����m<$��Ѵ��Y"����b�0W/�)4�l^Kۏ�a�хF_t�=��Jl�_�|Z`�ׇ /i$\�;���)�ؽ��j mg)�+���,�>|�Tr?kl��Ts�%4Ko�� .'�Y�}�H��>�U���]�'R�cWg�{`�p��_���"I�3.��l�m���[`�	j}��$�4���Xb7���:�꺳���W�6���6�Nل1�ӡ��9E;���.��8m�B���k�����٣t*�|oQ����o�t�������e���JF-<�mR���H��,*��ct���g�eg�5��6�|x2�N�H ���v_�v�ŧ�2a!�}��v4l}�|��Pu�)�ޅ0�ᱤ�t(��~?� ��m��'�+OI�u[#K˶a@� h���][��m�Y$?���xJQ�d�>o�J��<�����A2�����n�qOw.�3�H�����1�ΟI�P��)��j�V
 &�F����e��P?�2��c׿t�Q�gu�#�qt�å�s�����������/� ?�%��b��T���S�l�bnǍ	
�%�LVO���Sp����n�8�e-�*�L��m6���x�,�Ca5����|�-l
7��!YM�MRAˑ�����h����{�.� �+1����v��׏��\����[g`�z��)��?Zr�*
�=M�,����"ou^�"��	���A,[�w/j�"b)��$�������$���;M`PM�t)E�r�fK���LN����<:6���ﾽ�V��`��1q)v��r� ��P��o=��U��~�c�K.��/V��N�fȻH2k<7%`q��#D�%8O����F�-c�P<`/�����W�3܁U���=�z��|���Mi�Bz��p̽J��tjߟ����SV���<)L@��f6$���d��l���Ap:g�i��� ��A$�X�E���M�� .���tz��=���M�a�I�]�X�_.e��z�Mh<Af"�B��Bsd�N����;����=�>MZ����9p�S�3^3�kw"#�	?*�#/b��`�Z.N�噝Ra턃l����t��ƧS��8���	W�:T�N5	������1+*]����0�Jṋ(��K~8��$�"���)u�D�ՀK ���O|ԩ�>#��q�����*�G@m���-Ef�o|��t;4֗�NrH2s�z��p�!��e�����"�$XZ�.E�t,�{�B�G��~�N��p��jh�Լ��pZj/-ê�M���2݁����X�^����<�]/�wO͕tŌ�h4�@���Z�ns�����@�#���@�8������n���s���5�$�RP�}/���	�v'��.���QE��.^�,?�gB�D�UV��>���ٿw}_�*�JM�������C��5',MA����gCL��o�ra���h�6t��pd�F��N����m�H�&�f~\^l�q���d����S^f7��B���CZ�UU���K�u���h��(�R�v�zMݚ�������Q'�`�©"��H\K_��n8!�̈١67�!� C)vn��A~�p"{R��?W t]?��!߷�/�Ǭ�Xǁr�Xh/���+�q/+�l�:��	��ba<jbOr��LX��9c����4�h�K�(s�3�k}s���4����R��,�b2`���X�J�`<�2S���2�2U3�\6�Y��B�<�϶FO�]cn�Yu%�3������$1t"��:ve�beA@��H����ϑ���[O��?Ҧ�&��p���w�[TZْ�~���k�DQ�:�b������^�6����|�`~��}�\:��VZ��K�6��U�9���3Ԅp�2��)*��V�P�)�Э�{o]����^��XZ�'QMA��obr�?��m���&������y�KPc�q��X���,���T:j� @�|�Il\�~[Q�=�ԙ���������;6�2̋���y���h�l���sM�%n1'��.WB��XJy�,�V�r��fB]�eZ1��'��5>,���R	���K8/�P@��E4�C\	~t��"��PX��6�m*J�[m�?!�W��.e�q(�^VO��~��I��3��ĠK!�f܌$��.�KEa>$tz�%%^�߈|$�H��k�3��^`G��I�z�խI��Q
�okb�n��N3��"��N}'s����hq�W�A���le��G`����~��)����c�����h�1��)]u����!r\[���S��n8��j�V��nj�-��JZ
�.?�6���o'���{gu��O�!��iB���M��V#�����?״��^3�� �y����Տ�߂�6%�@�pmsZ-���|^"^U��
d8r}�L���ԝΈX��&�o"��8n}S����k2�S�����u^�|]Oڙ�c��W�Xڹv��jq��O�%�.��H-q�1�)���uW
X�����<q���U�Dub�7����Q�B+j��?d{=|j�Cy,ה%0@K�������?I��z�}�o�1�& Y�| 4��E� '���h��阫g>����i�������i���32~Y�����	z�|}\YoN[?���TO�?�Q؎󉡥1u"�����?H����
���m�ܐ�qA�C�y2_�5�p w����8	�Y�Bo����{���$�J�u���Y_�:���W�fa���WUǻf���<ؠ��H�9��>Ηa��.I1��r�E�W�I1������0�>*K�����\��w�>Fpީ���5��eF!	S��{�tk�`[�!��-ʣ���I��Sp6��7c�,�k>3bx,��J�|~�3ˌ$��R�p�s+��uX�ZE)C��i����3FWT�i�a]�!����#M�
�ѡ:<�u1�Z~��׌��<�-�MB�h�����_�	8e�39K?2�7"�pr�'���5��6u=����@g���vs��[��1 ���Yvꐀ�R,�#��W�<t�:ke��z��kv��	o����Z�1�7��Ӷ'���B��!����?R �1,�-Ɂ�����	�+M��tx�5GEzgu;7�ӟ�"�I���7М��=�9ߤ)�=fH;u�C���Pu��%u��ɌB�̠��'����u|�q��u	�a1#4�����\_W3w�!"�P͵9�@d5��{su�����*��7��-��˕{;<���Z6mFm6�̰��[�6[�pX�r�4U ����9h��}�P��HE�^����VН����9L��jd�R�+%���d\�P����&z�Or*eր6��LoD�Q �*f�?8�R�C>㊻�S��㈆�2Vϟ�L���L���'���9���Ɔ��E�ML#]��b�1�.+`��c��A�m��	ps���yH���V�`�R�F�{sg+���9|��{��Q-��g�C��\�(�.��D�w~�;�3<�hO�����������_�1���ӷ�!��×�/3`V����tdHb%��L�@��?&pQ���|�$7��\�oʣ+�l�0��~,�m�[���~�=2�!'OwE E=�Q4'}C�dO�i��"�eB�0��J����AW1ɾ�ԷS�@5��]�]_!����7!B�xyf�l�{ɪGڽ��)K���5~{e긓hw(T2�qd|tf��m�I����g����\."IqG�i��GiK�ƨ緿ob�����K���E�\�U��=�n�c0����p�c`g:>%��0�Q���/C��\ž	�m5�
�X�b��~8��&?E�����
�Tv���
8E���f�Y"W�A�e/�v�	#ڋ{��sɤ9�\�v��a��BF��㺢L|c�\O�; ������OY04�>7�6��ӛ�9��~R6v�͔sO�V�߈�����{:c'-c�~+נ��0p�=Hp���IT�M��U�8\adi�{���Di�O���#�x'�O6�;r��eFq�gx���標�a��3ٶ?`ʱ���|�oIgPo�S�*,"�cM2T��2��ħ�6�!���[PW7�����'֠5Fy�eҿ���Ф�z̔��u�t��z��m��&Gl���*��z��9m��V��L�p$L2lCч�k��{hݧlNk���)�
��L�R�ۈ��lwl�\�RP+���_��b=��.`�)����Y�*q%[���)���˵���YD>���H�ڮ���
b����*��:6T�lљ���G����p�(z���فyմ|�"�CFB'ɖf�j�[̭���
&b��B��N>@�ze8��}�@ʺ�?�ɣ�:�k���nY��Z_��L�r�!�w]ѳo؛2�[ƔQ����'>`���Qڷ���q�I�U@�Z���w����0�� 8�GFK��	`I��Y&?jFנ�uJI��*"8����T��}���M���0�i[p��0ϵ|	����s�B�f;$�����Z�I��z�/D�B��T?�Yɜ{"�O. �$CC�D���k�ӯ-_~h��&������������1�;��?�Y�z�P��
*�R��CGЀ��Y-�s��K��U6�4L�bm,�Pt���	I�\���i���|`�e�|P�E/���F���������2�P;���c�����A����]�3$�z55!t�Z��׍@j�>������tPo>AH�?���G�4�����<i:���z�YDA�h�\�o��ZnpJ�1�*T،-{��ʥ3����*�
��]�B��(� ���Ӱh��Z�h��+v:�@��y�v_K�w7*���Y:j�H���;�hEK�n�E��BȺR���a��藵�J�H��A�p�Ps�c���/�du��!V�6z@���t���AS���6ޡ��\�.�LDI�eAe���w.�>��-NBѳF"	�\�?U���K7����萢���������N���_�gv~������3��b~y5b��s�S�w���lSnu�x�1x�_��i=�}��3��X��$��r�{R<�{���@<!%�u(=��g���`�P��)�N���)&ypv��\��B����� 1|_���U�k��n\��ɩR��y��1ۦ�;.�"��k�x��5��S��yZ��e0	Y���s��>�<�G�(�o֣�m�I�nT�ڀ���Ծ�	rI�_���"��T�y&���O���W''b��K��O��W���dΛS3(D�N���Y7Y%�,{�y�����}�-�dw|����RɊo��#��c2v�v�+P�^o�%&�!�������LP,�i{��d�[X���5f1(T$]�Q��{g�>�R��L��x��6���m�=���+�E�9�Ѳ�o��b��ggP���V�
�fdH����pt�iTj��qVm����s�t%a˶�1�� s0�8u]�DB`s	>����ߵ$�lK0n��*�W�r|]>��)���t�,���m��N�-�����X ce�t^]�1S����Oa�����2�x�w�kr ����K��!��p��P��?��i�is}�ۏ�f��hR�/H�R'�i��X�T������e��)+i�Y��^�42v�4c9�L��������N�\ţ4ē)���+�����r�1�/�2��Nl��O��V��Ťb3�7����'�M'�wL��^ܤ{(@�c�����ޢۇ���U8#&�B[��ǂu�nLY�;�(S�ߖl�+�ïnU�&j*MV��_�~�G�0,�$acF!��x[B�$�_�>.*ݛc�v5I�UQ�^̊���N �/3�#`�~�H��cK-@8>�_L����[��g�_����-�,k� N	������Z9N��$���cZ⡷�'@^�N\��NdPBc닯��MJ�0�~_`Ε汮%�9�-͂�"�wX�"�]=L"���RU3��@���9αҐ��Q�)|0	0o��/�H_����ήi���5V@q
Q
�<�l�+���B�0�Ր�ᘀ�����ɽ����T���7wM2���f�,a_2�EX��0iL�y�H1s��g��|j��j���ͤ{�L%��fWm�A���'�LD�P<��2<ω���([�5��ߧBTU�Rm|��~����$x��빃��*2�*�ь;D�i�y��jL�W�Wa�D����s8�9�r}�.2M�I8N|6|Èx��Ӊ�h[g�%��\�B�GXލhf���	�a�$��>�k��^��5��HO��d�QF������"�sIq4�&�I���V���4���0�M���8�W��p����~|%�5��+�_qa"���q{]E� C]�=71�u-K�!������te?�S�&�?ΰ��D3`T�`��I�/������+#��{ȩ4�/m۬�$`mE.|�̝)Y��9g��n�I�ۙ� ���� ���*@շ��A�b��@�V���ED�@Ny��5�@���G~xRZ�����Y�]��~>����>�1�qJ���{{8��Vb��B�yI�J#N+����c�z��U�k)ƅ[�;��6���B�s;Tv��g���ĸ��2��l�|ж�R%���5K�:�o4�Ōf��~z�e�wj䁮�\���ʕzVތ��а�'R}�.oB��8o2����fӏg�mt�ƍY;�K����VB�J�.!���w4��ʜ�r´X�M��(YB���GsR"F����ff\H�={����9�"�����F��vuNz�u%���/���qYØK�i��;5��71�<l�U6�W:z'q7�.�%B8�c�7��B������z�R2xP$Η��s�:x��e~�#צ9q�O��N�m�M�@Րz�3l��а�JDD�����K/��Eˊ�C`��V/�ZF�[�;�O\q�?�����>�'�x5Ꮿ��N7=:����
�v��z�dIԤ!�TC������(�I�)@���l�����$�e���t���&P�/k�H-H.�? J���{�p���k��:�J�I����B�[�-����å����רL\�n쨥2rN�_�ᐸ�)�F��x�cA�"F���č��ߥAZ;�Z�&�2�)Kқj�`����|ys�:r�[z�P�7m��N�H�'�k�J�e�h��� E ��QV#�9�C/k���	4j`*3�e�|���LO^%]ߏ��U]���d,��ڦ��5ґ������vUt$x�,��ç��6��O��q<������|l}j��E�Nk������۩�嗭땪���	o~�K���uP��}�%o��O]�-�:n�,��c�Ps�0P�fh�MAb�VS�G��v�?ȋ��1k�I�5{uLq0��ݐ"��O��V��f.}V�h�+Q�����I���n��Y�tʼ����1�������B&
e,��>!���;�w�]����AҎ�f�,�ݸ	�VC=����ާ�Ԡ:�h�CwrpÁ�V!y*V��x�]Q�F��l_t�1:�z;�Yܯ�U: �@X\��y-�^�e]��9�Щ��T�T[#��w�+V�k�9��EB���rOU�ƛ�v��]����j2�^�צ���yfg������,����Ö dd����y�Ļ;ڗ1�N���_���{�7��ln�sXuF� KO�6��^	����W�������	�¡�.���ysQ�+	SaR�E?�!����O.*��G% ��R7J#��FHy������2��s f���R�yꦆ�em��QHN���S�Z�6��j��w����9*�|"\��I�T������<�OH�d<���<�?.��C�=,�p���iD����	�STz5�c��_ӷ��dĉ��Y�7W�[+�v�P,x��Yԇ����51~v���Rw���J[
�"W�]��kK��?�e�X��RNo�p>M�>A������*����mJ4�abƣ��lFm�:�ԁ�)�@�� Lw	��Uv���І���1H��#+���?����TL�Ǯ<%po�n1�ܯ��S|�zE�b���x0!ީH8�'y��Wr��Q`ҿ4dEd������"�IR懗��TҎ�p4�{�W�N�;4���)�X�}����T򶐱|����b�hS�#����x$�]fi��@�%��%5>N�j�x7ůB�aФm�8���oj�fU��h�^K����ͻ1�!�7����GMQ؇Y?r���'Ίz9TR�t�;9�"}�ɭ�WW�T'޺`$+c,�P�xe��7'B�t�)|���,��,�̋�����j a寂Z�P���:~�i2�W�L���}�b��0k4VL���������ּ�(1�Hn~��� ��K��Y`�����
�7�5�r4p4�9���9��C�44�+
s<M�8?��cy��J���g���Q�H���/�o�������EC ��|��.�w�u�#-#�/6E�Ϫ�}�6�끈h�,R�lw�������-���&��nZ� �5��i��UlŮ�Ӽ"d�H�u�db��1�R�cܤ�@�z�����QC%��	�$$�D|X��c�?[�L�8 V���o�Rc˴���֛%�K8�/������g��fy$T�"ȉ�|��=�R>�k�0{"� NA@��R_��3��~��@Um��@�ܵ6��z�t̹�f4�qw.D!l�ᣑ!VL�G�y�v;�G���,l�2St��J�=��q���G򝶘�dO�9�fVW�K�	�4�d'�q��%��'�����, t��eTuN�$�k�[+�O:�<��6 �t��ٶ�Cs�,�CP�����&k�PE���Fc5h���{}+�����`�����4�k�g���\XS󴮌<QDV��,=�# M��h7�:f]a29��IUP�n<��^y����0�fl����<?�
n�{MmL��r5�HK*�߂��y�M��_��i_ܐqOJU�,��8����+�n���?����f��9�vƲ��í�N�H���@��naH����A薎3���ԵK���J�m�i��1=x�ج���0��7��/#��Aˋ)J��r��w}�T���&yvU,`�ZD |���s�P2}�Ձ2U���?7'+��\=0 ��]��j��L��#5���bӲ�iO9Nu�����U1�, ܽ��HGY��g�呂tvu�t�e
�9}�.?D�q[do"�1�#�wu
�&�Y�����m��܃yԨ��X���[(�뭔00��m��ѵ��Q>���=��}׳����w^K���[ �q�si��4Y���{,E�'�F���ʸ�qEJ�vq�u6�eZፋB{w���W�Ny��� ��)�iu�a��3�����Q���ㅾ\%�$��Ź�*��:yA�j��h�=�5�����hE��_������
�[k=�S\��⢔L����M�8��D�#uʓ�pgO��#P���rA�Y��L���z��3�)ۻ-�G!!4Nxm���0�U����N]"�mc�,Q�*�s�Z�h��ӄX"f��D�)h�Xz��m�x'W�̭���S �usMέp�H�MmU�Q�+�^���)[F�$�Q �L�Z�1���\��i��M��a�c�����	:�j�����l�1^|����p��/�	S��Q� �h�G7�U+a-��]��&2:(�_Wp7/�1�`�S]b�O�zF�g!œ6j<� S��%�e�2EHM}�s|�!�\�"g4h�]�K�9׈�Io 3����]��u"K���)�/~�f=BA�
B�f;�u��B�	?�w���>���~���{BҎ	��3��^F'6�n�6���r�-���Yn�Ō�ﶿ��Y���輚�;�*��8.�[N�$	��������c�������]�X,�(�FY*�a�'gp %hJ�p$�4�1���zIj���yDP�T�2�����h��R2:�]�7t�=H�4�y���r��`o�*Ϻ�D�d:Z6�U|�7S�'�ɍO?�_f�X�gӈ���G}~z�
=�4�l�:\HBU�h\d��"ԭ3(���ũ@�v�Jx5��i��yߨ̙��1×�uY�  ��J�������F�;T�lہ�US##��3���s�ݝ�7����.�=<�� �7�.���5M:��x)����a�����,b��y�y��x��Cr,�tqP|zGd}-���H���f�0����?b�I �|l A�`��B�Gn��a��F)�ȝXz�|��O;�2T��]�{����x��r�}w%'=��� 56�Ik	�h��o��~����w�깤�����$i�? ?�L��_8�d��朿�����@��X�^��p%�)���/������h�0A	�vMl�6rc2�!6������	O��l�5��\#I?�>����X�E#����\�2��=鴯�EWsG�W��ZS"̼#�5��̼m8vT�=�-�U���@����NcA\Kyd�@�[؈��޼Q�;_������р�q��s�DTQ4I���h;@��8����y��:o������g�?���%VyǞ�dQ�����`����X BS�AO}e;�P��W���}�vҐ��q�@�'�e������<P ?~��P>d����$��ޜ9�#2�ܜy?�'����s�hT�d4&k����e��|�Z
�ؚ���x%�OB� (�.;:33�&H�Ԝ�&q5:�W�m��^�?�g��m[�d�c�<=�@��ǹ{c�ݴ��a���f.=O���L����$C��&w�Y2l���(RI�~����9X��88�p��T��J�i�\���Ѵ�l����hX��{Q��t�A;:�# S��J�+ȢV�-[.���/ T�پ�p/�J������hb/�t�<�Y7�۪J�:6'!����������X�4&��0�|�����T�����]��1��4b��]�(��Zc{j`����l�A��U�XY�[�:K����2�{W��M�m��	�,,�.�66:_iI�4y�*�p/��]9~l���>%)Q�rp�#�`��Āa㍠Ů�c�(x���s��Hh ��%���� ��DZ�P���WS��3.5���͢�yB◭^�f몔P;�.�;m�zb����C�JB0n+@���	@p%�����:�ݟMh����l�6�S5-eS)rE?9	� :8ǵ��Lٰ�Ò��a���&3��`�ÑΟ��FW3�bT/��:��j�=Q��9���1����w�*E���C�c��*�Xa���Zɑ&�[����]�i����c2��(Ʌ^�D��NK)�u}�	d�{.��
UA�tX�����8��|f~^��j�L��Ě�թ౗e�x���oH#x<a��z!Xk��8���w�9Y���sr��ݼ�2*�R�\�8��V��̭괗��̫ѱ�5ѧ�i��x��{s#���%c�-�����{*��[Y�
�TM�~C�&nQ�V`�G�|��3�Y�3i5�a尾3	�� �G658`���J��%�:��o<�j6����۬�f�(�î����������	��7u���.X׺?�@ߚ!1��ݨڞ���}��1ۑ�K�G�@�2�n���/��ǃ�]�S�mjU?�n��� ��2*H���vswKc8_��-Dfʮrǆ�lF��'C�g�'�a�yC��dm���t<�uW=�d;�xf;>a��i����ؓF���4�*�$������{}����q'6V5���sV#��7�l�t%�p�����͌����"���������+l�2�ic�����?��T�,�XN�(��M�BV�-�]f�ˋ,�b ���˹���l�V����������(�ʆ��ZP�,���IP���9���q�;�T�gɺd<�6��Y�q��"��X��:�	�:i$��b���hWO%�ȍڅ�k��,;�	�0��^��L)�U�}�y���X�k����Q����ya�*�k�_�9��c�3-�v��ϱ:F�U���Uy,1b6��׍l~#��z�#���l�m3�WW�JH�U�Y�T�"S1ƶV�&JR�`�:�y�:I/��`�1��BN�^��N�X��rL�J	#d�DX�ط����MГ)Q���OAN�Ϸ�y`}F���&~��J��W�G�>ZX��?�Y��J���I����r�L^�\�髉�{��^�ϓJ�V����.����N��T�NK^Pu̯W�o�꣉�?m{�b����!��ޟ;����e �9�B<�g:�) ���w�줜��88�Ɲ����Bt���"I���W�ҏG��L	)
����Hg��g=y��g� �ȏ(��1�����+�(��/P�k7��S?�7���|g;�5Y�����
�@��žљl��.���xHf���
���g-a�Ot-Suܬ�Ѽ����̠�G�Ԝ�/��٩��L��~-�*�n�����"�o ne���� �S����kۇ�r�'�W�o�n��J����Y�Ymy��o6���@IZ�)u{�W���Qt��f����dǁ�c}�+�.���F���MD<t��μ�Ĥh�*�sF�u�~�����m}�yX�S�+��v��*؞߸3��SfEZw�����T[D�k��9��Je��׏1�_��yxőA��D�J��#by��"�����%X�j���K�U�>�ٸ��g��54�w%!���d��n������Q.5����!�]��GMW��7f�%���ǀ������z�� "O������=CW�$�J�r x�`��};���c8���:a��Z/��p�FX1��d�=2A�zi��`'�[�vu��WP�;�و4�1��BY�QP�v�R���uDCE��>��0�W���vVUvMⒽ������?�Z���Y�j���[t� �<���4��0�=ֶԈ*�����oS��B:L�cO�$�1/.�D0K�����W�lk_���/n��"m�;�۠G"v���Rt�+������(k��bOy7�&1�pp��,|�] ���ɇTY(��g.<-R+��mj�����~����qmZ[]n�}�V|�ܪ���r�9��|rW���Ƹ��ES��z9㱉���T����wX:]���qپ��N������r�|O??��s��oz6����"mpq�~[�� �����̫&۫��՘!�D�웺��.�"F�v��I'}��z��k�4��Det �UN�w��p��:u(-��E�hA��K��6	/��A�(b� �N�%����PH7�$[����p~��ݙ������%�0�-QD�#BGs$����%6��p8�BR3�G� �C5\>`�a����d�fDVJ�z��,A;�p�S�o7�uaFw��{�yJFSL�K��ൃҢ/ߓ~�`Yb�jcM|�>+3J��1
���Z��CӉ�$  Q�A��,��F֟�Nx3:���6��F0���`v���f�CKc��EXp�F�L!)�-����.�D�8�ۗӯ2 ���
�������Clj�N}�%�\��,�z��p����ⴣ�9כ�8�X��CGX	-�J���Y`�����|6|�'�}�l5�!o�Ht*j��#�p����؃6���_;��t%�q`��֍{�\;z�z�	��??�`'
J��9���ѻ��o���O"
2�2WBR,��L��T]yL���uܠg-u��E)�Ng��1���m�?)�v:��W/@�X��	��X�{{?S:����X��}^Z�*�e������S�6���Wd1|�m ����dF�83y����k��V�3	�����c�V!���A�|���֭��AW	�õ����ep/[;�(�*V�6]t�B-�o������H!�%9�9�ODa�a��a�q�A���u�j��`gm�L ��>}P2+U�&q�U0�"�/�V�
���&n5<�Ø(�zs�rYo��&�M�-������r�\�R	�\��M����.F�ѷ3��j^_�b���I<������Mɳ%UF��Nk�B�Y�/
���Lӄ��uƑD�輻U-�Œ���)�1��|@>/��\�~����4��mj�	i^�B�Ռ&âg��aJK�{���ش��)V��G-��4H�l`B2�F+�SK�&yi���1*�8�2B =�Z�͸�!�C0�x��2ϧ�;a�����`�$A��}��|9l���#[�%��1J�� |$��؇��F�:�F��t�t�_F.���:�X���S��(��($��Nz�ǥ� �?��v\�jQ���w��'ε��%�AT�l��U
��)�;6 6��Y�Nǲ9��^���Ɠ���d��3��D�g�
+sx�+� �{@/�>������K�x�Q=��~�V��B�A������Q�\�>ܤt�Kd���'�T�8�\��Zj��t�"�)�����ؤ���4������p")y�f~@g���_�1UMP�P�Lf�f "�-\6���b����p��`:r��0`!����)���C�iM)�
�R�~�=�t�to>��s�����95�"��$z�7l���4�O���]�rڔe�~T�ã�}na¶��<�U�~��Cz��z�&�Ad4י�J����f�s=��#ܥ;+�g��n��DY�E���F�������tp��z�Ȗ�N�y���y�o�ڂ�iSV׉+����V��:�݁*�����5���B�F�: ������]�*���{��d&ru1�:I'�	��}C�,5�?'����|b�����]d��!�h׻�=A��3����pq�r���/�
��9[~^┊����X�cN�QJ���Xݑ�I��a�J���#�d����af�ƌ��E]����@^+h8����ccKL�����o�
Kp����20'�O)�ʲ����|��Ԫ��}^+���f(��!�j�w~�~�ml;�F1����T��8N��a���'�ͪB-����Vk1s�d�l��}�4q�7N����kzZ��&=�1��<P �>�ذh�-H�����![D��!YފKN�ek��fcǠ���V-�[�^ڼG�;�~e�<��jĹp��5&~J%p��%�^�
i����_�D��u��:�I.-��?�pX w��_���'��`�M��:�խ<���"Բ����>��'�<�=�-<�S��yMD�����#�\6��}Y�ن���.�7D���~z��;Y�QH�T�ٯ:b�XD����|ˋ�:�΂���ՏN;��{��~0�U8w��<��p��{U���b=�ӄߦO���ފb66Q������`���t�iAiw�����v[:#���$T�&#����m�Z;*�����.�_��c�ܗ����1�����FUD�D��_�]��|zQ���e��Έ�X�O��V�#��@?��7p�HC�H"�dg���&~r��O�Y{9����+3n�a��ۢj�v��e�g�����O}��_�<�lw��oV)�{�f���|;���d��)⌶�����j1,��^�.�P7`�I����MA"-�7�OdA��:L��[u�����{���wߤ<�s18_!e�@�S��~�&�Z��+.�3���Z�����v�a�Y�v�	t�9�D�V����rgKm�$4�!��h�w٪`mMD�0�z���o�&8�?x������Z0%��>{�r�up'#=�B�z���w�����ؠl� �콟-��⊣nz�O�\kY�K��MR4�|9Ä	��$�u#����]:h�^�)4������;z�&K�c�����/E����^H�b�����=3�G�y��d���pR-�X���9ei�pʃ�L�w���\�2�ꗡ����%U0�KK�,�b��E������˙�f�6��'X@V��H�$Ϛ�
��2�B#6ޑ�e�����ѝ�om��м�Y��x�:��yk�AmK�i�zf����Ͼy׬�B8( ��N�|:�.v%h����?����}!H�M)l<��=��6�16>������])�%q�!����~H/����r�lN`�1H=��e��GT�z�0~��K������R{���]N?��]��A�^�V0{�Q6;'�q�Z�m|N�|t�������㻷4~�e�]���s�+��G��%{����|�N�IfAv���1!1�|�p$bö�%�~�,�i�.��*���|z���{�< Fƞg�󶓽��Ƭ�d@3`@�$�g��/Q��;Z��!kU��*.��Z^�E���,au�%�B�Y�܅,\���(JT��S�9ƍ��B(�zr�(ȒYY�(KH���e���_�Q�I`I�S�t��U����<ȹ��f!��o�N�j+���6�p0�� �Ɓ	���m���T)��%�� �V3��`��:b�����T�ȱ�4��
��\jyl���� o�+�2��Ҙ�� �a�����x�+eBx��dG!��\@oͨS�ܲs�9��DP�;�@zf̓"5ʈ뻴c� �M�c"X���L�j~���N�NaW�� Jƶ����[���W0�u�LJ� ��� VLM�3�n���pM���15��#�c��uY�0>طW�8bK�"�����`���o �l@�۪��(�	U�{H��M�2��.�*n��`U��O����?4w���*u�Cy�w�/�zSp�\�
J�%��[
6� �aQ(VH��p�����W�>k��[R��H��p���}DH����o謐���uy06�������}`�$���#���i�;L��L?�
\�LX�6�F�0v2�u�6�p	r@,�Sm%���Qt&]���ym��E r�IQTa@D�#�x�q�Z�"	h2�f<�,��H�+d�輱z�G�n�p1X�����Λ�	�o���b�YnSч�-��b��^Q��P��r+��u���:��D��S�`_����o��D�Ēr��~�rV�Y�<��ka����F}��4K��z��N7�(D��8ط"3(�zӆnQ�6������Y����/�����[H�M���a
2�@.���Y�L𞂔�v��z�=�r�A��@ў���L݀���m��v��ֵ�irq���;�Y�A� ?
1���0�C�#D؉�S�P�'�(�N��l�40�L����0��4�Sƈ�꠺����׻t5P\qo�8�4M���5��vBf���x���@�8��\���K�1�%��ǹ�
�Ь5��qG>���x:��`���F��v�/탺���ҙ�nՄǈӱ2����V��j\A�"�Q7Q�_��S�l}E�۷�}��-��� �����%�G�Je���QA�����D���|�����Z����^:��\��[7��_W�^�E�5��ڃaR�N�t1!۽�3�$0����,kۣr�P��;8���+)���Ѡ;���G�F��n۰�L�@ϙ���д8��Nȗ��s*_�້i��(�.�Td%L�9��N��䪣�{|�J26����4��\�ͬQ6~�*�W�H0_���+��^a�E��[�le%�����I���$���,@��snd{k㬏^����PJ� ��L��?����ى~��r�4��;Q=������v�&)bA�{����Ξ-l#���5\���nԃ7���ۈu$�kH��n�����,GF��^sМE	����f����cBݏ��z�{�>?׎��B���C��R��L��:�Xr%���jU��>����F�k�����8�ں���t�Ԫ���y詈��e|5�;u���V,º��yV��:)!�L�/ۋ;����4G;�1a*�$���1\ghg���ۙ33�W�P�͘j��X���~kҕqf��;����P���2��%o�C5��
Od�K16K�Ti����ӵ��iJ﷽#�c�V�
��lh�3]���]�\!c�r,�����ͮBeA�hy줩��@��*5��� ���C��q�7�L0�.���-&�r^�|�����+2�l�K�Z�IRπG����ҟpJ�˴1�tFh�L1�	y#�a-԰��RK~�0�
��|G��8�C��&����5.m�Aʌrcm��b�+|�kɕj��=$�"��n��!1���i�?�ǎu��G��:���kMI����z���FE��%�hI'����y�N����/�
����3�G��Yp��%l��m���a9~Y?�\�����<3^���K���\�v�>~Y��F=#�S�L��!Z$pL���{uɵ�ė��;E�l�Ա�Q��B�$�( ��n��?r^�+���@h���D�!������F2$>�s���,��O�]�{��SA�^�=����&�m������R8��G��F~Uy�0L�k��KL�	��UU��m��?�>aZ�.�D���=mR9YY�L ' j�h$�������~�� �E��ӑw-�~"#��[qz��'���'�>}x�U�� M��'������t2��.��8��"|�fy�γ�$$���M�����?���hjf��X[�L[$as��
o]S0��"��j�Y+Zn%����������݂W�|ψ�+I��=�W+����7�$�]3�꫹�	N��'^&��B�%2a�6r��!�uS��N�@����♱: [��9���Fz9���&G	�߽��G����JD���[:�Uq)S��~
�_�XN�Gۋ�qU��a4n�h��HQ �۰<oq�Խ�nc����#h����e?�2��u��!U�պCI��x��܉���K�?*��\qi7�q��w<�9ͻO�jTL�����~�Vtq�ؽ�Q�� ��<�쮃3Uy����\��a�r}�&�d���8�6�r�QW{X��7����F�2�=:7��&&��`iȁ�zuǋ���M��@��qݕ)G�8��6G�U�A�lv�T2�@�>�3~�[ ��볠m��ip,q���IWV\n��V#�AA�G>����&<(�r���rF�k��k�
h#R��C��i������y�^�!��r��{�IM�[�'�e/c���U>|�:��h 8���i�()��f%a�����N�ś�2�O.�fge{\�z���²��ے����x�Q�5��:�{,A������y�����<���ǡ}�Y3b�@�w���X�i(��t[-��{*RF�؋ɥ�}�D�_'���j�j�޸�3m�R����4�0�Gl��q	�KsB1�� S����l���P�'��D���XP�ʀQu�� ������9�YLY)��:�_��]����
l��<�?���k���2�as/51T�g�D��N�L|�PC��I��0�mβѾlt�\� X�"2>���Σ$�T�Ӥp�������AjIg]h��x'��	6���꾤7�r�'�j�󼶦1���C�ol�$4 ���n�c��S�{|������f�R���;���@��ab���ㆽ��Z���Y����kՒ�\A�V��Ѐ���(�w�Ǟ����ǖ��hn�]g6�����$'�!���w?�f��]ѧG,fȤ���x��ڭ��ĒV���# 鎞
`�ї-K����=���3�ִe3uV5��I`'eZ�{x$r �T�J��:����+^8'�˯'���� �|�/_�4�8`���������LX�\� �M��k=\b$33�d���L��VMy�ѳ;�Q_]aM%���(�'���J�X$2�G�D��LI�+bf�s�cr��Uh6=/�Z̶�~Jt�Ǔ��t�U�ܺ������؅�N|m4��Me����%#���}�%�<]GU��r�$%���g�0(�Yj��ƥ�J֝_�KT��#=%�c~�"l�^�����6���`G��h�X�o��(���4Q(�)Pd
'a�y�9�$��FV��ꮜ������
H`] ʧ��S�2�jc������Uv���"�������}�����X�)]qX�x_�qZ�_$r��B2?�DL��߻<��$^/�N�����+�fLD?v�SH\�ܲ���\���G]CA�O�K��U���m�Z	]��ʕ���ф���4#l_FI���X�7BzDL�ܝ�	׳�X2xhy��œ���I8�vȕ[G��?��'y'nOc�8�B��PN��V�1�mng�#���r0��KBnev#�]vE�Ȉl@Q�1^�>����K:���1u�(���SϬ�	��[�I�f������B�S��=-ޘW�6��\�bL��xj6]��v��:.Ϡ����m��b��.�@
�6�T�{�r���-������l�!�M��h8�
�dJ!�?��$cj�$�s(&�V8�lA���2��E˛a��T�U�G��vE0�c�uL�$���#�F�n��A�?g�0�2���a��5����֎��Lh�YOF]��ZII�����IW+U��pʎ=�%
2���}i�)�0?�e�̳F٨i�x�3?�����Zh[���C��h���>O��/��''ɍ]7'�y�2Vla�+�\�1�؎�)�>����E�����6�K��#��s��� �*�n'�+.�����O�+Y��P�z�2�'�A ���S�\Z>�}HY��=�7Ӹvx��hv�i-%���?���L�B��* gNR�M��a����.e���"�"�B����%Cf�\�K{h>�Г-j$�e�鴵��UO�����Fa0��[+����#�GQɋ��+1��p�ٙ^ڙ�~A�H{��Y�x��4G�Uңr߻8���ca.z�ON�XxA��m��m��I�� /+�$���I���g�|a�|q#�Ӡ!U���))��=�H�Wu[�-�i�:�u����a�0�S\��W�l`�?ϽKו�[O�m�����C�_�"�Bt�J��r�v�Dk�s�?�N�"�&����RyU�Fٵ�e|
;�You���a4
��M���̱s1�Jߩe�%����}�}C���~k��Ԃ��F�}C� �р@�sق>�f��^�7���K��4����e�l��*B滶�spCNG@W�G)W-`G��tJ&��������{97�����4u�!Ƶ�U�8��=ļA�Z8�����v�)靲H����$�d���[��l{�J���(��˲)�I�?Y1��U�!E�IǱ녈�ӴU���"T����y,j~����;�nR��q@a�P�����HR e����=�o�[������n*��>�Ei ��\V�J� y������x5��1�@PWoB�gկ��y�#�-��)?.��c:E|��E���[���qAGEz�؎�YF>�硫�T�r=p�i�A�����y�c�*���U�'�<��"�$lZ�Xl��&��4�����f.�PX#�[U5"]�o�Af|��x f��wW�Y� o��ss|'`]'��== Ze�������[P�7�<���LӜ�}�ITFx��D<`�@����(�UO��?~�p�3��X��U�����ʹ���U�!�>;�Z�5C���7��R�5ެަs�1�o�τ������^ ����/�cA2Oߨ��	u�9�0�E�K�U k����#�[��>Lo��ʑ��,��0�?����fbְ�wR�^.�1���i]�����Jx��'�.�>��[}��~*����t:BjT�t� |�����W脉�?7�M�&7�G��"�<��}a�d?����Ɠ��'���E���Cⴚ�o�ˮ؜��ٻ���?[���������vG�fJ;��������s�N}��0)1).��.m��~G��-�n6l��C�h6�k�n��D�f���� �km����+����j�>�6�a�k��7��R�rI|���K�p���r�74��κ(��w������E��+>cqtH ܹ+���`�^w��hőP���Y0�f�N�m-2+P@�����dۢ��h�o~��k�����M%.Ǌ8�c�1)��}�;����]/?]���~���S�tIJ7HH����:��)����<9ж���9��D���F��5p���f䟳�'ߵ�[�ϖxԀ@���Ћ��|�8P	iv0��w󂠎ma����g��>Yv�9�q�zy�U�Dѯ�G�۶�y��4M��c�Q5�3�u;�Ouv�D*�-P�C�߭P	� G7B(Ғ�#�%�;-�<S�B0�J�9�v��D�zJޔJ���S^��*33n��O��񂠒YIS���ڕ���<m�P$NKbZ��FC4 ��=!~)!�%:8�<���8]�7~}~<4Ǧ��-^W[j��$����\_��l�<��	�F^�b�Ǖ��-ʪ^��1F�]����R:d2A_�쯘p��"2f�i���|ٸ A�<ZQQ����
S�.&�4Z9*UѢ�@u�[�=F�ZW��d�|i�^f�.6���hz W06�"~B�=���˔�r]�Ce.3�]��=�E���E�2;c�n�b�7[PuR%������q=��~l�.�H�c�d���H$��Ӂh~�V�˝nHCi�Z��B��]d�1�s����c)����뻛DSb��3���(|Jo��h�<�M�#��Ek��a�����	�J��LgQ��=<�����c���`�_&�yroN�04"���v�h�n9��K�?s�,M3SZ���]1N�H�8D���)��1���f�}���&���4V~�'v�4�Z�n�e����W�TR2wn@Z;`��ƚ��t�/��wc�H-���n�sL��R�e�a�KCQ������X��R�~Z�J����p�8���k4\��MZ�*��n�fT�Ϸ�u`k�M!zd����ʆ�?����>��y*��������l$�����#8?g;�n�#�>
6J-IJ��õg�N�!�gN�fS��X����ETꢥJ��d��G�
s���mHލ^��ND�,�z�wM�z4��v�}��s+��6�3�60Y:)5��/}!��Y9}$-����W�+��R�ҺJa�n*)����P2��i��BTѼE��stik�XQ�`Q-iX�3&�F�C�^I��5��t��Ħ�]+������Z��dSz�Y�V�б���b����x�pQq�X����R�]{Avt�5��+����	i�O�kCن�>�B�v�� ��l�W��ohT����O��D;ԥO�d����'z�u��a]��_ ��K�!�W�9o��+`<��_���	Ӱ�OڪL^\s$o��A�ž6*�1��p�9�M#
�ln
�Pr�r���&;���:�� LU:����2�D��R!}��h�N�E�.G<�ց'#��O��Nhg���S�:�`�6�t�q�������i]?�fg������q#��� ��}�Gd+V��a�Bp��?�lz�Ɔ+x_���2'�Wd��^�/�����n}E��zx*D�Z����l� ��.|!��G��%(�����8�����u�]��Z�x# /��k��qf���'q�T�ɏÏ�7\�\��@�������|ܺ<��ޝ+�C�b6{a�H�x$m��b-/&�[Zi*��ٗjV}+`�ʹă��d5<�,���F��۰��*�KA�j�6m��1�X��a�<j/�����d��j��+�TW�O:ιxay���?�1%�H���jK�c&���^�� *Ž9�T�Z��W�9�ۋ�d��V)�5X��*�l�AY�ki6��=YF��q
��U:U�(��6&�/�&EU�?�+ ��l\���}"������-&6�;M��ܣrf��x/���n�*Pbb�OĜ�)+��W��x�?�%������E��B��
	6��z���~[����a���+�yK3/����W˪�v�{ �m/(���蚢G��{��R���M�M��=wH+el�b�o�����$��כ�}�a��N1���e�Wb��:N$��PjA���3?��eXN{�R��򷔰�۵u�0��+�O �?nʳ8��2����J�-g� �����v{�~c�<)����;�^O�$fp�������?� �4�m���[I����^�T#:��蟃יJu�����Lt���q�d`L���)L^3rl��}��>p#�ݱG��UQa����:��	*(.�֕�G�X�%Om�p�=ZJ������_� y��?Z���1K�Y�{�h)�ZB�~X ��A͆����Lg\�����w�IQ4�`J���2
?����8߳����XC-V`H��U02��6�A<T%�H�~���߳P����E����䜰����E[��s�_���FM&���f��̯m�N�����v9`�')��ZT��o\��Ƭ�$�h	<!ґи�q���>�B��B�����e/�6��2�� ��w͙t������{@��/6kuMg�ʮ�>��� �a]�q��WGEV�����n-)����uI�zԚ�R�ȓ-�*�ɢG'"DXޣ U�Q"�RJi�<��]j��g��� r���nC{��z���I�|h�=�Ծ�O���oZ`�ǎ��Z�绌 �f�;��JU{�a\�t�3�Vv�oW�	>�i��Ye�d���J�w�M��x&`�����X�;�ll�����4�D����k6^���y�.���im:H|r�`~��9٭U���I\n��g�����a+�c�^4$d��ˣ�1���)2����P���d�u� fv��x��j�o�(<p�;'Е�N�I=��r⮗�3 ������B(�������V�L!j׈�>x���=@Sz����(�7�)Ʋz	v�	����3><>e�m��R�1�z��F�ʰ�)J�Et�66��!��3&Q}��~R���FR���R-�9�O,S�s��n�`5b�Pc˰�tK��s�9Xf��N-��_�Z~p�`}�l $��׌�?)�縅��ϟYc7q��7��/h�}�L&f���2��Z=��%I|5G���0�����}���V�.�[��O�U��$�؈�z�$#U(�'£���"�W��P�g��a�u���&����L�4��T�7�{�J�<�K �G:Y�M>@����,�y-�ߨ};�r*6e-��$�<�=��4��1羐�W�1&��%H�#�-�+�opOʷd���̓U�I(�ii<��C�����VT�q�Ծ��6��/n�\:�t�ßpw�)E��u`;A���fw5p;��u/�\2O󟪞#��ޡ����9�,S��g1��USc�7�X+4�����[9�����3y��{�iW� �Ltׁ�IB��UW̜��6�ן>�MT�FJ���t}d"�#���H������Dj�WRt����R��G@��pt��^��ۼ3�uԐ3�OAs^p�Y0*$w,\!�[)F)k� �r��h�o�DC�T=
���N,8WVa��s���fS�<��Sl�ư��u[3��ODIr���ǽ ��C�˺$�����(뙌��	��j ��=wNgbV��|.��'d&���K�e�����=T��0��l_�j�E��|H�3�E������4���Ԙ;i%%kx#l0�9��yUNa�ץ�Z@{٥���WɈ}��i��A٪)�E-��3�l�e+j��8�{�b��X�@B��W
��BI�ϲ2�{xg���)#���݆�7�����ҿy��3�Ie>��P7+�Ǽ�ȧK��R�4#�vp�M���+�) Kl�����}�2��|��O��|��,�@�.�g���.���������~s6����(	�f�@fz�*��|i�_6Q%	|k�l�Z��(޻g��8���9ț�R��㒇T������A]���aJ�HEf* R��-�X�)�ZE������a���`q_�{�>�f�>��"��ִ��̷��T�<*�?KȾ�ȯ�����p��D���̄H��l�)�.uF1�rG,��>�2fF����=	��o�õi)>�Qq�+�8�<Ñ�g.�w����`=`��h�D*=B!�9�銂�����T���ϐ����Za��s����P>�;�-�O�v/w&���X�|G�%2п�SeR�M�k��nX��7�z�.A� 2��W�6��WAR4<��ݯg'�+�vh�h4��f����ЪJΈrx8�N���t��}e:���{�/�$��e�8MDtXc͡	(� Q���ʸ;]�|K/eW��7���g�~�҄9�u%�S��h�yk�ʔ�)��T=��Ke]|�܂��+�����ՄܡR�@�Z�H'�̷����ȃ=P�pameJ����ɽ%���h�� �ߍ�tsD���>t~eWf����iь.��mv������-�SY����'BO�cʑV�Q�n�fBϖ�S���o"j�,: �Wy��۶���.ŧ�h�8X�'S.����`��7�����[�80:a�S)h�u@�/�k ��,U��˨��t��0�:=#�ɩ��Bp��\��j��QkY듔%�7��� ��R }ݤ�d;���]�!�L����%Ȫ���0KLh���J,�O���Q���\>8�j-�H]�V�[7*�}�Isk�O2�]M}�R�Smd3do�E5�ʜ���+���6qۮs����?{��A]F�"������E�CXH�\m� ���r�y_���偄T%�V�<�o�NFk�G:�'{x���ٯ�FZ>���=�50���_&)�ul-.���S�7𒥤c}��r��.@(���2���S���u=-e���Fn��q%S)� ��^���=��ĭ�C�5LǠ"^�n5�n���|��*z�4֐��/?',B/���a;zS`��l���2(��Y���35��"�����$yi�'C�$�ք��g�ډ�Q\n_�x�����{fDyl8~7� ��iL����-��J�1���E�����}e���(����uq� C���6e���w蜪"B����%��u>~���֏�#��?"H����,�d64I��i(&D��Z!��*��N�򙽸>A?����(תl�
􏟳jG��9B�GP��=>�H�ڣ��K�m�p��<�\�<{ݵ鞡M���6�^c�Q]��t����Zu90hu�;���?L��*�-�;66R�'��Jr���bq��̿���=�����u�s��OiZL���\��1�F������߄��V4<�'H�Տִ�?느��2pC�z��uV��n�d'C{|qd��vG�t~�As���_6��\"M��/w	��T#���E/U�a`�n��lS��ma����ɢ�1.���c�&)yd�})>!�R�� ��@�+���L(oKSm��wj'c��� -	J~V��bq��w4�A!�F!F��s�⽟�M�����J�i�U��ޣ1y��rH=p�qf�W��H@;���>�W�W4�4w�����/��zj0r=��R�{,��0��XcҮ�{��W�v8j���m噝���R��^U��U=vwa����K�,�P���i2�=�!���LI�E�قi��m����t#<$�d��ϐ����w�ܖ�ݱ�15eA�5��;���r�kjn��%�f��J�}J�/�5!^x9�W�Qd ,O�����ѡ�U\�F%�n�%S�6^�w����؈�&��%8��Y�����#���M��"�Pbl��߷>/��<rЍ�9$��b����R2�3O�e@�ϰ�o�Ns��OTi����
(�oZ ��y#-]��Sl�,G~����i���+b�@@�T.N ��=�lcE��|��-c6�y�����t�.�V�c>�(���#�%���W�N^+4^� 
Z�5wW����K���;�+p /��33�NT'	xG�`E�NS="Y���Z�(������MM ���.�qC6�ނ�tP�PV���+C�o������*7�W��͇iD�-c���J���f(�&W��yWfx�f��?}ά�6�FX�\�G�&1�[��;[������ƎS���x��b�+�����u��~r;B%vc�L��Cs3{d��_��پ���R]�$�P�ES�үg��1���)��~��-X/C*s���*g�(�#kp>�;x��dS�Ǖf<]1&p��.U=/~�x&��\���N}T��ۍ����C-n���'\V~,SB0h���-o0��4C?�X
"&�ך�|�%
X.z�n��:�W����}͈a�iS��^u�L�r'
��G�Cv5�ひ=p9�X�q��F<"��H��^,V3���
F�i�?5Y+@��i���<:��x.:4���45�y��+����ЯG��O�EҦ���e۪*��qB��I�c�&L	.�b�a^Ra5�z]�TYXrk��fNSGN��
���VN3����bayV%ۤ����E"� L&��Ʊ���=�\�W6Y�Y�7"����S��p&�Άz���g��X��{�J-��&����I�|�A��G�ոrL �.�P7w2Z�el~���9p\Y��^
��7�+OmU���VHD�>��L}��o��F��b�I�>Ϥ�q����&"B��ٙ+�Ѵ�b�d%.q5�����Sڟ��E}aݘ�7L
���NH�����GHN��0�l��u���qE�����'�;�FNx�*(�.�n(�
��E2ry�\r"�؊v����HX�������Q�,����/�|N����$��&u�x&2��?�&TrWi�v,�! U��+�΋oAt|�,W���:i+��Gsh[�S��<C'y@-�EQ�FƟ��W
]3��%�|��� ]A�é�k�j��-�x�{��u[��W��@kj�H�����C�Ԍ����c���ژ���upP^���>��@��f��1>͔yH���2{
�W�t	��%a-�%��ڿ*H�b���T���L��E�� 0J�.���=�qQ�tH����W̉r�}�QF6�t��b�!g\�����F�%� V0�٢q�	�ъ�b
1p����'�˥;R)��Yؒl���г�w~�Jt�{B��URx��>�'h�hh��1��ð+ ��%���X�95+�1zу=
?V���N�ԗ��[bƊKJ5����'88�hj�\A�J/���!�f�Œ��l\���'���>����i[�Ef���}����]�7F����%���A�V9��O�h=zE�E�*����<�{��N�m��t�Vi[��p
xI����tWVL��{��a�Gv�I��#�Y����΋M����Dc���
c6��3T�;D�W<n��=0S'l��u��K�nbh$c��݂S��v��LP�����U�;�#�{H&7�o�_y"� ���R�	��-��N/���N��z��`�v��r`���-�ʞ�)AZ���d:�*Vݮ�>%!��_zQ�K��	�1�"l8�? Ƽ�=�� ��+T%�[�%ClJ2���VP_����Qץ3>԰���'	��
��+������1MA�?�rs9�a��RA,�P#p�[ɣ����6�,��uՐ���J�LOo`�Ѩ���
u<(��֫��
�E�"]��*�S�G��[%�4��=�;Pa�L��/9�#��R^Y�˅$�~�	@N�Ob���aw�e8R�r��ĕ�_������]��9�]]��{;`3��a�
��x#JJ�������D]}:x�����u.���"r�幢T��%��
���0;���j �D�~,�m-L��q���c������3���[�g�K2�����.��H���J;CH�r5�MV���@��U��#������J��������'l#�� \���!Ș�Ln�6 �����2K�វOML�>~�oZU��W/�[qHo��:7E�~A�^bd�!�g����8E��'?��a��[���tƊj�5A�#1�E�|/�2u�>~��]�Ȫ��7�M_��A���
��}��C����Gm����?Vf��M��8��W�й��&k�n(SvG_Ad��P9��m>5�ʒ5�|����n7�9$�YR��89��FP��􁾓��rf�ܛQ�r���=��\�(�hk���hFSp�m Z������ؚ�9���Z{�d/��[#�{*Ŀl�=[�i,7e7��l	}	�V��-2&� ġlBB_�"w>�d���(O��V�۳O������ӱ����:�4���L{��!�r��^��x��!j*�|�9P������f�[��e�Kڥ<0'��f�Z:�&}}�QB�~we?�(�-��`Fl��|c���6���G��v����q�[�G�PL�꫎Ĳ�M7�y��N8nP6^)�x�ɜ��b�L��a������:��}su` ���m2|6��Pm���٧�X�=����r��E��������
��Y�����R��8T́K�_Zc�l$ޠ÷\(V�[6���I����[!C��sp�Y��n"O|�A����<KI�]��~��%i��٘��Ӡ�#����#���D�paڳ�I�z�G�1
̎��m7�5�AjY�������A%�=&K%��y��j�7 \З�g��P0Z~���TC���j�7E��ndv�B�� c�_�*�1{�D�>
c����GdyYV��w��)�w�Y��?�'�~8"���E���h��DjWUN;�a!���K�8_ь�S8xwE��I�C�����GA�B0E�Ų��\B�Y���h�Oog������H?���ɢ�6��E��]����UJ�a��f.v�̆ D�ƢVo^�{�B���!>��ڔ�Ju��:��ٻ%�(�qg�E)�����;S�'��J �:�C���-�&�4"6lS]`̗�&�sT��i4�D�RF��]���n�#x��ٍ����&[x-�ZT�,n�]�<����i�~jk��+P�D�!����-�L>Bf܀p�uZ�4��]�e���;��|q�阪�n�ć���>XZ�|��`�6�W?y�G�s�7#�� �F"HoN�A����|?�tʯ�?r(_�>�r�Xp������!kŘi�G�0e�j\�a~hth1b?h@a����G�>,k,O<}��kY��U�T�ms�`E������W��<ZI���NKאa$�.N�����L�{��y8���`kA�粙k4^E�6>芐3c�E�g��89� H7Z>E���e��G�r*[�}��U�fJ>�������'�p�s����8V��g�	z�S<����+�a\����?��}���}~zО��R�5f�q_����K�N&�u��&�^�L`[�:�n���K�+��Y2w4|�% ��Cd
����n�������z&���doI�'�E���i�/����0A?!�����]������ �����p���J�������_�J1=L��í��e��(�������"�
;_�\����\�a��*7�i���]b�(K�(x�H�t�#���m��u��֧�8�*��~�p�Q�����A)�]�=��FV��n�"뢿�9��沅<�l24[�F>�O ��(�����ޱ�J��n�F���q�&��w��T�|���t0\�t3�u����H��?�#��)PrC�4��~A�W���R��9J�����4��K=��䔥E�^Fr����Y�D��r5�b��*Y��bq�"�	Y�P��,���	�Tlhi�gJ;	�rr3����p	�=Ě���|��Hq��F�w	��y2�8�g���c���.X?��[�����:vRڦ,A�R���׾]�/=��i��M��z�C��s[k��W���]NԽ�I�����x�f�7��͆�	�u���Sq�"�7���&6���� D���ogCl�� �!�-LP�j�x_[O���Y�/{�����Yܖ�05һ�_xt�$�҈;B�Hj$�{Y�&��/�!���m24�!ZHJ}t�:���@Po��V��@h?ٛ�YZ�zEx׺�K/�>[rr��Y
�F���g筓 %=JMЩ�標b��e�sbh�fͶ�O���	� �����>J�����&E��d3�`߭j�&��A +ɰeW��U챋�	=+&���v�Q�i>��t���|��ި�տ���"���3q�z��q �w`%�~2�T.��!Y�7~�CU�ޒ���7���ţR�1sA5�\��+��i<ᛑ�q��~Ny��)�j;�F�A�>{*D`��A�r�z{Z����]��y�C�~�``��� iv�h�管�2bQ]t����Z���bq���-z������~͂db�]��r���{qs��~�2�8�L�9����n�a�is�>ץNv�Ze�����X�d��~ς��L�4���?���/�.C+��]�&�Xu�p��Vb?FpP���C>�D��e�suk} ���� @�m'5[���m#"�����J�ׂR�Uq���|	��S�g���߈@X%."��!��W&c#�b�I1�p�����  �ÂH�E�4�!�N�iI�5"xx{��w��I��
�E��^�w6����T���%\b��M��
J�\�\�x?<CI�	6kL���T,l���L/Oh�,U�;܆6�OR�����a~xP�����*3���FO-`DU�5�oֶ��zaPE��uq}ɜ6�{��v.�{��X7�Hw�"��"�؀14(��L��)!���#IS�w�V���t�z��}k����O\���7��<��@qv����A���-xn<�CR��gtI��T�P+ķ�j�T��1GHg���C�#o�����?ϓg�95��+@ң[^-\�8�~��#؟��K�
bE*̇&�6��./_�CB���IM(H�C^հw��/��Щ��i'�<9�2�����w����m�T�ˌ�
�L�gi�d�̜�P���lٝ�/�H��F��2���р<z��d�zD63��a����'�%[}]���cЍ��X�%��>����J�ró�ڨgr��p��,v����@g+�G.���療tO��
���f�x���.�XG�j�¸@=��2O�����!>�H\�o�����(�R��7��EW�̇�T�=l?��Fp1��g��J$X-^z�
�����Q���C1w�)i �H�������	a1��r��.� ����5��c����8�������$�2�E�Y����^�m�����)s,xȤGh��Й)�F`(��r�,4�Q �E���J�E�sJ�z���1�t�	��u���#�܆�5�FGx��V#+~dS��b�N�	��ϩ�m��FD(U!D�&^OL�bsr�����-F,r�G�$�^�uI�z�+ٟ�{,Jr��>�*����0y��؝�1L;�^B���Z�(�W��]X�/��<u���D����<NpaL�u�p6q�R���Cǒcz$�C�ui���8��q�|���u��{�f֮���V���_�a��A�7�S���l^�լ���ù�|���4�B���(������L�W/:�@���/t��;�����Vep��L/{f��qBo�U�����<z��ظ����bOT�f+��pb�.wZi�(���u&���}�Nq/�PA�?�6l��(+�Ys����,}�+�)��r�k�����h)�mD��UQ��I�=a�Ѯ� 쳏�)/e���,�́#��5~_�cԢ"k�ۇ���ZYg]��}Pg�^���w]Q�(�12D�Ց2�X�4�b�WM�||{�#F0�:�(���]��O�a�ڹ�G������>,Bƨ���;�0'�<���J+9zAY�c�� 6�iC�!���C<#iw}�P_��%�Y��r$bD��Ifvun*�x�Nq������3�}ŭ��_�YCǍ�{�3�Z&ˌuGR�̀l�&D+� N.��=����ZVD��=[TC��˅��GTM3B��������ˁ�Q����+��<�t��A�G�jj9�c*'��D�dt�`$�o�H�����K�KV�U;�ч�3�D\^ϔOX��s�*��[a7��6�4�V)�!�9�{�CWu�g�;�Qw,HR$C��L�5�RgǦQ�'��ɣ1�$t �OA ���^���q�,�[#;_�S�~���b}A+6���.	k�̅����k��8EAR�>��U�-�r����>%��i�����m�2�
�de-$-��
��q����1�ē��J�����D�d�Z�����%+���X�ӡ�j���H5:p�5
C�%f�h�1_�}c��G��J�a糹�C�@�!$o�g�F�\�%@H⪖CG�$��C ���l�k�#D3SF�}��=a��,�I�I�Yn.������F��OU���PD~E#���ֳe�\ә\�����|���� ؼ��8�o�W�륡����X�b��_q�����z�/��(���O�XT�M��=	(ȡ�T�3�e��*?��y�)ΌwZ3�ڰq �R&U��qB?�Ӄ?�0$�z�h�|v�K�Ӓ\� /���(�z`�,�Q�6�7�����4����N���i|ә���C��X� }k�]�l�ط��v��͊��s\F��,�0�Cd9R0�&�ݦ}}:,���>�s4n�i���eD�a�Jy�N2t�=i$+ya*y��x����BcGR��KT`�H�u"^]A�������x��K�THK!��h�7�4\5������R��2$�3#9e�z�5�4���2I����NIρ�|ӝ��?�z>�<�v�@��^B��H���7��I�������8,A]��Oϯ�[Q��6aew��󷙔
ȱ�J�Ione�t�n�6p�ҽS&UB��K#� x��E��R
ݷ��/�����|�܅��m�f�Q�¾|l��f�w�>��U���zz|��(�n�J������T\�i+�=9E�fV�+m⫶gkMo�qc#��������n��3DF�Q���-��{=S��:+���#{uU�E�Eғ��B�w)v��w�s�o�u-u�~�u9��6haOU�X��zq;z�wË�|��A2�W�pJ����Z�_F��C��2����_kvܜL�PfŪ�������V�?JX8��ԓ�l���a���8���Б��n��1�]h�^a��� t͞\�O\�	��I��å��0�Q�s5{K��īZ�Ai�oK���0�0,�t�	�2�<��5T��w�~	��}5c����M�`_��)�`��(������*����NꕆM��_��·�H���8�C{	�+z����C^i�;�����=2V��IHv�؃�n�<`kJ��wʜ���z	�G�乕��7k���J�]�i�����+ے����TRۖ�7�U��{ �m�Li�q%p-�1v��VJ�ת�F�FFMb�c 3���s}�P��K���~��9h�Su��-�~c_����o������L�@]�q��-_��gNrQ�����QI�nZ�	�?��s����[؟j�n�L� '�ŉS�"��M��{���&	��N_=�-np��v(^v�'uG��6�>|��Ǜ��kg��T��9��A��?���3�+�<D�&?	.�������A���<q���mPRL�R�����!�0Y��6��*Q2��`WBتD@VI*m(y��>������>OH��H�Bʧ�a]ߥ��MJEs�#tǩ=�������Q\��#����#�G�!u�1�0�b`\�&�X_�O�(E׌��[����
*O����"S�{{/5��Ş����Ve=��w��_!"���[嵪ٲDV�
ўxc��\wM�߽νC�v��Ы� k�0��{���%��OSO2��E���RE �+���=2q���Kn�A��R�p�R�%�-3���5軮�9��k�����O
���5�#AP��P��=|n[N�#fZ����>��[�R�PU8�lje\�ewX�M�ht��j�q�9g�C)8�W��e�X��;*L���ۋ��|�� d1�T�0����OΟf��d��*�M�������x�P��c��[�x�7$k���}��*?V�k�pR�#���;dk:�Ik:[����E�\ЀT2q�}`�e�g2�π��j��"�	gJ�\��Ó��H�p,�������fo�i�Vf�!^���.:/]�-�ʅ$~�������?�@�@fUm� �æ/�U�C�|�i��>������ׂל��h6�Z|�K.|X��?�\�.���oD0�=+exUv�y��n�0�a&�pT���Ǹ$*�)g�}i�;��v�RoGs�������E ����g�&�������G_�.dư�]���	T�6�(��V�7���_��_���>,�Jr������%����Fw����W�?���7���W�����-M�~o�#�*adOM��g�2��|Z�T�Ϲ�)X,������3Y�p"�8u5P������|6ܬRYD��������+���D��m�XaQ�}~7����B���P������8��@��u�,�o�B���\�݂�0c�i�@��\SY��>���J����6@�V�2\f���}I����pz'X����"]�XLuR��%,)@�ȓTF#��m"��,��:��P�SG���$i�:����X�^}���I��7�l��$6��!8��3+�TQ���d_&���,E9?��W��xF�G(�r~(�slI�{�GRH���ν"O隘l(�d	U	O(~l���&_g�[1d�\rf�C���L�У�e�A���&qJ� �����:�5�W�Hx�� Gz
�Rac�Q�	b��<��7�Bd�_�x�`���a�RD�q�����u0�(G��-�o�ٛF��6��^����k�ѡ��fZM���_�¹ތ�~~������NBm7���������R���W �9��6-谱3�3���肳/�D��K��q�Iy����[1�������7#���ݤ�5�[�� �n+�ӂ���CJ�N���tՉC�}�]}�O�^��>8�q�XR���N|�Z�h�ݻ�?��ͣ�s�Y�Z�7�����n\9��@��fr�����9a�rҠÌ7M� )팆sc��
F�N ���lH��%����#>���~���ҳIz�_Y��}k�LE�2Yy����� �ɷP���I� �l��
j����R�Ą����
���Zˠ(���-)��!b$ӆ�V�f�Ea1|d�>��S�@����7�b�F��.x�]{�;����f��6����}�.�k��V�������6����nN�f�4uc�������N����f�vP���zT���j�Ixe���F�$(���Ƚ]�����:��+�J-�w�m�˥�-?��o=��IPP����`T:�.�BG�51�,W�ר����%N��0�����_2�6t-�� ��0���@��󀺗	�+��ut���(l�P��	�w��A������I�,���% ���`C��LD+�9:m��1ֈ��ѺO߅+0�"n [�9`������Xk������gS��!R^vak��-��ݦ(�N/"ӗ0�P5��<�֓C��'�>�N0�m�?d|:�ksB����wI�hR�����K��E��L���2��a_��;qtV�@Km`�CA�Ȕ]Ğ�cj��=���U��v��>nH������x��.��;ᶀ8PL8��kf�q�y}cٵ�3�Q��G��c 3�!J+�q����CpN�ŝLy6aC\�w�U������%H<�S,][#n@G�qw�w��=�^���x5���=��C�O�臻4�6��"�&]�q��}��YZنX^��a�I��
X��xTch0�+T��� �~%�(6��ނA4���h���K���9Գg�r���RCT;z:�Z�3""��0�ܺ0���N�o��򃍦�����V�=ru+��M.:�y��鮿G"+ �@��a�c˺5q�_����h�D�鉸�BH�s24�F2B�:�֮� ��i+f��}�B��t�Z�d0&-��=��Ο����Ɓr���tc���%����U:x�E�?�z>�T6��]�\��$�D;���J �។<d�Ux�<,*Id�jXϛ �j���mD	��F�=�h˘�Cƍ5��Y9w,ڪ���~bC���KE�l�ʅT�q�nÛFgW9�VZ��k��G�u������9j���`�#��g�[��H�$,�+:м4���!���]�D�ӹC���n&�WT��Z���\��31;�"�-��z��Ǻա��i;��TW��+��M{P������~i��AJ��J�f>�-��Sz�� ��P���#�"]*ܱP�;�/x~P:�E�z��L(�x8�
ƢV��R�|��W�Rgt͡�b��
��PKTx�,n�%is���9�c!�w�zC0.z�>��S:\���n"�/�6rMo�L�ͅ4$K!8W
p���ͽ(g���G��q�$RD,������`�3Et�[z����9�ӻ���}�w�vUM$�h7+�@��`A@@5p��w�{x�/ԑ�0JȖ�������2��e�خ@1�l�(K��5�s���󲷜z�K�ⷯ����q)��/ƣF��P��N�R,9 ��ʴ�>�����i������7�\W��c�'G'��P�n��T�GQ�3�����L�n���x�zMu�ˑ���z�1}����65����|�y��Q��
��^�z�]�Þ��h,;Ԋ3�&.�3#��x��|Z�U;wr�~�5�.N�8��g�+�@D�oC��	6?��v�Ѭޅ�uy��G�xMC�69�%%8*
����S��=��M:ֈM湏��+*��%:���u�Rm28�6�`/�ٚ=���|5�-˒׽�S(t에���55�G�h�&���#�VX�ц9�|2x��Ԏ\O씸���4&�Αi��])�mS���R�_�6/���n�
��u������|��:������M�l@�H8�]D��L.u��G�Z���HM	y����Nf����P5d�6���6�N�H?�_+�qyg�������Mh���ϬR�-`^�&�@A7�y�4��~�5��B�sQ���c$�~K�����'D Z�ZqqO�ɡ����`&R�U��:�B�E�:��i��0�ɸ���#�l=v�~\D����	�:
�WH�e�S|)�@�/?��}��WR��%���*�VIHm�
<�W$�a�-"Ԙ�޼�6\�;��3|;�(Ԯ������8�-�|�}���s��>Ϧ���,m[����S@�q\�>"��%C��}�r�C}˙�2N���lVF,N��'��^���XM�9����r���q�g
�@�SӖ��;��p���Zx�4`�B�=V�t,s��EO��&ǧ�3��>�3�P�RDv�Z�M^��Wx�C+)�p$}��F9	V�Ad��~u�}�|/����]�!�+n ,�8�7SV�r���0T�/��V*~+���#&k��_�����yb�
�3v֜�#4Ͳl;�2׶�r��h>��lf::g��'���]ArgL	7�)��êu΍�^Ըm3C6q�~�լz>{�����^	ٕw�J.���u]����l�b�p�n�:�k"ԏ�����,�L��zS���T^�1�5nms����yY~ ����D��Y� Sf"C���ٻ�	��fUaUȦ���r���3�..�1���s���ϵ&b�����F	�h�U\�uV ��r�.J�f�U� � U7�#��8I�\�jWQ(� �j�H��d��YF��a��[�"{Y���j����{���<]��h*�?�����]�T<U�+�_S��D�L iS&�������� ��c"��f��q�]���{�Eq�*�v��1Fk$���U����X�G�U�^�4�N�AN�����̃�N�2s�R8�*v�Ş�%�E�܍��I2R_���T�ylx��c�H�����w�X{ܧ��U���B��G1���g�]Z��.�XlC��u�a\�;\KdX�]���fhl0X���7���>��b>d*�C#��ںc��_��Y�)W�,E���V�[�*���/Ts�g h����X�1�˿�m����t���I�(�9LA3�އ��x� ��|�)�PI��M>��ѯ4F(��\����W�w��h�v��� �ʀ*V����W ��N\9hO�7eVlc�]�f���� ��H�������uN��P�1i7�g�Q���q �o~�D�~�;�Tky�;�d"o.����zu7BX�q x٢���ǲ�=u��]o��qPsN�/��[}dtc�{�+`�D�JS[(�׭'�.#�w<�4�?�3v.�n��E4�FGԲ݋_{�^��ώy�f�|{;<6�S9l�ks��2�aFN|�,�R<�r���l*�XMNe�ܞy�:?�,͠v��a��i���M_|�����c/���Y=����R#����b��/$�����p����JX�i?�!�BGO�lm�������f7�(�]�� �q�U%{GZ��ǀ��n�RST��+䅑A利���K�zo������=�z�rXC��8��_���_V��3��a��zjOb�M����&j;"ѝ�q^"� Q:�C�P��}�})��|��r���$əd)����}ԥp�;v�.n����`'��${�I֥tP��*�]EV|!��Z���4#W����c�eG�UX"w�S2GcaCyI��)Q#��&:�q!�ń6�a��J�ڲ~���+X.�)��
�U��<BLU��y`:EQ(�Wr�ggZ�Aw��jX�"-��Ѕ�� EJ�bz�^����c3hŬ�dN� o���;Z^���.i^�{�]F~�JE>�r����QKl2������G��d-Q���D��p�F&;�$��J�zۈPM�d��"��C���D�g{�sz���i��$�з��V"�7Z�k��-�l?}D�E䂱��� uV�!ж<����L2iPPn��|�P�E2�\�=�ZZ1�|<�q�B�1i:��GWF�e��!�X�<��7�1��X�cU�|e���W�|H��q���T���Ɖ�S]��N�^P��q���o��Y�����H�|��)ւjބ'8�ZY��H}��`�w��$+Z}�B�<�7�D|%�.Hotb�����9���أZ`c�l�ͼ���.�.�`�������wT_oq�۳��\��:��T��[5���A˧�Ң�X�[��:�V���8��8��.k�B�N�
g�lBb��@��]]�Ѱ���Q���Ѐ���}�3�H����}f5.��!(^�� Eʹ�zݕ���u步0�Y���Wo�D��jU�{�az��c�� ��/�n��'Y�$�F�(E��fV͚�=��aH<SO�^�`�C�����G����9�>��
�K�6�3]=0HW\�(`�c2��b>c�XG�=ԣ��o�i�9]�}�)z����\NN�0?5��-U	ߏ%�� �?�p�Y�t�w�(2sg��<#kC�]�Ak���3����!�1���cT%��_���P�K����ġ�YM���>�q3H��V'�YT�z����
�*�賸���������ɱ�A3!�Z}�/Q������J~%�|g�$�^I;'����Wu�/�U������@x8�:xp��6�h?���JŦD�5<���l���|��,u�M2��J�h�l��7<�x�vi���a����.��@������sbC��@�;�°l�Q
`Z�{�vL�����t�ּ��}��n��>�2����F1���"v����:�.�F�uC�  ^�V}d
�?Q���s��d|��z`a&�s���ڻ:�.�t9��m#shEf������ALnV�Y�O3l(?	S�D>���Qnv4�=kG�,@�vl4)�"�k�>7V�>�]�Q�G�����
\��͇p��+i�SDV�.�=R�2�����\��4��S�k��ԽTpVd�����ƅ���W�zp��/h��]R(�^����ts��a�?��q���e�w�K���5ĊV�*���4M��N`@^^��f�<�0���M��T솴R�81c�8s���r��P���W��!<��dd-���NruĖ�;��ǋ
)|�=M�3d�r.V;�k)x��丯 -�e6 )#CL�=��D�� �|��芊�!�B/&�5�[}�@=]�	*t����M�K���$.b��bN`��j��h��m�h��%T���
nJ,U�p�}޶os�մ߄`��CZ{��
` ��m*��P,ѕ�[A6
��|�0!�F�����W�&���rO���bn`p�*�W/�׿�<j0�� 	M�Q�_��7"@�h�!��_�g!�S�KG�}�\��{?W�}<���DL�Q�S>:�Xy���,��1���D�ߐ���^�x[����F/$�F��
�/ �B��e�h�OT?ی�xM��l������I�3@��S_�/�2�7��V�t�9��Ʌ掕�?�DL�>%�MY+��h��\�V��n,���342mj?��.k����7�2��{�+=�Dz���v��4�rJ6� VÃ��q�+N��BQXK)�8X��N�l`�_�(R�D�	w�{Dy��(0Ϝ��c\=�4�H��o���ẋ�F�f2�oT�Q����MH��"�S0��{̼�E�m�+�Nಅ$uW��lҦ&kL/!~��� 5�o��H���:����&�G=�5��d���X�
<�@���Ӆ`<pъA<��1ެt��D��Ɵ�RL�tq錙��N,�n��� �B>á��p�)�@�ȁ�\-|Q�1!,�+~E�X5��n���5K	��^�*S�d�6~5_!��С�)�g�}2�)V�R�n%,�������B}��4=�郠�	���@��%={	����y#�ϙ���a�=��zR��/@A\����wq=q�:�i�����y�Z���VȬ��RI� 6���MK��~�~��%�ݐb|�}�T��SQI���?�R'Rdv��7]v�1����� �G.��~i�Eu�>2��4 �Ӟ�Wn��2��|����W�e���t���C�)ѯ�r��A�.e��8�7�g���?gO�@	z7P2��ؙj����L�lS�T�4�9,Yq'+���'C�^'���R��$nط��oo���J�y��1s��u�џ��2�%Q�*a�C�����e�M�y��z���,�3.&����m��^ l����:�ϱ8�*׋sդ��GGzI����&K��P�{>xA�yw���Y&_���?��-�Ҭ��c��Ic��K����`��|�i�_sx��������mg�X6��@�����v�_��s�c��6�I��a�$��h�6&q�=�d�x�@��L�d�b+��T������]x������-���Oe܂�`
�"��>ًW��[ʟA��:,��T�	���o�x5K��3m�ARWN�-�9���0��s.�H)g�X�)��&��E��_�nB�j����M;�<p5�I�s	��xZ37(7�1L�Rhg��0��>X4���k�?+�P 0��U~b!S*���_9�>�^/$�D���<�'fq,�,�V�OVywpݏl�/y!~� %�An��W���B�#D�,y,L��|��a�JG�J�T���j�K��>{�FV�u�txg%+q��Ɇ�������c���fEu�K���x,yfz�*�5���y���Y��ώ
�҂� 9?����'to��!(��w1�`o.k�O`�r�1 �H��L��ߺx�2��p[ClR^Ώ�)��r
<[��l��𼶈Hy�_|�Apb���.���q-�דS<tWf�w�r<���|�d*�C;4�����RH8��{���$Ly-��� B�ըs�Sź�*a��S�!���i4
��FX(<�&��3�riU���O�O>�M�E��gj���s���= ���}:cK�!���m����k}�t1��&�')��B)�����b��t���`o���c	���`O?�|V�-_����C�=���$w(�w�D�����{Ķ�:j�J�&�a���Ŝ��x���/�2��i̦�Hq���,�A@�׹����t�o,�$�� p*4Pk���<��`��t�z.���s9(�����+����D$.^�Wx���t�0� �y���h�+�?p$6Ц�i�����pz1��0�B~)x��(X���|�i^�%��@����8�d�0��ۉ�Y���ߚ�����\[��@���-hLn��Z��G�M�A��1�n�sW��0�<�˭���8���
��ߒ-��yd*����{B�.��d3i��epI{
�`��Y�J�Q���&�.{��2�kD|�e�į/o����J��i^FH�vJQ�i�]
���	a�Y��Ԅ�E^�i�WP��|���K�Ql���������m�V���!�-��lg��1�����L���PI���$��#��Ѷ[��� ����Ժ���o�`��<�1�oߣA�	{��[�ێXa��O���k21��>��[�?Yl碦UrudyT
�y�S�D�6���[���h�e]��G4j��t`�ʛ?�J�.��O���i�`��L맣��iX�+ۈ���LŔ��hwr���G�"hwR�T�oR�SgB�?��G�{�n=������P�1�.�Hb;�`a �έpƵ���������)���M�Y��BS�R�7�*>�V�aPEw��4rD��(��&�������=}�%�&�;>��`K���b~�/�+����:(CJ��V�1n:�Z�J����܅�(h����-�]�N�?L5����_�h_�(7r��V[�ۢ��U��O@#\ƌ Ecj�k�]��T���2mV�)���q���E�w����`����Zn�/=�oIϒl'A����5H疣îW�Umip-�
��â�|�q��?���,uʾ��a��*��oOEObkl�����49 ��hɞ����%Z3��2���6~>37��o1.�����ܭij3)#Sv�Ĵ�^���2˒�fb�|����b�|gx_k��0k]��TJ�����)�:�-gdB�$o���L�C2�ઙ��e�J`�]�oZN@�|7%)S?e�%RLLӷs,n��]]�t'�4��dc;���j���s��ڷ3�Zw�橚�����(
 `�ܜJ����ejн�2�ǡy�&��>�W�`��<�r!���g�9���������1C�-����{_��� ��eF����s%����x�:׺��p%�D�4��ȓLyD��F���߁ţ�e��7z�R�th��]���}}7ɯ�$��R�/&�^�aqpo�1_���
��|��n�2�pz���D1��껀V��>&Ƃ2!�c�p�c;��R3��P�g�8�l��i�������>nf�G�8	<>b� ՠd���4>���P)M��T��}ӝ:rC:�<Yx�aY�4�>�n+��*��9Ӳu��]MdR�U�W)�`�8s8ܱ]����Qm[�$TS.c�6a�p�*���Ŗ�!�_�oeD9����ƅ F�}F�}��i����˳?o~
���xܖ{��0%���c �ˣ�Nh�}ݱ�z�5�.�����`� G�c)2	Lm�)�#��>��'��������#��,cZ'�a�5��Ƒ�[�>W��/U~��?L��Qzr�xy]ͬ����w9a���;O�;o�}�CO�~u�����⸛E	~������4n]���\.����~���G@@ n�p��˻d|-�8�jt��`��|�����f������0�(�&�.čn�1�|��e���^�X��k�m�Dv��t���Ռ�	n��:p3e�w%���b������F�{�����"�J: ]2�`c�<�B�\�n���R�84��>aԙQ��^曃Z��e�'ًv�d>��S���Q�g;�"�)./H��bm�,W Nk�h����Q �?b;'�n�F�X����	�qu�^}E��s[w�6M2�PS7d��������1�H>��x��Qi����HG��1><�&�tAk�'���4�C՚f��
|3����$�.�,j!��5�t�s�)�M���ή0�h���}��~�#q�l�2Û�������0�o*�m���p�
P����x�2�+Ɯ���b0Q��й��sD~�F���r�h
�v.���ەA�x �z�<{��Q<�x}g��qS�l�]�]dl�)ԅW��uK'�rU1m��!kk�g��8)S&�vgO�\崈VDAO�R��Ah��\�9����-&�$�\�h��,�_��&Y��#E�� � ������#�uh��S��T��p=б�~��l�x�0G�t��h�]�Rn	�[��9! ��6��_/�2�T�@h��b�H�}�[@�Z������e iA%�����Ҟ��3ޔ��]�;%�d�K���Ɉ�S;,)f
�ѕ���J�?���Ǻh,e���7��@�wr��̟)�o1�n,XN�5]��&@Dq�\��þ#G���;}Jbh�|�UY�����S:��c�7���!�D$���N�cW3� ���:o�SD��,O�|ɾt�X�Vp�zq{�DV'5�OW�¸��N���r�lg��2���_�\E�hv��t�`�'��!�J��_�#�mf�VO���ƌnH�'C��� ��y9�m�y2�)]���#(��%� $^s���;R�!�=Ob��[��'��)�����E�~���[G��:�AS���xA��}z�?Ix�?��؞6�.��shǘaZ�"˕a}����Ru��,�"��tb�����́S�N�g9\�D�h-�j���m����w���v�P�ڷ� 8�� E@� �,�����:l3#�a�v�u����k�I�5� ��2��Nj��~��)/E�B�G�/��Eq@���E^����NugyMO���(Ƒۀc,SnYɽ�R/�"X��j��w��T�����`�szy#) �.ݪ�!�}�5?�0`����&��h�"�.�s��s���My��N�h�I���ɰ h�Td��2�Ayab����� �$ը�Na��ʧ-�@X�Q���zi��:M�9d��'i��{�LrV���}��^�Q���m�>�[*Å�����ǨO�dW�ؕ���<��w9���cv�����rP�g��/^*�+����;�B6�U�<��
��?RADF���5��b���J��H���i��`�n���I���8gR��/\��;k���t�OeBJU�dL;F
L�i4�Ĵ���� �be�S����K�5(��*u~����q��|�,��{��~�0����\YI��П7�'9D�O�x ŲԲ�v�֘�O��oA������!���[�İ��E~�}�!s)__�����j�-��D��I����ցH��3y����LKo��J-LhK
�H��|t=�s�P?KP���h藅�C��b����II0���f�O�(MI����[��\Z��i�n���g	��O!V�.,ʎ��r�	��gUcq��S9��]��КX2�Dp���
�.h�/�n�J,�<8|&#�c~H��R꧋�����Љ��nd��Y*9�f�����!{P���7{���U������47G]`'ɡ��L�
�E�V�C/�Vep��=�ÆP�Te`�V���3�f��n����ʱ_,�:��/�K���-Jy�[薙�`��G������=��ȶf��}�A��,���3X�7/w��
(Bx7t�,��g�[��j`�l���/@"H$��nF깆�-R`2G	0^y"��A�lq�^�.�8�%��/j��58$�n���Ku�#	�J�?�k|䓫��JT"=�Ҝ%b]D���^�J�l,�f�b|91,�s��/v�)8Ϸ�zT��Z�:E+��*�,^�FN"���ȒN]� ^	k���x~�ߠbr�xf�9:[��A֭�?LD��HL7���-��b���2P�k��I ��n��	T����ϰ=-��J�JrI�Q/;i�]����N̉�J�{���_V��Ђy"'E�šE�O�7���d��P�z��`��8s�k���y�@���>��ю�Jyd�8	lܫ��d3�,�շ���u��A�l�.��C�V�߮�XJ>�5���·kY��L��/R��β�0@�"}WTh�#���6����Zq��(����.��B�����n<RE9����&�e·�
 vvr��b������FM�)��`�#<-:��Җ��Ro���{ޫt�(|	˲�����r����l�0�f���x��M���wLT�A�J��bL2[f<��F@��RU�jLX�S9�"�"�1V�i�d^Q�q������LȔ89�1٘�M�"l�U���\;u$�a�Y���OV�,9�[��|�m{
�3ț5������GFj��?�,��M�
�7Iv-�l���l���a�v�أ��Z���
`�T9�1+���.'#P�R��)Bd��K��Ԃ�u[=�6k�̧V�B�:�A&Q���r9�9OyR���O1��A�z��W������kdd㢫`0x-�곒��K�+�Pl
����yu�ϼ_{���q��Z��~L��O�������'3�7�3;H~�"���r�7�%()/�Ru[����?|���=kbzF��Bw���?�;�1�2,��ZՉ�zM�E���$�x�)E�bQ���Ĵ-��y�5b@[�fE�o��Ca�74Ӗ���;��;��H������`~�gL�`���.|��-=����v�RN���g)��Z�3���R��?�	U��p�Нs����_�l��v����8W�չ�8��Z���v�Ɣ���DaNp�Ke4�Fte_�ÑWdO��g�VU~@<?-����7
�MM;�mHa������͌x����,��cւQZ5�P��u�++��k�s/"�h������C~��-�d�XN��v���b����X�%9S�g��Ez>�"E� �^�Q}<?�� 6�	2�-���� a9���ذ�Av�Ǝ�#@�n� s�U'gB\��Z�c��~��n�Ci��V��_��2k��;]G)��}^���+�^N]qpuN���a)h��͝I�<���?_�O�"�>j��t����˧�bu��09�Y:Dణ^u��fQ:At�s��C���%�B*Qf�pȉ�2���3���uhPT|���좚�TL���s_��IM{Z�f�*����A�wue;:DQ�d&mX�Ý���#�0%��l�-v9�� 4���s<5�Z_���]5��Z�Ѵ��!���ټ`.�)�
�o��Zｋ�u\A^q�*M9W��!�?�]0ޣ� 9����[���,�2s/�P������G��c�JDm���c�1�n'�,r��bi��s���\\���V����l@���F���=.�՞A�jMO
Izi���ʤ⁇�@�/}F�O;�,�G��c;�N��l�1�U�f��%��{�E(V}4z��w�kb�l�>�B;7
`��4l������D�C7m��5�1C�'�����;S�kCV�'^�s����T7<G`��y��ĉ��ׇ��3�_����缲=9��j�on���h��@��-���!%C���*P�X㪡�57�2�da �	���U�������8T#�>C����4���nkCXV �qE��� �n�ٿ�5(�=R�������1��������i�o��Ox^<K={���;���7 g>��L���n֛� /��< �#$��[��8e	Fwd�g��o�Hv)�Vrp�D�[.�E/?m
p�V��4���ݙH�<С�i�G�W��\��@����#��S�I?�UT�@��=�^n������5}6MWY�z�Н�-X 't�@��Rb�QH������]h5��u>��چ�Z|�%�H��_�'kw����e+�6�q�"H
�� U���:\hB�!)JJ�0�{�%k5�z�+�y�j����&��3ƿ�j�_��mzn�h�]�M��B�R]��f,3���
j;tt�k\�����ܶ)�-m�N>�Z�gs�Q����_�Xu�	~������pۏ,��^Q^��s���\b��OBņl[&���q߷�Z��� �K;]}9(|l�g��t4��?�
����$HTEd�H@?Spx��������}�����Y;u�0�T�U�bo���w�����C��/�NYO���L�L1���7L���]/�W���0�U� Rcc>QĎm.�H���s�{L��P�FB�o�˕��e��35�q-�2t��Bk5��c��nH���M���^ �Gb�}	��:����"B6'�+����{P>���)>��=Ʃ���k��'�?q"�b��3��	w�G�) 5����u�G�ύ�5��V NB�J���/M�j%��ӧZ��?��[���>� �V�����s�Aú����S��whp��ڔ�z�h��������,�X]�I���(��Iq7V�i�Msf�t[�j���3i!�v�[%��]�ڿ�D��Hh]>�YZc��m��ʲ���B1͊F�:�<�������!���6���\����)��2���H�O8�(^{�����9}#�+�#�Jz帨��O�����|.�ȆM��?ﺙ���>,����j�(KY��]!x�i�^�D쭛����YG������}8�w0�s8���~�J���B����M���M���`0AXT�r���^Ҟ�C�ƵG����Y�ۅ�˭��o[
7�\<
���ؽN��O�u�nk�L�1`�,P?�'�	N�]��.�\�j��I�S'x����5�0�(���Y ������si���"7)��j��@'_�V���]|sS�"�7@~ Ȥ�1
<��ߡǆ���g]� ����a��d[U�-���ͽ�X���] V�%���##x�����%��D��fF�	R����Wa���}�sf힥&_B��ޣ:�9�8P_��N�8,&
��\�	�� G�a���d%�,hl�~�X�b$�.����W�X���W�K�.�'O��aY�v֩�L�R�7�&�׀�4�w{���7�i�]WD8"�a�{�.�Hub�"�v(�H'��
��9���]��3�~#AJ#���sz�Baý֐�^��T��g��Dc�I�J�
.��F!����7���#���w�1��1>��bn
�e)�)[�hn�e�'��I��
���Ͽk�ۙ�'JPZ������ۑ&Pɽ_��6�����K��@��^+�~dq�w`C���R����)�~�*�]�1%�;�:�QM��������xY8L�U�/��S��0g����MJa�"X���[�Iv�V���:y�\@@�Zd?\HY��|K
�A�ODN�����P��J�V����Α���թ�lMV�S&#sÂ�������ʿPJ��臽O�+���b���#�v�B�k���'�=�2D�dHwk�2���&�kM���6=t(fb�1�\R#[p�0���v��f�$�s��v���A4%���K'��k�e�<6@a��5�F/#��T�2�m| � �@�_?]���bW.c���y��sni�WY��x�)��&��P.�ec�WǺ3?S�����q���_����l`��}�ᮜ���S�@��Z��R�c��1S3Q�U*�*KE�zY1��aF����d���.]>��$se�����䯿Q�BNֆ#��b�V�'���"ס����VΦ�~ë�\\��>Dܐ��2뾘�G���Ŭos�y�ᚉ|9w?�y��f�Dy���I$N}�gn�A���3x��Fp0\3|q�+5[A��Z�s�^��>҇1��*�7)���GFCe7�{��2�څ�M�	F#� FO�r�-����H�@d?>�yi�n ����b#� )p5`q_o���B�湭�D��3�#�!�>�{!md�0X�K_�����P]gd�
iQ��_=�e�RJ�)t&3���|�R)��Ď��?
 pڍ8|�	��'n	Eϥ��aB"�Cq^L��%�I�1��õ�!����{�8\
!�58&wg�GJ9�=�*ʶ����=O���,D~:�����1�:�Y��K�Nu���䮸�^��H�k7���R��ZB���ц���I�*��םt�Ⱦ�_�tKT̊�(�{�J��4�P-���;�?D]^os��E�Wު�zi�cvQ��Z���C~$@��ЯX�E����ss����%��"�S�hgq�S��t�b�8�o�ER��&�S8�D��D��:�O�K�θWڳm+���cͅ�X`F���U��B,	x�ϵ��,u@�ᖅ���}Ϯ�~B�EΘF�sE랬����#���l�Dl!�U��#;i����ek��u��&�F}$jӨ��c!��(;�)~ɹ��O�v�։M��z�K7�9�������"�mY$r8I�MQ�r�;Kկ��6N��b����R����I��6�gWʢ��������
yڴkܤ�1ƍq[Q����)ҩ��� ����>�9�� Ҳ��6�G��yd�f���W RyI%�h�F>"�Y��?�d�n].����#yM����z�ś����B 0-�����j�ַ�D��I���䊹LU� �7���\�)_�
G�*&�		���a�~��-����d����(�K�|�-��S���!���-�n�K�Lc]D<���jUGܩ����� �������_�z����'�"2:�_rc��3�(�F��8o-D� ��������5��46�=�h.]�Ү�'�L�Yx��x"6��vҙ�Ý ��YǑT�`�������n2���2�'�;CK���٢��= ՛D���o�N �'���M�8�d.��C�{ i��PG��8ZvL̵�jf�:"3��ε��w��'�oM����#2n�r�Ře{&�����x�NhVg�Y�a�琖
ע�f�Rƾs{����OJ�y�p��1��@'���_\���L �Sb�� ��Ȧ�Ru��ٍr�tAah�Ƙ�y����N��EP��cC���QJ��&����34r�ן\)
�@��\onA�y���
\9������6|ڎE��n�����D�I�ea�� �Dh4ÇFvt�����ρ��yX��q�ثk��Ȏ�r���6�'ۘ��D�?�uޡ����0��d?忶�۬,�����ܭ���Q[?N�V.��>�ǲ�ܙ�2.7cyӨ��@)�}XL&.ru}$5���.z+!�i��|�P<o&�H�� ����{���@��%t�pZ7��٬��I�Ւ��X$��ba/@���(;�>0��C��'�{��)��������$s#(��#����t�U���~o�G_�;d���.\.��$����OA!��aN��5��j�1sp4�pw}�Ј�sx@/��Vu�S/Ż�@dw�=��X�P�ӥ�K���/�$Ix��G$T.^�Gxݳ6�_LE��r
��׎���ۗ2�a�<[�Q��(w�{Վ-��������[i���Z�wWJ��Q�c���s�c�v�1=O�Į��!WTعC�S���q�|��3˩��έ}��܁)��ܭ��?���l6��/P�C��Fn���H%��frr(��^re��$��y5�ІSB��^�����Q�%?kADܶ��:���3��I���\	������e�{���	n����g�{�2)F���_=����kRfu�TNa�|�qa��S1�b�����n�u�k�Zc�R���s\�~�U���6��K�7���*U[�-xy2�p't ����vw��HV
�)��Y&��H*�PNe��QSa�T�2�}�E�H��ߔs��WSg¶&�T�VX��R���S��r<3����eV�I.[�hh�^�0&��X� n��]��mw��-���ZwG��]�g�|-��!S!�|0[Ժ(?"��˾��3W��:��"�� ��w�8��(� ��KT˼z�_�Ի@�&�v�;��}I0��;N���U�����O��������x]B^��x��!�j<4$���rh@�!
l�0���ȕ�\f���)͋��̵򻝃[�;��[�D�����Y�Ј\���<Q�)�����vD�U#��PoYJ��8� ��;���עCYH't�����}��U��IT%�ԃ��@��},�u�]�sH�m&�_t� �Z�Dr��U���KrP˞�kn�
us���4R�؛�V�N�t�ԻJ���~=�
��Y�Bb#�7� �FA��������d ��x���\Ln��Y�����v__>83��>0�Wٟ�VPiP)�J��˕s��7R+��*��pɌ{�``����E&U�`l��I�����d����~�_3;�Q?Ȟ�f5G�5��Q|{��1�b�9��bx�j�Y	5��D� �s�+U�5
���"���X�'�m1����\�e��iPӿI?)b=���݁	s��!} M�\��M@�`�%sݒ����I��l&1����TS��^1��S���������	(�D"h��ܦ��଎o������ވ����T�ҍ��6����XIY.7
��^O�]�C|1��}��auD��O╾���o���ß�B��9�x.(�b�x�3��s"/d������_
G��{.d����[���.ͮ���^��W�P�f��NDU��{��e�i���Jq:�&�C
���ۧ�I:J���̉��03b���������P�ern2Zh*��.������s4R�'*ʜs��?�v���E'������3�0b�+����	�m�zy^��u̭(Ł�x'�I(_��<D�ݪ�=�AϦ����u2~�{|��X�Ii��],"ʢ�GS�i8��@�g��]J��)��x�N���7I׼3ZZ�j|˵"�袇�1WThSz��r`�����WՅکI�����n6��҂��a�i ��oUs@	�Eh�8�2*������D;��9@�<��g�&,x��*���w8+��*"ów�»7\e�����OJ��,1yl4ɐ<����QQ�(�΀2050ECo*���-nSw\�Ꮛ���O!�}�{?�7]VSE�Q��~�����=654�\�E�t�v�d��KH����c���Sk%���A4���%h�{0�k����v��ة���a��8��pO���hU5�[2*�ƾ��K��g�x�?�W�l��Ez���_�uŦm�$ް��ؽ#��@���1�V`��	:�¬!^��
!�������\�ޠ\��9��I���:�E�lh�G�ფ��t`?�~�
?K�u�\ ��G�vM ��ء%(#��q��z|i��\�1|������>�f��[a:L������`
ۡx�p'���L��q������$�0�H��`�ߑ�W���6�Dn��#���A��|t�m��{�K1>�����G�ɗ-P��"�h�6B�'���8�����8���5���E�{��@ P����b���W��l��&�&"2�g���=%��-��g2�46O��:`-��kZ���Wv��D'�r���	S��V�����G��A* ������^�`L�51�y$��(+Pa	�g�\oJ��UfL�P >gRc����r�B@i�>3_�2�٠$�%JڀW+��l��?���V?���2"�4�>D�wՅh�d��m6�q׬�>� ڿ�/�.��SL�U���CCp�
-��hw3Ň=w������|š&{n��`(߲�,ऴ1�S�{|�ǯ�=��4s��_[ͥ�ƣ�m��ǂ�c)�7U,��p�Om��r�2�i�ƋͶaK\��Bݨ���ߠ׍�B`�)|3�4�a�4Fe�`F;l�"ļ��pX��.�w��q����*���z��LmWS]��zG�N�/�����te����8����Y�BU�-��n��(0�2��f���S�}�^�f�ds��I�Հ�pk�z�����if��
��3]�/����6װ���Rcj�t�JЕ���Q���M8֢��h܈�o������4)�	����ߞ�}�'Xʹw=9K%E�����0%?F�Ჭ�t5ͻO�ތ}a����(�-(i��zڮ�v�n�ǥe����;�F�K����b+H�ε[`��%F#�5P����|3���#������m� u��wӍ���~���Nx+��5��w�𴤀�'�ql��W)Q٭���rI�+ѝ��-}� e����V�������K�\+f1�Ad&L�2 �
�`c������ /p���Q�-NJV`�OP��!�b��=�!�\��`R�G<|�u������B
o�
�-��BGcN0*�s��3��o�K����|�a�p�1u����VW:kO5<�r�M+����ϊ���SA�� �x�R��
�}��୰��F7!O٬L^:��Ir����^�&ҳy)Xa����cW.����i�r�U��k�߭mő��Zz��Q����	��e����t?O�t"�D�Ud��L��Z��M��/;��\d�=g�}�,e����ub^>T��:L��[���`����I[��瞏�|��f^��6�*��@�+�2�YS�*���p�Xut��������ۉI�Nɻ����쥺韍!.�[�p&.|�I��n˚m��r��ֶ"B�˅Z&�]-R28P��Dr����xѴ��I����^uRNqF�¢���;�T��85��mg�4Ċ~�^�F"$Z;�-N��W
�p����j��3PD���w��(0_Q�����I��H;����}�`��Ŝ�?�S�lv�9�QHJ5p)25Iq�L=y#|�񏦦��M��ot�e!a?�Y�>��! 笶�8��i�F�����O�Ɣ���L�R���F0�Hbm�a��?3�yۍ���s��Rk>�K�����cW�b2����hjm��/=ٽ1;0�&��E(���+��k �]dw^�z})RN���Z��T��
���q�R!�\�A|�#��TL=R��ėƶ�<����<t{�:���2��[��{=љ�R�|�I/H�!W��<����D�����|W$�E`a����7i��+�25,����}*z�ժ�k�D�M'�"�`$�Z��A>l#H�C2�(3o�>��>>x�Ō���#ak��0�sC݃��K�XDlG�L1/	6ïv~&��M?�m�[i�gx?��<'?b��M�\:>c�۰Ϧ���vDP���b��q��(P{��Aۉ�ټz�j\C�v���l7i����G��M��ia��'�cX5v�
�x=���Q�7B���|��Ms��q�yۃ"h����⣮V��`L8N�YA�iCn)��1an���.�A�%h�}�y�-B=ځ��㓻;:�O#^�:%��6XB��}1�Vb�Bh��s�����߆�n�.��p
RL*��&������^_�V�E���%��sp���w8<����h�^
�o�N�'sy���ET��>�!�Rb\��{��6њ�;���q�B�����*{�v�&b��({���U\�
���9ޣ!(ثwU'����,�Iw�rI���w-8.y+y��lHtqLR&F�V[����ms���%��S�\0�v�8u�wN@gH��I��P���iK<�#�5ǊQ'�����I�/�%��/֍�ĿS&m6m��իqm?�^�w0�#��#8äx�705Vv�Yo���E����O��Hu[�5���:3��}�	�Lِ�@�w�bV�]��<3�x��i�S�s�P6'.�H����Όxm�}�ǵRXp4��[/ci����t O���u�[�����8���I
Z����+>�,�ۊ>�ЀzE+8��cl)<�=��y /��"_�S����^�8a�������lݪ�hm�����I���
�lO%@2�Ԍ��ѧ\mz	!�^�)�ؙ��p�T.�DD��T�s������"%yJ���'+�G`�)٪E��ʅ�J�uV�)<����L�����O%J?�X�����L����q�[VLn[�����'�Ƙfx��E�#������ڭkS���q�Fl\͝ѡw8BF�E!���r�?���x�7����+���V��t�=�a���xwx���u�*`���q�5�8����!@Fn�˗~���u�佝��4���$ϐ~et�S�:�g̽�A�Ɔ��a#X�U����Jt��^y�Ǆ�'%�ȗ�4]�/��&N������D����.q���Z'����e��a�/��@����]!�껚5� q�bNdIX��o��-˽p������))�f�J]BW�J����#G���"��RA�q�ABۧ�+��[�����i�i�K�ؑS��|�g���Ě$��H��Ժ?�^� ����=b��A��BuXG+�0a�u
o��&���naă��Bfe���)�ׇXx~}��~2��4�P� �@䵇*j�b�D�B;"L���@:0�#�3z$ǵ	1R��~n���D[��?w� b��(rz�r�o�Bs?�9axz�e4D2+���U٧�:ʪ�C}� o!���k$���m�W�d�����Q1_�ehRFD`L�ĸ2����7���W��V�6���,����_��|	�v���RA�zS�	&��QuJz-����O}c_�j�ig��C23�8z�܄�U.	���`s@�؟ p��*Α���B`?,iiZ�Ĳ#�+���j{T�� ��{�J�U9	���$�]t�o���T���k��O�������Oba&ݸ��o��yU�'d6�^:%ZƁ��ݕw�)�H�&��Y�PD�W�qÃj��h����q�W�|.oh/�F9���\�?�m|�Ա`���0�Mf+�fI�VRWEl,��M=�JҺi��m�;�����B������P�{F����G����V	��Ѩ&5��S������I[�<2�O�6���6���ӟ����|������ߒ�w��{���]~��GSk�ǰ��ۄ_U�����V@�M��<�:���dJ(z��;AT�(����"�o-թ��<���f�G�j5����T5������[���X3I#��)n�
�y!4G�v���1��42�T&����][�[�>�|�b�s2C���#�|{��?^o;h�N2Da�����\l'�v�Q�H���ޔLG��'����-f�Y�ԣׄ٧���yӃ�sd�St�/�����(��������b�Q�
�#����4qd������a�E|�%�Ϟ���GYy�8�(-�8]$� ���}��z#`;�.D����|�4�u�H�q�ƕ?\ͳ�u����0��'2�q�dU$1��$�4�vU�&��	����><�ї�d�X���rȔ�(<��wX�����£��Ň�8�I��p?�TM�Y��F<vZ3i��\%}-�)�Bz�����p���d6ݍ2��� �e>f�*�= �{n`��c��q�a^�P),�
��k#t塅��CI���+�����z��@�KӵK��@:끵i�#�e���vp�)��8�� i�(W :"Nd����b��F�C1���� 獈r���C�y���B����^�twg;Zڥ�r�5���o���@-���u��zTm�<9ʏǏU/{�pT��/!���� h�4!�o����ZMx(�6S�ppZ݈�!��/�	S��GB��DLF#�9 H���	$'K�����l[�$��c����͎5 �~R��|GN�/�`Y��ek���׋Z9}ȳK� 붴���oɰ-_�1����-� �X��U�*/���a�_��#5���#��V��&PG�]J#A
t� �9�$b��!F��.n��ɬ�@����X1�\�6Z6�Z�* ��n80 EKP��Oe��zp�:����Ze��c����h���|�������<<@/�������V�z5�iI̍�=�Z�� oXd�$Ia�W3@��w�_E�N�fw=���#Vl�{M�F�6_��"Nx��\w�r?��k�i@�y�C?��5�?�!�K���[S�Re��j����P�Rψ@K�`��������wh^y��+�ai�\����ޝ��� -�o��X��g(E�RO����@d	 7|�m�߰�N�T*��&Kyug�TP�%�s��>p��m�\=��DGCI�'��C�[&��m��9f�z�C,N2,du%J�ޯ���]q�OU���P�udt/��K��|��eO����wS�~.�ff�*��z���[�TF���?j�����?�؞A���~Ё�"kp����h�X��T��V��a��CXp�F�=x��=���V��_��w�V0���,�~��em��x�/刓a?��a$6�%@���EW�7�!b�'a`ͮ�6�No�$�� �J��!��S�W���7��c�K�=^��k�,��oyI߳��da&Œv����")��gL��{m>#�Ļ��ovY&�e�^��̗Bs��i�����_�e<I���>ӜO�&���flD��k���c����������!�J�����M�u:�f�LL��E�P�$^|ʕ��9�>���m3��I6f���4R��u�����$f�;�w�|ހ���&��b�?/��r
��s�G�4q��5I+kVkk�Þɪd���1�N\� px�3�FS|�dZ�I_�-kO�N�n��k��v���<�g��Y�L���������x��t=!n�E�k�~���4��V�#�g"S���_ٯp�C+c
@���_�M�/h+BKNb=㨹�lC^T�4{�hАC|s�0�UXGV�ѡ�& ��5�F��.Y�^ק2A�n�u�_O�z5jEu.R��!gR�a�Y������(
���^�\p�Eot��ft���""]�/�w��T��,�n���,��񦵤��ȼ*�L�s�a1���(�l��:-K�ԣB�L �ECQX���ޣ��5c�C����;jx���f;}�ߙ��
�be��R��{9�C���~��<�Z�0��7�-���5�?��Wt㡞�?X�:�~� �n�b";w���$��4��&��k|�s~n0�	&��~�Xx�7�!����E��d�g�J�j�,�ͧ�� -Z�c���p&��-�Q���w�$\�Q7�-&�-H�8�K� r��x�{�Χ|�H�%c�Q����s�p[�9r")2�'�T9.�ɪ�#8�V��ȗ�����C���g��Y��q}��/��� t�°�XTE���Viq�*�\1���=�횰<�H�!ғ?����:9���8���lH�96p��'W��TBȗΗ�xޞ�A�j�E�x=9������l�Z���� q��P��&����$uc�fE��"L@�K��i�C�瀤�j_�jN6��	
+f� �`���{Y\�����
�D>?�c�nCF��Ѐ[�]JާiFu�k� f�t˚5f�����ڜ@x��#:�zl�:�a�r�=2Ǐۀ�� ��=�:ʛ6>r��D?��'�Q(����Ϧ�����T�ԈD��U�g��`�0m��h�B��5t��ܼA��~]�uԵ�O,|�6_��|�郸�c���t:��q���r��^lۋ�MdM�h����K�%����LG�uE��Q�2�P�$襔|l��3�	h�v�AZ��_J��T&"[�����&au���􀏦Y\Ό��զ!��#>}E\,=��K��r�h�Őj�����eb�<��h��SA&X�����e�@:~��=U��;/<�L����[vp}���Ҥ��i�P�<�w	��'숉�l�� cضRV�j���%�k��Rr�s ���,e�6�dA{а>�s<��}�7F�ݗWOJ�rR�1ó���j�� ��@D2r�cwj�ʤ����%JT4��!�${S� #���G5h	5~��qN��}��Y��"�3��	�'6���TPP��>��9U��?�W�*���I9?h�^����s��O��B��sR��܀f>��D4��p
���/�#��$�Ķ��	r��'�;"��9=_�YlٌU.�Fӧ`-�:O糣Ƌs�|ʻL8�j,��
��O��0���x#�����l*����	��;�����L
���L���;��kOf��~ ��"ݷ�r�.�vSK��D�V�D�I^�8�{�5Vi���Tq5oa���;����tm{.�<I�s^:�������Ӎ��9��TN��bxGo?�
l��#�w�cqի�EI�/UĐg��9��H�l��cεl�G[�_S�=c���IpM�˂u�d7���S(���7\ �U�~�h���2Z�������W6�6V�=�����S��L��,ϱ3)�]5�R�K�:زʠ	-P̲(	1eql�S9������,����4Ս����6��dd��w���j��5һТv1\��N�:8���D�1 �.2���r��q�\^T��[{�p��,�\�E3q� �G8��gh�遘��W��C׻gB홀@4DdE�h��D�'�۝�9/{AoG>�Aʳ���1Xհ�սqΙ*lM���v��qFHF{�w�}��&�4��~M�fSa-�h�6X=�U���W����c{T+%ݍ��u��lJ@F�ngK�c�΍o��w9������z����	�}_,�Mɘ���� %��>�I�Α-��e��nm�n��bR��~����^X/��e�FI��˦e4cA�S�`!@+dɰS�
&����z���O"+.)�\�M�O�>�m^"����] A�
���#�d|���b�:`���o*�
)E!fﴴ��u�1:��s�{IFά�����6W]��7EAP_�q�����K�k��\��g�$�:x��޿Df�Z��fra&���KM؉Ǥ�~֛[&Q*sR�b��ǯo����_�e�:�6���OE�*X%�7s��珆e��&�@B~ �FA�k��7�-�	�Fr��^'v��8�Q=oK�4��$4i��3��Ϧ��]dL;1��j�S��b��b�Sul85|�-���'�)��W��� E�_x*��p�s��
�"Pҝ��f3(�G�}�Z���%�Ac�c���a.�E�=7�z�J�6j��**o�\�W7
ܒL�z
����ö�V2�;��pl�<l�ñ�jo��[��:OWz�����/��t5 �)\�?%���Jʭ��Xo���˙݆؜��8�6�S���XgH7(�\E�1�\�!��b�Z�uXE=�{��
ؙ��]b���TZ���ek�jĬ��z6���v��'�%ֺuPe@�kl��+2%�lg�_��sn7� @U~�|�Z5*;��j�RN.�+|�DbA�2�������X#H%W���]�M>U;�s$�z|ǉŘEBK�f�A_���$�ꊆ�vp}[d5'or5���虣b4���a~"��ł���o�e�� a�+����(-��6�j	���X9��"��kL�^��W���뗴��t-j�����0�:!Gv���ur!�r��B�tJnˊ��2f�>*���E�W{Hh�T�'x�_����Ǖ�h3�ם� �N��'�)�]����}Խ�;,[�ײ���׳l�w6'��J��0�4���U�3�˿E<�N� ��B^���Vg�aN�07�aI�>�w L�	����_�,l�"�q<�U=	�����$Z��q�8�N{+�����c�F�E��R���ɽz�`��\�=��{�{m�'��x")�w��ZE#���S��>n�6�T"Z�٭A֊��rf�-��+����H)iv<�v��%i��K8:��O����&m�Df���)1�����T��q��ȓ	��~���TW��=q`�}�$����4S��Uh֌:�SZի��LOn�
+~�v�ͭ�m�F$ׁ�m�5I(�xs�:�9�v7��Z�I���9#�LxS1I������g,
⑴$�+�<V	g�yȃ�?gX�3h��nl}U�����Rj�?�TeZ�̕E�C��/�� ET�bBuJ�N���f��=����g�� ����M���=�S�{+&Y`��D*��f;E��F�3��q	*H�)dP^*��:gc��2M�X&	���be�������J��YG<�G�`D.%(��#]�m��<]oa�cL�a߁��������,��[i=їV{=KG�
k Ǡ��Ɗ�GV��8^��b%w�A�q.P�� ����q2;,^%Dܧ�W+[r"�i�6��e��YOq+/�e���s\F�l�C�!������Ta��,�Tȹ{=�N���SU���x�c|�N8�F�_w��Zi77_R\�ri�QP��!�ٙ\�
2��;m &B�k�l�d��x̺$n�|���@���o�`C-�Osb3}��E��q�u�Ҝ�Ԡ�pz��8��3�<M�He�3)g�e�5K�%�Āw���$��n��N��7��4�m�dJk�����O�V�P�����Û���y�"�lM��Jz��o$)$Abw��2x��59�$e���T�&�!uST_���aю$��⧬%)?��z*�'/e��u�=�)�|���jP���r��������5knθ��f4?a�tV�5��R���O#Ui_u}.o�)�L!-Y�����pAb�v�>Y늓�n�齜M ��y}�W�~�&P֗���}8�`~C����@�D S��_�	�v�nk�.~d< ٿe;L�œ��i��*A>�K��QG&��	�/�[��dƓ�H)��SW�Θ��/B����S�-X���<�*�ic�2��(3Α�6Z3�}jf��-PC������Wz2� ��}'�4�8�:�#js��8�tI�u��E��uF��|�Yc�����_�O����F���nl��a��$�+M�p�^��`?�)K;����Z�[l.���?"�R���1�3�����Ԕ��ɱ lv���DfXA4�Jű)��f<V���d�?�\%�^D;!o
+Y��~����V����n��q����Ud��m�"�������<O��Tw��Z��c�{���w�E0qp%Ѹ����A�k�$�4��[<0�Nn�Y�6�?8��ʫ���鈡�JUO���{��J�j3lm�	�j�����v�ډ|bI��P)���e-��m߇�K�+�诤��.=A��Z�4�6/�2��̱u�{9X��,Fy�s�9��p�ã-���ՑȞW2^�`qJ���燸aՏ�#�����V�6 B9�Ep���0Y�N0z�2��\!���i̵:9c��a����â��!t��K�VϪƲ̇�F�m�Y� w��if��V�o bR 
[��_��7N�K��u�PmB��h��$����蹺��[���K�dط�O���o��(ȣϽ��s�/��r[�&EG{�!�8�e�cկp�yT��W��<�M��X�r��PZ�������>:&���k�[��İ��o��@c�iT�W]q���犲-���5�R�����[ߪ�s&���� � �6�,m��s�1)�I�H^��|�����~�qY44�2�^坩�\P�~��1��vr-��v
��Q�F;��������9C����S�;�5�%��F����V��j�A�Ըd���/���S�����;��͜i��n�w�_��0��ݏv�DN�O[�C�����
"+�-�[4���h)��u�\�x���+j!?G7�S'ͱU����	�yxOR�
�j-��^�OvD,F�z߮]�{w���dꫦ�+�N�]@̑�_��ȥz�v�D(ߐ������Q�m|GǶ����$A�wV�)�Ge���oz`@@X~HPܓc��J]A�(�����nkP�)Q��u�8�Pc�� ���2��C%c��.!ê��^�R`ժ�5h�a'�G�w3�q�VQ�7��^�b��ڍkGAk���j�c0��A�b>�R6�v?p� '�TL0�L|�B�;�/e:XPHN� �v�J���uڠqi-��넻W.ce���$}y1mށ������ᙝz��䵟�6�(�Jh� �3ۧ�>Z�Z�ϗ8���{��ڭ��u5:f1rh=�hA��ٯ��|���G`/��+ ��Z������CZ�7L�!��swOs4�^*l�@��r@�E��,��x�+�4����}B�J��B����ntԭ���s��I�[��8��)	\�X:�_����Ya^���Q&\��x���j����=x3�7����.-t��l5Qsm������6� 2Tg �E��#�b��B����Ԑ��N����J#��0Oˮ�>��R��C��
}���x�7������RD�A�窟��#�Y��Ԫ���Z
��L����i���>��cT~%�A��0t��Dy����p{�ܢ��R�0�$�`\P�ஜ���)D�o\p#��ω̜�J��t�vD�Gn�瑼}
�z�郕B��6xbC�#[�I���u��*�ycw�T��T�@�e����B�"Ł+��#Xv"L
T�y���7ī�Wt����&:,�m�l	� �-C8���y�ؚ���۪'�����CZ���2X���s��H{'��u�4�app״!>����)�K�ng�X�����{R��;
�`�-�%�G�?AL���VT[�i�	���2x_ ��N��a&��Jp��4.g.��m:rLv�6R���	X�Ǵڎ�8[ӂ��:��BA�#5d��ķ�V�p`��E�r��g΂�4o�R�JPnq�y�
L(m=y�B�8~!/��B�:7M��N� %�7a�
�q���9�<�Pw�?n�0f�!E�I��)�п�(UY��˿LZV���C�W2�R���o	+Z��?�;(���@_4R��&��s��EL���T�"K�8��5+��-$V���"�@iw��V���xnU��˕���=p+މ�Yic�)h�����p��c���*%}D�eW�:;֟���Bak�˸.�b�H��2��4VǦqS�F� �� �{�_�����E���R�Fί�K��1&��.�e�G�8�S�2-���f�ʆ��A�p_b�9�����MM�'��uĲ�Ґ�ŮlFje������G/q�Xsu��^*rϨ�r%�L�M�cQ�&Co�������[Bn�%����jp�FGs39�K.L�c}T'`�+Io�F�m��Oc�pl$%����E��a�Z��0r�c��U4�8ׇ�,{�&C6 ���OE�u+�~~�~���V@+F������o`&��t�S�MlNt���O�P�b1�m�5�C��(�8�~;��h$��|��[ҨV;�@�&��#���`�:�LG�ښ�]>�_�ˎQt�z��i$�1%�UP8�'��?r��[�7�S���v��a�8����Z?����@2���4�sݪÒsu1*�Y�@9��J�D�vz1u�SSV��Zu�P^I�W�F�S�\.e��T���]2����}	����r�Ѿ��/�f�jvt�:�#���#y��[iK��ș�Jծ�y(�g۞�\�F���HS�����d��SK/�}'�s�p�:N����@�uŗ*ﰬ�Dy��L2�q&��YkZ�;	z�}{�vB}R�(��1�X���WwN6��� n��^��1���*���<q��\wV�i���-����"u�N�q5�ԪS�;k��y��X�w�b�F�5/la��'R���d�j}6V!"9�	�Gx�h��$e�)�C��/a-R��/�ڭ{��h+�/R���&��	sh��uőװ��TXx�1L�W�R�]K(H��u���kF��5��_P56b|�uǯHmfM��+�>՚F!ʠ�Nߧ_�
��G����,g7��vΆR_w�:x��;�f_� �&�!S�I\;��."w�C�q�z�eidL��sB�c	����p����~�*��ITכ�Xz��!B:m�`@9��ѥ_��z�;�Tɕ�V�͈ޕ�3�'Jny���Gm(�cAr�E[�4j��1O/�Ѿ�Dh��0�����ҧ��꽩!���ً��3��k��������^�	�E"M;�L�I���%�f��mml�b�
�\H���)�Ti��N������ǈhF�[�G��ʙ3�)!@��x&/�^���6!)R����͖�G��Ha����� Q��|�YQ�#���D�D��u�{�e�'$�$�K0kmT���=$���'��2<�(!��F�=+�)��Mm���D����y�!{Kn �"�y��$�Y�Q%�}��!�O!+�&��F�l�V1�Uk���*�'6XӅ�+-G]cG��� �=d� r��q7_c0+#�3+l
NJ��k
a�}��ˬۮ?���/#$��Y`�i�W3�==�,R�ܲ�VO\�J|�)GX�W����=p%!�pj���d�^�p��H%T�m��ȉ��&�2�)��T��J%�-o��֦��4+Ǧr컜�h�~C�s���=�(���Y�>���c��ץQ��� ��[v���95��CR��jOxo ��HU�����GR���K�i n�I3�-���[���n��'5�����Ph��0t���S���6�c#����8��<@�����ܧ�}�s'e!:W�X�D���]:�y��:��4&"�n*R74wr�By�k�����-ȿ��CS__}��
��w/��/B�Z>$��k�f�?��x�O�rָ|&�rr��/Bӫ���|	gP�G���IQ�[�Tdݍ9t�W�yF���lN���N�[���H�?3A
�i#�a	?�6Y�H99��4]`-9&��_�]��.�d�� �.*ˑD����D��N�7x�xȮ��h�������)�X&B������g��g�V$�~��U�Oi��ٳ�wf`VDa�b�&�RqU4b���"�ȓOݗ�ٺ����j(��>���Dp� S�dZ�}�]$فunc��/d�?O��a��%4�����\�"��6�<v-�_!�{���UN��J�-CZ�e
��A��2�q��X`>�~���;8n�qH��K��]t��j����6ȓ~\�a�r��1p.rv�2�c	��%�Q_���r�2%�A9f��^��3DQ@��?:�v�,�}��/z���Bv�L{<�;�ז�#�������© ��?��E-VCd�+��tb3v�3��,ފ\s��:���c�_��0B/#���ʶ.<ݖ�MQ�� P�6cS*7Ǔ��|�]����M�p����^٭4NH���y��9�,�����X��W�~�M��D��x����k�i�D���P@Z�@�z�;���\�Lʁy*u��������Z	y� ւ1<u��J����i��ҡ|��T#�Ɔ2`�#���m��4�*�\�N�.:o0���ss�і3'e���oA{��!�  yo!�Պ��`D/s�5^�0�9�MP�x%�.d*��vM�Ij�-1�p��q|-�C���c��qPE���M?*�p�#�sh���1בt�)bFXm6.�Wx��AV{h������]�PZg证#��(s�ɏ7j�^��_�t=;D�<��'}>���a��ƴQ�2��E�?1�� �����v-6���1��}����^	�a�eJ�ZKqӴ"P4��zL �q����yҊ�Q���
���*{��ou~������aV�%�j���`����C2��^�;UA�T���6:Gw�Մ���^j��U�,�ꬼ8m��3�sj�o.�f�O�b��V�Ű}K�}�%o�GL!W���Ķ�U�b���~G9\y��ZsY�h aj����N)��lȼ�-7�;D�SC?Nc+�.V���`�G�9ɼ^;t�/�X\�{��b��^b�/_<s�q��Y��H���"_>�U�j�8 �C��d@OT%�Jz:��	�:v���?^��=�c7ޒĽof!�c�̇Ct��O��|�� U9p��JF��0�1p$��x;9:	�zPL�]��J�ea�VP�}�M�kbJ�;���^usE4į���J�b�zL�F��P�X.o!��#0�	5�r��@�TQN��vq���٫v��CD�q�����t��z�T|��@��.�`�E�H��k7ڨi9��n�J��b����A����ʭ���20��3�������ZP!�.���6Y�ٙ�{OHE�u�~P������3�Z3ߍ�����֫�٣m���P�{�����7�����3��|UJ �ݰ���f5E��\S��Q���'�nR��9���Q�c/C��s����U#�o��5!��T�õ�G�?�����(zN�+4�=�D���s�nc^�ZSEkX�bwKͮo?��]ώ�fYҕ��֩���ѫ74��n���u��������z	�aүƴN@Q��؄nl�����J9��cp����	8������a�zX�7�>i�}!�*��^T���\��h��&�B�.� A�2�"E*��x���m�qMf&��
��c������(�Uq���K߸��C-9��;̶�v(���l�d�d��N5%� S�;+�
��I|�OQ���X8IQ�H�+���T���� V�y=���Ye�JBӞߪX�!|`b������:���vR����I�a%� �y7���,��^����+�'
"L5y�G�7	�U_j3����:3��S��K�8�# mϡ��(��u�F*J�G�P1X��
���n����Đ5q �6�t��Ni�8��Ï��ok�Η���N�w�~DنA�H~�X�S��V��f�c�V���Y9��Z�x�z3��tB���/��t6�G~~��Ko��_3D�B��[��w
,�L����ȓ�E���h#�1��+�+�Y����28������v;���)�1��O�*>��s�e(����[���4ݾ������o��$��'	�	۽�Q/p�嬈���N��!}��`"�D��\��f�|1|�=��]��T�&Y>��Us�3~/���6�sS6{g�~�����d}Ū��t�wQ	��n��}��Wi]�����	�Q�XZ�D�ٳ�s��_����҆�Z!�*��d��BP}���A	��o"K"�������8����i?H�z�t���5�dT2��Oo��U�Ag��=��	�3km o��~��ZĆ�[���DhX�º4�ذ��H7�w����
1_�.�X!�\/gD�}�9�W(Q������e��lb?�I�5p�^g�$]FdF7�t[�x����[��?;څޝ����b��>�a���$�������������F����cc�r6�g�2����8�>[��˃��8w�ޚ���(LU�*|���d�������Ӷ���1��Y�M�	�������������w�Y�*�a����Z���&ʕi�im���p���w/u2�6�����MY��tb�dSлg����v!�N��)�����oTɢ������4��^�
���:pm�I��0V�&�쿅�������G��ʯ��R�]���-ϑ�ņ���=�A]F�[����Kz���/�U:�bʻ�!��|��{�����i�#�ҕŢ��i
/��:�s'T6�-��%iZ�wo�؊ qD��
�ଡc3�	��w��J��:�%�;�(á���T7�.[=
�:B�������vk�wn�,�����'�"Z{�>����t�ǎ˿�[X��!:��n��,��US���k�����*ӣ:-�,}����2),n�{d���x���l�K1/bC���M"�o�X��%K�f�x0�_�������=qC7Y+��%�i �f�:X��%�Q��E���&�C��:7&�r!QLZ�I}/��jiWm� =�^/�����(q�TL�;��EOgq!y�o�2t<!�!��l���<��Q�XS{q�x$����ٳa7�5���o�1!=VSS��G�92t~��\c(<��Q�K�v����s���}�o�}�����w ,�义�R=社�f1f&�������m:��ƅ��h�%}�����IІʟ�[9�;m�;'r��sH��B8�Ԑl��q�Ѓ��w���j( �	='�2���#:�%�y7�J�FUN!���^:+I�e1x�g�ʤ{l�c�.�"��p�]��;{R'����A�Pް�-��`���Ҹ�r ���a�E�V�~��]�J�n�6c+mz��J�S�<�-��0�T*�x�@u���2�Up�g�����`��x�C|&������g��6j}E�1P���!FT�i����!�y��8�Ѫrnʺ=�����,ie���Q��Wm�;�{����j�rY����<�}��� 5n*}R_�(�W%AF�3��eio~�N��,��=BV��C��[iy��cUֳ��XH�}�X�n�2���=�\gg(ޞ��U)������P9	��d�yں�Ƚ�zY�BV��vn��Y���f�Ђ����]�[����:m�;|��	�!ؖ�%,h��H�6�kE_���]�n�u������E15���<�9��Ĉ��P��s������j�U��]6�I�T_�2��N��>t�1y�.b�/ej�Q��=!Y��o��+5vtf�6�%���`Gmq����M)	�|����5� ?���W�i'S6��H�~���+��f��B6NeK0Vi*������#��������܃=e;�1M�.k]ۄ]j/�R��߃��k�ƭ�`BB*��j�c���-�ǫ|s�+=0�䊍k��\�x�6e���@j��m�nI|>\N��kR���:�?D
���>��u�,�Z;
*�/��W��S>��7QXn^�	{l,T���L2)��v)m[�v�ub�=�,g��+���(���s6���'�F��2)S���8[8�(�qB�!UjV�����3+D[��ޔ���X�����\6'z�A���r��sVt	'�:o�X���H���	zY�I_+��fe@"喇d^�4 !�Y^@>	F�F�t��]�P���+�y�E��cv	8��������'���#���~�q�OEnB��E���L�k���4���Qx��7��bw�}?)�̚�0�v O��yM+�>.s�N�ph͖ѽ�����dzj����8Y7�a�m"#QpCZВ>���!��7�*��ܷ��C�,�P7���;n�T�"�Sy�{���ʢQM� ���GT_W�<�������f������=Q��z�ռc��P"|��iB��F���-���Ck�{R{�g�͕[�qEd����96������ˠ��'����[��pܡC��[ꌷ؉x�W8[��a*F̻ �=B���;��"����ҎC�
���<����<}d�l����g��	��9�e1{����U
��gd��� c�U��Xu`��l�L��p�Z�v��9��p�V���e���Ū���T(�(����'����7+�IL�5�tϺ�s����7�M��� �U��*����`��� u�/<^Jc��3o�jF/��2��k�0�N�za�J+'.15�`�nz7�w������	S�P �F�kK"�o�1���4���7gL�}��fw���D�)@�-�PY�9�B�O��>��`"9�q%��ʹt��h˯p�	)����'�J*�)�:q3:9��%X	j����¹�&/7Ң聧7�Q�F{qhX�r�?�  
�Iěl���LLxLH��5�^�~�RL��˙F�!6BI����uԺ\�A�xE�ÿ �m.�GW���8@|W8��p�.�h ���姀mh�@��G�T%�4��Z-���BSaSp��S��#D�*#�4Go?(3늼B$6Z�\�L���py�I4z��:�"�B�dR�c���b�G�;[����|��oP84<�xFu��~O�F<n:�����x�5Qw��b�X*!Y���qG���}���s��|+��#:���Ͻ��:m#b��%��9���⩆]���`?�Ύ���ie���Wf���d��G�X��j<�ʀ��e�͇~�|�B!;�'Uq�Yں����`���:,�2����@�����h.ʩ�-+�p�������E/ժt�%z�A?��`*���L�t&���������J���9�F3����U8��wK[��hB|p6�8�Ӄ��\h���)Io#>pU�Q�2�_K����9vn_4S�����xE�؉",Q"i@��W�w�z����f�Ķ�ZV��Mq�bgʋ.�ER��)Z��wKu��o�l�1O�v\��Xz^�r�B����'�WGGM t�T�*�1���.���O�ظ��׷���ͯ����{�7�`�������-v��fh�O+�V��������p�E]�|2�3��J���E/uǥ�or�g�3������Y���b,1X^c���8C������1Ɇ��u�W����vlN���T���t����Jt�>m�(�lh�1��N$�Z!�_g���7^��6z� ]��[�7�}�4�R7���:�l������#?��E���#m��>C.�vs"�/)�
�a��f�20MQ�[��Em�c6��G��(B�I;i3��R=(���ߌ�7د>n�m�(��&��v�7&��;�����S���� \��X�$��$1���B�"�w��_�1���9���mn>���w�c?��ͤs]7 �b�^{�˔�a)bY�E#���"Gs����[hz�''.#�dBmAϒE��p�q<*�F�_�_ߪ̰=0^�����9l���:~"�-��+�С����ם�j,�.�����S�����b����������^��{M��4E��ؾBF�vB��Z+���泥p�2�l�H�P*�^���"^��y�靎M�m> <�E��Q�I����tt#]��k��9�`�66���i�����<Wv�̽DW�	|	+1Lw7aE'��e�> �iu���[�Ȳ�ˤB�Ox�n��c�1*2Ob�m��5Y�Y���������ˤ~�r�6��'�ﳯ�I~7ZesJ��������ܔ����Z(C�z��@e�P_-��I�.�KY\27�h�& v�\�o4�£$�v�5N�q��+��h6Y� RSl�gm�X+�C�1~]F/���P���RR����ۨ�':�>&���W08�)u�p����s� �őcҮ��ؾ'g5fI~@A'm���.6ƍ��,�S��쁍�B�Ta
-�U�[�)�?��7b�#=�����W�p��O�������D��Wy�P�x%_��s��{�Q	ڋC��Y��n� qd�L�����'^:��7O��v[u���3�"Q�&gu�eo/e�� �9H��_U��-8S<�\Ĝ��gd������~��P�:�t���զ.5QhM��^�E[*���^h��񽽁0T�W}ɝ�/�����*v�؁����1+��J� ��dI�61���颻����~�P�zߐ�g2l-��:y]���W��"fW�cw�� ���ܓ��| wH��5h��#���C��ߊ/�($�x~��Ih�ɚ�Y��/������0�z,�˻k��%C�C5%nO�@�+��"U��81|uˠ�P�������BƢB���,B\�H��Id,��y1�l'f�%�񺝩ڽ���� 7�����ͥ�&�F�g�%�����Q�Y���I���> ,D���I��ܞL���뼗%_NטI� 9�0ñ�z���K�~�9��_3���]
�z��	� ^�>�����՘���".h���Km<�,�BG�sU����fjz,H���9΁��ݻή+Jw������c��-K2��a f�*�J\�ݔ�vk5��	��cYOM�J>��ޣ�uR�h�>��H:��m�7�Wh��C���}�ì}��5�c���tN�BzY�c3aV|�%�%�j�����N4:�����戵W_ӽ��u6|Z.�ʤ�g�㗂�\�TF���,t���</t0QW �M��/��mH� �"��j��tY�Њ�1�Аj	-��'p	����S��@bPTB��R��� W-	w;hfK���:[l ��5ņ�^�_���D.�Y��
;��M�� !��)�I��������!P�"�T��Ca�\#�g���A�#% j�o�����9���"<p�Bز����ȴk۹f<�_�7�҂g%k#�R)�%vA�R-1޲4͎PH����_3�P��.�����4�U:���t����9��8}Z �?�6�Ebeq y���i��viM��G^��f�%6��4�qd����j1�M�t岨;Yef���3	��2oo J�D�bm�h����.��m��`�9S����7�t�^AT�k���H$1�Ц�]]�mF�-x?��1v�=k�����y��NS][S�0� /��x���I�����m����'�d���~޿:/�}7�u�ey��y��l�޵*���b���І5Y�J�`�`3��UȦ���=>?�K�[���uy��]�U*Wլf%�y�D���#H��Wjy���R�DWpyX� 7��gN���}�0��n�AwJ�>�b�:x�O��`n�5p9��K3�z�z7������dy�}z�
��u���`wj澰"�������#~p�١��Ц�vq�n��	�ߞ�4����i��'�>�Ẏ6�Z#v"s\#�_a1�~��ܵs��5=c�g?#O^��x2�]g�><c�C*���n >R�V~K��fJGLZ�.@{t��h��|�(]�����lnQ Q�7��3,N�$����5wz3�ߨ*�1O�J��b]���e"1�~p����������@?֣(uU�2����@�%5��C������[P�ɘ��N$�gl)��Q�M�G��9�;�G�[�4"o�ԫF���������x\����#c��A��/�d2��mPk�a[��2�/��Mc���$vɲ����x��;.J(���R󀎞��%C��=�Z6�C�UxQ�ʘ�W��@�yEa��Q>멥�o���b�!�^L����ޜ8��G�Doz'�lg ,ZNT�|w��3᫕A��z�nF@�ٜ-��>v��zm�������,�8�c��X���;R��/ןH('�d]�Η�c�Qzf��CWFHu��du'�^�k��\�7tr��]p��*��NTO�E{D�Φ�YO����P̡�;�R"�u#�7���g�5N*���Tl��BOZ��ClQ�h���5
\��(�~q��e�p�YIx��L"
���l�}�٣~�sQ �=(����՟JH�O_xly�%ݘN��� ��3}�)�;�y܅]�mmu�Ҁ�/�J��~��j��5��P�i�a��h�JR��ɪ1Bw��kY� w�S��
3zx�	P���F��a�sVlh�(WQ:�Ƈr͊����fu�w�+]�9�����˥p�"�38K+/��R�'	�TL-0�������?ŏ�7��uq�|`�:�z�9���u���12�I����*�9e�χ��/���^�f�<��E`0S���x,���3DV.�Z[^�'�9�KΖ#Tym@�Cd@X��v�R�o���	x��b�z�
�Y@2���U� �p)JbĂ�H$xj,f1v�����xh5m�A=V.�*�PA9J0�Qa���`��<R��0;owԟc�U�͆6�q!���ͫ���M�%(+ư�ǹ.�u��w�Y}�@R5q����Gw�w����ݯ,�}&t�`Tƚ"`:�^@v�I��b����ᵋ�>�����P�WΕ�:�V���%�K�Ɂ��`���;n+��]�5��R��f)��L[#��� �I)���Mh���p���hj�l��l�P�Eh��$����n�2�MҜ��/J0LI��F{�$(��Z7�c�+ c�.\J�<��p���w�+�5a��g�&|~�ҵ�t̋ �e2/"_��ڭ�?���$�ی��$�Z; t���h�R�*�n7$��QŰ�C���y� ���\߬�:��O�C��'7�DZ�ߺ�O`��AU��9����3�t�,ȫ��s�y�|uH��c->��G_�r��Ie.�4 ��ۆ��M±� ����n�p�E��q��"�To��j�آ���፼zO;Q���! 7L��̓�ǵ�=m�[�,�,�é�~lӖq M���{�����r�P��-4hi�?��˳[��ߥ�
�	1� _A?�ڀ(8O��8�Ug�ynX"�]�9����F�=#��o��A:�{�!���Nʫ3,�{�h�1���Wgȝvq�<�'�'�"0s�Z.4{��]���a0)��{j��ܫv���W�,��;�|���i�:}��F�^�=�?�xU��mQ�P
o����0��o���Y�p?� o�aŜ���!�Fb��������b2��R��|�qtzt1�	����"Ж��o�#�=1`J�c�j]�:1���0[q�+z���;x".+�/K?����T	�p��3+f���%R�X��Z�����N�@u�����7�������^2aJ�L��Fo듈?5�nU���h|�T=��R�>��v�A��,�$��<��i�@��8���h �\Wq�ɍ���p.�f�Lp�4��u蝅�Q;.
+X��Ȍ���	�������&i�� ᵫ�!_'��{U������{[wz4���_v�҉�I >�U����3�C�����.Db�5:�ZW+�;�����3֔�	P�E���M�CZ%�1f�a\��)S#��@(A8��+�}@���t��^m/̻iMie��<����X�>�r��5 �CCLޑe��T5����vd�[��I�n�H�� �
� ��Q�w�I��W�dD ���6J ��8D˽Q{���e�&����D����?X<�h2�8*��7���t۟/�\�iח�$�mq+��u�0��>�h��˝��̣Q����T��9��izm�ˠ���C8���ԏU���EU��y�_R
�XP��F�^\z{����95�"�/�K6Nh�,�Dw(Jn����C���dWRMy`L-�0�~���'e⣋j�d<c��
54ݐ���f��8^UA�_���SP�sJ(G����=2��u���c���Q��-n��6Y�Sԥ�Q�V�ʰejG���V���]�.��?u�c��Y%9�%���������L^r��q��4�j>8��l؏^iM��y�,���e��ߵVLU���ȣZv��Ty!�1,����A�*G��Ȍ'&s.VPF��Cj����wG�}����-�����Cace��nJ�`�\䟶����nas[�O�w��zO�	�������c 1��KY��g0�����'�Dy|�K��w�.��
p�۬_�s��-�O84rች���c?[�����M�L��A��z)��a��2;�S8b�M��	�tƁ�޾����h�'���7��e�*�K�1�/Y�3D�Q�ik�-�[����F�7�R.�:P^��(�CW�����:0i]n�7�a|�(b���S��$\t6����SI��d	�ڭ�5"�tt�X��{6��=�:"&�Z��8E���e��)��%��w�v�4eZ���>�f�0���~G�o]��s��G���xhc�X3�#s���YP	-�C@��_��)u��gCI��x+�5�mGS����0����E~���A����T1�1�ƝF�%�|\͠ͽ*9�.�:y]z���N��2.g&
m"9�(�
��%S��h�
\��9*�N'�e�A䦧QB\���v��~����}-������!ê0�O��-�c�A�+^�5.��j�%��P�pGim�6���"Y�������|�L	��ٽ�#iS�d@r�/k	��'<uI�.���dH��*���K��J6h*�	�^�k�Ӟo U!l���s���T1K���>��t~�i���É�
�ξ�s��v�Ve۱�j�"s�[!�zm�ם����pEP�> �ѿc�y��7�g��gwȡ�	"Mr>��a�R�D����ڞ�[���SJ�M}�����G���QyĈGY"{SxM��(A���b���~�d�|�$u��=�l7����=�Z���K@�1$M��Ym����
7��a��~z����ٗUM�2εpUǨ��h�/K�qmmy�,��^&�մ�0�B!R5���`պ������X��u|A�z�]!��i���'[��4��r��Q�Lz�>!9zA���7��=����
%��٠���Q�%��+ ��I`)٭rM�Fnc�$��UW� ��Y{"kf�#\WP�a+w\��E�G'�Cl/��v!�6Ws�dw�#p��l.8�)��>�%�o�{s�;����cutq@
���D���)F�覊N��qe�)T@��ͧ�q_y�D~�#���}���N��ĨP�89Ȅ���ĉ'4z2�L�9��'Fb=�E6�f��c�fG|ݕ�!��V>l3�/RBk�U��%�A�;?�o�3��l��R�ˆ�~�}|#���!۬{+��k}S��)����gI�ԥQW�\{%�`��]����r#K3���h�.Y�P�07�]�Zj���SJ{�w�(�L�n��t�--��Rэ�>(A��#��_8q�����I?�A�xg��&���R�����?f!���&t%���=�~���yPq�5u��^L� u��E��c��~È�_�ԍY���SzS2�lX%�r6�d�%��>���'5_�Θ&�i/���*�wp��a�V�a��i�q�=��,%	����%,VU����N��hq����|6rT��[�U��4!�0.�Z�tmj3�'�ػ���>ƚQ�7a�*1��L����7]��v����'$�Pѝ(���ҔM�!e�(*cH��غ�촗��X�z!�P���/֯i2�=Pm�!�@ێ���_�s���W4 >��C�B�V-�Q�c�n���[1��F��kɇ��{K���;�!7N�@5���&��L?dD�:�v`�� ���E�oo�H����⚠W��F��O=���.��+���=XQ�����pW�}G&Sʅ����k0���k��V�6��"+���պ?�|A��6Ӌ�[��L��5&mP�~�F��3f#�	x��ǊR*���봦�oP㍹d��Xj*%�[��XD��trYLR����k��7�����}�����?	��g�F@@�0B��Do0S̙p�D�Jˮ��88|���������p���/B�'b��	��Orn�����¶5D�6��l�<����,7�J%,Ț=�U��*��S��*j_'T^�W�e��ݮ��7�:.�;<w�+`ga��"	
��S�0��Z���ԩ|����<��v���d��G�l���#�B�u]�T"�Z�W��[�Y�[Nk� ;�\���v;�cwv!G�/Y/��waH��3LN;�o�s?�u�����c @���a���W �؇��aUaC,���^֐�om�$���R�Q�|�WB Y�[:�W'Ѕ�&��N_�_s�� h)8J�d��������,�c���&�g����v�VV����0Ȱt�l �F�z\�+��uz��� ��W����CefqS�cj��k���ĲW˄esj1�@�!�Q���?�H��^�(�
�q�v�Q-�sL��*��R�3�m�%l�E��]l���O��T��,J	>h^�Sf�ׯz�,̈́֜�L[�Xj��\�lg�����XY]e�=�0h��lS�֊��%B�5az���맾~ʗ( ���_�<k�9�. h�UAc�D�F�g�E�=Y��R)�2X��s�*�IH���&aB(̖bC��!QƲS��e�BGX�KIE��R[S��A!��ơ���`�;o<�O���8��}sg 븈oQ;ӣN�%5���3�.s?��t7����+Q�=B}q�7�4δ��8��K8u��N�yxY~0s0p̋E�j�k|�3��Z�g�3�mޜ�+��4����|�XvQ��U�7?2I����,g J�2r��|@�	T���oS��laWW����s.�I�w�v� .e��k3Jn�X�ܹ^WC�����L����g\���9�lnd�v��ҏ�LDλ�xS������	�?��&��D�G��&k㵠��<G�y�Tne����t�������@��mf!��A��<��ݻ�|DU�c s����V�R�q��s*�q���� O�$��|yQ�_,�|�s���萸��tE���zo��S%X�N��9�����쟰�d������}!���0Ow�+P|��f��&�����OQ�'��%o�,�_���:��}t�a}�Fs��r�;и����X�r}Y��P���aku8���w���w�6�m<����vd[G|[�\3	��y�TA"S����Ӌ��J��M�4,#`uۧ"��ȉ�#V@�G#��`�(lE͢�k��g,��	{`k��U@�:�>�w��t�m:�Ӕ�_��#�N�N�&X�d�M�gNk���%��<�
ڨ�q2>�Л��̼E?cЭ�#y{4�)��R�Q���r'��)��޴"������]ָ+EXX��\S�.#�����U�4���3�~K�uy5IR+>��p����pJj�O�'�=�qyM��R�&uʍ�0cb���T�c�����";u{�������xc�;i��Na)�gM�%���"�S�򼠰Y���3�_��V��d�eU�9%K3��6Ԡ!����É,b�F|<jr(�=D����a�`Ƞ+��be�� ���8|�'��X$ێ��>z�vG���>3��;���X*#��������Y|.�sN����={r?@)}��1���X��R��t���b����h=8*���.tk�{�*�
8$�#��M1�.��о�ߖ��*���U1}�Ow����bVX����t?��-;��Q���e��P�@z�Y�u�%&�jQy�c����36��+V�@fCd�Ȫ^�{E����'�f_f����,��ER�#]�����P-�c��v$�wfs�$�+�G��gi6�]-���HS�QB?b]4m0���<:�_$!a,�腫���R�8
;,��M�S_ƴ����ś �o�8�{M-��\=��$q�wL?����)
tT��~k$�4Ǒ���I���t�& 1�;��ʛ��!���66���Q�th����R�A�A]ϵ�aj�2��[>/Ȯ�F���c����n�l�v7��;��T&�DRqYR	��`��>r'��Ru>*`�4~.�2q੽�b�XP�JA�,��i��j��4Z�a��l؋�:X� (ػa̱�t�	�>.�!/D�<� u, �<Qm��'���I�.S��H�,��aM�[K�gx5�Xx*�cAo������-Zҗ8�U'�D���3��f�#v}�݃Ì�$�f2��P�2ğ�J����݆M��ln�{#J���5j�t6���&i���S���i.ZUPǶR^�2�B��+����:n�!�=�ثb���s���jU�,������5�S,ݳg�.B����y~�jo.ǌv�z6u3��^
��R�-�~\�Γ	 ��Z{�2w0�}�7s��×pWp~�Q>�GM:�2���A�r1�8j����Q�_3��]����x_�K�b唗��n�8�o��Brڴ]T���`[uF�'I��g�L��9�':�L���a�.�J���p� &�8o]o >�4�m fqr��/lJ!��&�o#O��n�4�ΊS�d�|��9tj.�[���6?����������u�	�o���s2�h�*mC�r��ݝ{AV�5SN�[�'����9���X�e�D����6ҷ}��1#��+;Ʃs�ǖ|���h�0n�kg� s�S`.0@��L%��"���T�+"#��kJ��e��Ҳ����`��)Y�@�~��5B�a�v��4���E2�~+��dK<�M��
�/���\��]P�@�<�1�~=�b�Y^��G[��W����c���O�w���b��F�o8I���B-��Q�}?u$�fs�䒌�U�Yad�Z��,*��q&	��:z�ǲ,c�Wp�A^��k�^LI_���m* ��0��m�IІ_Ӆ5YC���X)|!Z%��w�����CP8c,�^rȆ�ׁ4˶�@���C����цޅ���WeC-��|����I��e���y�=E�F ���}C ���<�f��Tzm��1dMvey:���O��<�v��H��Z$Ȗ�z��Us����U�j��:�x��
���fK�{�j=�^UM�\b
��Dr}K���`�4+;w��17�r��hM��W��n`�H̙z��o-R��7���@�����S�����/&+r$�]�z���1�udk�4��qi��m:f�b�E�K���;�������mH���>����s��Y�>�%�QX!�>x�jF������%,��L��� �E����W��]�y�X@&�mB�U�Nk�u����~�3z�9�9��i(q4t&3��]���O0��X�Q�0	6bTw��v��PSJ��k��T姀x�ȹ	��k��b�n��5q���xZ�(���2��������e����"� �hX�X��%;�&��ô����CW��>z�t�>�h��V6�X��\2?�\�/�`@��Mk������1?_�J�^��������8�k��~fg��������;�K�$Rx�l�XU(x�70�?����/5� i!������W+���Kǘ�Q�"�޽�����W��qn���^Պ�Y����	��]&X��s������1����t��Z DG�a������#����BA���k�(��b��K/���J&Ǭپ-{�$�E��4&»�v� ��U|�[� �W6�a�9g7���ޠLl���k?ݨ�[TU���H�.���!2t0a�({�%8�͖{e�\�P����5�i�������K���g�Ä{��шș{�a�4;��9/*#�z���c�(���
WOY�S�+P?��+i�Ӆ:�ST�� ����a���s鑛��Y�["��Ə�,���Z'MD���t|�{E��g���d���D���)�~�(�1�zW��a�\h�1@S%ȃ�/��S�=D4�]�Z�0N�5$馃�PNoSVy�:���H��W��Pzo�����cɩ��ͷ�q�|:>�v�����YB\�8��g��;n@���g %t�NH�gs0�P�������`bg�����q%�@R'G/M�4+�� b�.R��ym&���zfQO7<(�v���ᯗ���:P�mL����,V����!Q��$��EAt#�	M�)fn����đL�O��lr��*4��^JqFo�H=�Y�}C�8wP�`��إ�$ﱤj�Ғt�2��K��ݨzd[I�dꑎo��}�n��O	'�����D� ��Rp>
5a�2������?1��]]� ����D��f���PlC�Q�&PؕZ:�Z�b��j���v�j*=mی�>�D�_�KH�w�:o�������b�ah��烠�[�_����W;��/�b%,�V��BH�"n;�EQ3�H�P-mB��䤥l-�}��V��.	M�cD��y�@�Wɞ�2 ���,H��^�$y���3���[ �,�u�6�9��k���$:x�l2�}k<4'{�H6����t�eE�Dܻ�/�̰C��=��@r6�S{�Z���[N�א'{�Z�%�H ���[!oO�G+���Ƴ��؅�/����7�n�h
��Kd��칱r�~0j��RVX�r���d��v�
�n=\�t_���76��V��t{v���,c�ê�,�i�\���>�+���F+�_b�m'|OԡS����PU�ϗ�;�1�tu�nP������|_���5-q9N�x�%�Z�""���͍X��1q���A33�_��DsWih��Ш�����I�[���Svaa��f��.�s��e���W��Ky����S���(���2�À,Fr����(���e��O̹
��]�)V`��Ʈl_h�g���d%��I�+n�&@�/a�	1�D�7F[�I�!�����ʽ1�,;iB��	a���s�ز�آ�����`(!����>�E�˩��:�0��! �5�0�ƫ�Q,(�r��ͱ��r�� �;r���-��2�<����P��Vx��1��.�5��C�h(EZ�̟��_�Ҏ�d��
I�~g̡�g��c�	�{c����q����o`�ژ���2�]5T��"��a�Zߚ镒:A�rrh47�MH�7�ބm1`M��H@����(ȭSь[�%������(*��\r��@�OҢ�2�,>:ƾX�)]�6QߏWh^�'�������v�]�Q��%M�R�mmF�x�Bգ���8o_�:F̬i#&��>����,�O������R�*��фCβ����|�����P��ѧ��PqmU�DȽ�/P�poFT Zk���+�@к��.�=)B����{۝��N�G
�pܓ.NѴ�x����3����ʇ�!ܪ���OMf��AqNt�{"��X޻�o����ܤ�?��	e��n>\ L�$�(6 ��Y�[,M����Q�W_��t����5�;,1��n衻F'�y�߲>X �D� �iԦ(ai�/^���� ���z���hH�J� rH9�{t`��e�R�*����F���������:�I�&9�mY���g� {�B{����ʰ��#?s��y�@��,����������nY�IdG������m[w���Hz7�����iTW�m����@F$Ѿ)OnQ�(Ak- k/��B�#�O�#lJgĸB�4[mI�6��a\����u,��Q�΋a�j���Mt��L�_n
��{�Z#��L_N�3W1r`Gxtq5��f>.*S��~)��$>Kz�E��Il&R�79��ƹ8ba�!>6�>��}x����SZj�w��:��%�O��aZ�Z�>p{(
��߯�;�"�RΔ|�m�+��H=��h#Ӷ?e����L ,S�uf�qN�G,�T6k������t#�%�+\��u��І�PӺ��1�N!7vp�H��zV�nQ�p2�2��~�����E(�[ܗ��"�dr�OČ��"��h��Rz=��s���=�[v0h�/C|�I5��-���.���0*�p��;�ܩ뜢�2�����B�R\?a�E��+UN���	2{g��,��5�ա��+]��pfVHi�ݴ�ʋ�d��r�غ6�Ҋ��f��\��/�F��_N�=4���v���:�p&�vE�G�y_42�,�:�xBd��>�g}r�'Xf���s͈!��A�lK�,�e�2H���F�b���k�D��b����v��i�%����R��E~�舤o�W��fG��p��.R���rL��|�Y� xE�a��'� .�˪s�Y%3�L�������	�!
Q���z`��o�efsvlg��?�ȥXg�%~���.� g:^xP#SOQ�$�a����k�H��v�28o@��r��`p�)xIzC��ͷ4~W+�3;�����ю]x��e��٘�f���d�wc��E��'t���Y��0 \�����c9���D�j��ˇ.&?���;é�ƛ�K�T�j���ds�E*�A8�~S�vmPt���_�%79��˸4�͑�������9�=���n�)��#��Jw�8����j?�b���dĴ؛������!���pU�����)���l�Ǘc�
���J���˛��of�|KDװb�PAE�윰�#�0�q���KhBgZ	a~;(��"�I�G�$n	%ˁ>.d�j�J��Q�(��R�uė]��E,A��{~}nE��w��S�����o��������"�N�m�g#�m����� �F�ac��l��i�J̬&�S�U��$/z�sc(X��Y����D�]{H�L���c��)/���5��ř� i�^H�@�o� ��ָ,&��_y6���	��bU�k�{M�'�<EBy�	�$ͩ���".��8�7�f�-(�L�3���!����
[�qq�M��+.���e��ZQ����a?V���K�����#+kf��xB^	�/&�E����[Η�8\�V�:ɣ�G�m�>�)}���):�t�ʇ����R0�n��Wv�qI��0�>쒑S6��-�{�ks�GpՒS�� ��k�ܬ��Ŕ=��xTkҷ=�.����F,�2�.C���)��vFww&e3i��(����G�bY$L&7��o9IRj�v�?m}ATJ�������	v9%���7�p���%��P��	=���Hmv@h�lЁ�?]hzmo�]AT^��]�\s��sސaEHf��q�_Q滳��U��(�����V�v�8�`\�h.�D%0����N���x�8��$t�}Ǹ�s)���3�V[���/]R�7L;��x�J����^�v�ˉ�{�M?�Mg�t׆u�y�V��/�4��4]�!㾞���p0�6��oՕ�Al�{�9�f/��������A� C�	�1��~�(��5Va~:0�.���Ǵ��"���Is$�����&�U���kO��ʪ�Z�p����KqE!«��r�9;G���ᛁI��H��)}LK	6 Ó�q�d��f�M�����!���)�f�-���魼�h�����y�q��񾛠��<�}���=3�F*�e���8�4!��Z����?���o�ԉ�)�W�-�\[q�����t��ZG�x<��$�g��p��.���e[���`_xg�X�"����W��q�B�$�Sgͯ������{��w~<��a�V:Ȼ�}6�۰�8R��0>�i7���=��!*��y�a�Z\>(�5�׽L���M.v��00��>#���k��R�$�8ʞ�GL�.K֩�Hʹ���֜���n�A�FhP�:��!�d+|��������V�ҭ����r��ԣ&]���z���ן&��N6��xl�䃗��3�8���٠c&�0>�I͍��>�A�0��g�pZ�\n��.�W�Lt	fG�ק%����! wwK�;��
�Mʲ؞�]�N5��	��ah\���?
��a[䐼�2m�7e�GcE]mg�p[*��=�9���W=���_�{y�[����WS�&�(R��vxx���{ӤH�����(#7��r�v[��P��?ԨZbk|"��=���R���#,�]P�1?���k0nwē�e��4t�Y]Y��������pR2f�:�m�)쑬5��*���2��'_ k^/{c o�/���l���Vz����s5��(~i��_q�웏��2Mp,7��\�e��ԭb���s����ԯ�,��Ec3�A��͌P�A[��J�����Uv��������,�B�.r&�	
6X�G�;�"��������@+�c��&x��3��|��*�t�\�\��<�J��biz0��������^v$_�9}&ڐT�e}�>]UH;�T��VC�X���
�Ʃ9)�q%�V!9`��.���>��ďB?���sc���x���Zv#��?({��D������w����|8��d��g���d���K�D_���h��E{����4T?Cef���˗��N���eG��a�:G���*4UXJ�����Ȝ@s(G�-�#�P�.ҺK��0&|���,Fyܙ�ynU��|������Y�p��*Z���|"���< ���ݩ/�������9���4�X
3ON/��X�\ɤ��>jl;;)��J���譎�l�o �T���n�7S#6>y#����֖�ڍ'��[(����iIT)��#2�����[ĸ>��1��+w�M]��I[Ν�����ESNqw�W� ��:�!�8Q=�$�8�xB�1	dŊ��m����^(�;�,!��{I�q�R�bnoĢ��n�߸��D���n�Bl��-m�x��w��J�^��0!��VK���[4���B����T���H�ZV�(�(�a�i�\8�<2.�Q�_g����y�,�0;�U�sN�u���{`*��q~�\��@�TL\\x�٩��)��8˳�E�J��Q�_�d"`�i�?���V��L{�!�o��'�j�"l|g��aM-�a�-�e�ew��q����@R�f�yw<��ܧ��!��O�,�� ����@��	���x���b)Я57>�\�Ţ�ŢI8�v�(㼤^��ڵ������>�ASj����ͩZMЪ-y��u��{�a{��8���o
q4��I�ȗGT|�ɲO��=�A�V�~D���\�#Z���J_�q�o{#�
�<h��ڍ��H�.vyo(�8擘$���E���@���;�#�ђ����d�de�Mq�8؄�eu�	�:_���ӟ@F�W�k��og�f]N�3����u413����i�p����w��M	���GZZ�~`�Fi���^e���!<U��������B�^��V�Rc�&
'n�w/�i����Z�5�x�x?䐧Q���E6��;��	{W��;[������L\�~�N@@��W���T�5�=��* �k'֤���� ��L�E�+�-��JM��_
MVU���z-t|7F9���%b� ���Yw+�v�{E�`~�Yk3y�wo�T^��{Լ�u�N��NԢ4��ޖ���n�>���+�tEG^��������hHS1U��4l�,D2K�uQr�ʂɬ�0����<d�e�@�G��87��h�#ĉƉ����NM�(���<p��?6��c�?!���P��Ȱ���>b���<�#�P~�B��J���*B�}L^|4�CN��\!d����)���� ɹ�:U�0�
T���F��A��Yu�P N	(�",���5���)�.��"3ͦ֐�ʞ6x��I���!�)�j��1�c���?�����>?U�t��j%Ҏ3Ww��a�_I��多�/�w��.n͙����;�N��F����H,Bof�gM �|b�W�Z}�M�iJ��Gx��������;�����o_��t��6k�6�����	�c��_��� f 0���[�x���F���d������W�l��g�yIa��i3c�_a�HH���?����f)�ΖjK'�_a~�;��Ƨ���L.6���֥�eG0��+QQ��*甼`��p��F��4�6 ��I�/�os��8����Q����f$c��M��jN�\���
{j�5�0�E���uX����`��g*�s�8�<�˛�of�v�����y���'�c�^���l�Ck����[g��p�;�n�R	-�O��TW�A"�q��R��_��p4��Q�Cά�%�AE*^7���������L�*6���E���}���Γ䂥�r�`i�4��(4��|��_� �A;�w����
lB)N�v�M�na��R�6P��iW��NE傶�K)��k���&Rr�@�cɊ@*����Ք�V?�b�1:�4��r�9�e��+�C�D=��L}eS�]��+�_͑�VcR�Q-`����@)�&�U2 ƜP.�I������1��3��f\���8��5^ʣ�`�%�e��],�MqA!
'���42K�|4{B[�UZ+��b&��������_ul�S�9��ݴ]��cnZJ#f0�C��������Ѧ��ۺ�A���
"Ő�N^����l�Y��I�N�j��Pd֋!}ag:���RW��I��x�V����e�
�~aɍ�ܨ�U�j��f:}0���GS#�81�Z�F��������Kצ���_q!���� 7�EWue<����v�d3�����+5�/*5!m\׃�uEw;�ԅ�����v�x6\����}D�#b6��j�p�� �{����:r�O��dR����C��7%b��
�	Ff���ΙTO¬�����jX�o�X�@*b�'���g�TC�/93��$�+I��?}�w*QipՎ"�C3� R*�wq�i��-�*�7�ZlW��N�n�B��xYO���َ'�yK���H��{\�㛼
=j����e��5�jf���2���`���v�^\�A�Ӎ'xZ��:ƒ��l"�Ү�Z��?c�+�٦RZlU��� ^�(�t_���aˇ���!ޔ$�GH��{=�V��(�9ܫ����h�=J���+��)�YvP9Fy@��9�eZ�4�Q
��M�_���/�ݪs_��@�id��w �i�)\���b�Q�hf���_��e�,L����_��>j/]#~V�n`M��`0��l9r���Ι�"�	!IL��x�4�$�U�=k��0�����8/�66��L�������6�5*�ul)_�m�+ � C
�X%�o#�r�O�OVRV��Z�u�n�m�8����F �t�W��V��dZ��+7\��%���<���6�A7�4��C:�[�=D�H�[��s�h�j��p��1���O���Q�D��|=!�z�
I<VE#�Y��~4;���I��RIF���i?��S]%B�W�F9{����u�$Ԁ�/���t�bT�j �<��э��XXb8�W�ci�̏u�cM�5�v�Z��S���o��<KB.�ק7c�����(��=�Y��X^��ʌ{�EG�X>�1����3��鬉�2�A�Q���sa�J�|�M����\Ҁ�Z��d�>��Z�4���W8��^��4�y��6���p�|�����|��pF��(� �xꆴ�����������14s�L]���I�O�n�޺�L`+�J���GI'�� ј�#d�B����H�ɀ�W��}����v�~�ɏ�(q���˞�a�v�t�-��]��m�8���_�w��!��$�����i�\��qp]��6C�1ɍf��M�������Jb3B6�j��f@�<�U|)�K�y�fL��@��K�n��T�������N�FN:��v�5�0��lO%�� "m�~��Yb+����w�] ГN�#�C����6R������O��)��}_��ClQM����>U�Q��8���0��Y�G�Xש�u���~�^i��l��L(���D%<��/���Q1��"o�h�j��|����ɿ�޽Vкne�5P���rP���F�^��iM�G�aZP�4N$d�y^�˴/�j��<��N���b�Ӌ*k����i�y�20�?�Dy&���;����~�Ƃ��[����'�fOR ��e���N�)8��:�b�:���r�%<"�D�]�U���c(-�7xs�k#��̄a��Z����
4�.��wI�x��`�R¥O�R�l��e9�_j�zx���G����p���;���P�i���S�T�B.�(����`�OdQ~���V&��zk��l���u�]<I34|���$��L�#�W�{�3w��q����Ɗ��!�`��'���|��Z}��;#�+yEk��L8���=x���,p���ݑT|w?�m�$�X���L�������l��Q��y�)؟Tm�ϚR�T|�W6��lϵ��yԸq�6\��2<!-�h��h!�CqV|SଈL�:�-E7����ݽ�Q�Ps��J�R����])\�\�a`����k��V�4�S�/���1�i��i�l}f]������$pS���.z����7χ�>���ȉ�f@gH]��}"Ec}����G��	����Ȑ{{!�vϘ#�=:��ȵaб��Ġ%���vd9�BϏTW���|��IBV1����{�[LDcc���*�qf4��5��H�?�y�0�9��������c}^��0wo��u�7EU���F}nR����7W8��;�_�U�	�(������ �]ׂ���X�����n���e��� ��qޑ�
�Y�X��#zO�O���?nOû���G}��N!�[�$�G<�8�z}���2��,E$��N!�n����s�f��0<0��[�|[�O�Ѳ��3֎�a��Q��y�k�(���$��&�MFs$J# �ϖ`�;�88�ƨ�GY݇֘k�X-wRRF��=g=��7�+�L�ߒ���	^���-��i��~��T
�O`ie-	,�ȹ���z=��� �[��[�Վ��q�ݝv{\��<���T�@�s'��9��LM������e��2/�KtZW��JbѼ{�����r%�B���F���%�~�Bd��,��]�&W� ����P�B"�>��b���nL���m�>���%�WZ�UH�nE�!X�?��E�~x#�3�g���+~1&Y�*�\9��྽����ƤԱ��ވ9I_6��aB�;#k�7��;0z�]�*+1��vd�7�� �/C�'��y$�{�y�U:�U�R�[I3T?a�d���,�$)�|Vg���DCn����cU(�%�_՞���z0�-빯*���d��� ���+8�y+�<�U��5_O3�-D�ILAԍ��*w�uY����)({�E�ܗ?�o�s��Ӊ����SC
(�x{��6���^����ɝ��a��)��>�]%4ҷ�9X�!dUS��rcP�����C�(�N(�R����FIZ�&����(m�|��ZT.�X/f�A��Ev1��|����ғ\d9� 8�{�
r��n��=<�/Sy=�H��(�r4��|&E=�.:Ld�=>�/��	#T뤓�:�O���R�ƔD��%�~��EbG�o�R���M��d���M��0�:�Gy1��(���kiJ|��rO�y��R�в�?h����'ط����m�)������n�#:�<��;�É�x��r�3:�b��h��#�J�K{����p��YQ߈8(A��3fP[uT4�KJ]�b؝�5�z�b��/^DꚘ%r[�J7�zz���\�� p�O����Z�m/w�����/e���?�r�<��g��{�鏣�{�U�X�w|2!X�3����n�uf�$��_��"!��S��f=_Wm�CjKda_�8AX�? ���G'p�A�5�+��Q���!�G�7�/����8�>0�����<F�ɛ���E���=}�H�a�R>H��7c��p��Oa�M��h4;O,/zO-�<�.Y(��C�vm,E�΂=��'�\��s��)ƈO#>2�]�b����X����3 �D�����|���kx��j]�z��N]�BSp����[��)䓙���e�w�Z��1,�o�/EANv�D〉�8�Bp��ShC��A�S@���p�����FL�{���'�~Mr�����JG�����4Ra�&�\���w(/�!Q����!��Esh�| ����N�S!�۫����~B@��W�-��qq�9�*i����Q�m��PN�+�I����߸���3�bV�M�xa�p�yߩ	�Nb��KO?�Pzk4�S�ϱ�R����2	�Rq���wb�.6H�]�wJ�'�6���T�ã*�3�R�����}bc�U�60Y�ل29b���7��(�����&jJP�?E��=C%�Pׯ���&j9Bd��o]A��X��u��(h	�Ȼ�bh3{��^��6O����w�g�G���B����_h��`g�Of�ѡ«�����0�����}����2s��wV�/�36L�޶e�a��M���:>� �x�G�6�����~�gE�a�ꤪf�z�x	j���d<����I���3W��,)�(sb�jށ,iy|���r����Ed�zkg��ɇ_��A���t�p���â�|��u���S���Ԙ�-r	�C�rCM/��\@��Q��0>��Q�ؔ+����A0Ir$�6@^�R��a|	j�v�N��?jo�dCP%�%i!��cb`y�#�r�
����$�̇ �s4ԿY� |F�9��{ߖV%:�y����bf��.�fl/!�G�����2Ғ�LȊ�D����}^�n���تҮ`���T8�b�z�?j1@�fh��O�^�8��5�,t��>]��Zݐ�(���ڑ\��+����Bq����P�2_�&�o4��W34���m��X�bn��X�^4
��Gp�itD�ق����Uy��4vt��E q@���bUf �8�du��HJ�)_�+hb�����!?5FI./��催��9�匫b=TN�bas��ʏ��)��E�FϷ6!o5�"�M��������_}A�6I�
�nӼT��[k*M3+�w=
H�\��R�횺�f�&�j ��"�0|���`�@e�eWjtϱ'e7��Ry����p9����P�m3�M�ۃa��C �XQ�{P��΋�E��׾B�w�%��Ȥ�l�-����YN4W�.2)m�`uWi]�	�pO������������(2��6���9r��7�!���9 r�/�;��L�)>�?�K�������nD�G�f��z
)�因��������┖�|��H��-pG|c� �+Oz��^�������n(=)F�9 �Z����c"�}:��QO���BR9�#F�'����MŔQ��)m�k@qa�����[j:r�� p@!%����U��{�*�w�1���L?QE��3��	qov.�iUA�d8o�`Nꖡ
}>�7?&���ҩFt��� �V�:��pkr�m`��k�`9[��2yێff���+�!�-��6<����C�=D>��vdſ6��8+� n���;�/������;�Hz+ST)�ä��$�]�c�Q�Ҵ]�È��S��*E�S|��T�y�R�f��l����@śe�6��W1-=�����Dc{��K!���gk�!�g�?�1_D�FM��h�~��wu���������RI��N�y�����i��Y�E��)�⹛�����yФ41����~�'�7�����7�qb٤��*"������k�Zz���E���.k�ڧm��v5l��"����o�C��Nq�0Ȝ�`��DE���#��I��@��l'|�����b%i-�웍�P������ob��^�AJ�cY�yeh�n's�><�c�@�V�̆�<K���)���>�Q4��)�3j��8�V�C�#�����.ig_�|A<�\�����nne����d��!��aD��M�|�Hp���iQF�E�' }`�5����O���>hb��,ǟ}��/x��b�C^���dK" �m/ݽeC��CV��!B��#k�)@��~V��	q�����u�����_��ۈ��=9�|=��<BZ�öֳ<5CW�J<f��>m����dGy(�h�N0gZϸ{��Y�C�=/���[qt��3�!�,�~�����
P�5�5!�xG�$L3�3dXg{)���¸�c�I_W v�p�`��I�� �*;�	�����/.�.%;�6��[,��uS\���`3�>-�D@��C�7�S7 3â�#�^�o�'̊r7���F5pr: O��O�=� ��}�����q�����}�~J���j�iR�~��GQW�@ .p� �'__�.A�_�k��4��ٛ
s���rV\}O}�dzv�-�°q1�M���'w�Ŀ��Һ�xgf�9ge5ߥ�T�҃�7�������CQX%砰��8��hlތ�f�5� �w=P���U��:Sc^O��xQ�"��wV��h����W������`�<�V��<�h����q�İ�AΘ�kC(fS�K���Ev`�B1�e�������+w�e�s�h�t�Y-�-g"��g�n��*P���w���C����*P4�6�H*;t��ˁ���!.G�#��G0!����#;l@�=^n��e��m���o+�!��x�g֝n�rd��U��-���2Q@=�b�ߒ���跟�+B�Z�f�N�{�j^~���X�3� ����+og[�jQ7����)���w��k'���MNěǤ�VP��@��*���Fp<%P
-�:���&���<%�+��GV���|!�2�_:�x�&��2wt�-��\k�.<(�ÏA�y ���EV=�g��"p4A`������ŀ:o䄇���O	�İ�(�h6s&ߞw��?N�=��%@GgF~
rl�Ku��ǈ4� ���988������V9s9�ړF���C�jw��7����L0�SZk��Y��T<�tW��F�cW3���=�ylz����VJ�ǽwg��`��`�(�i�~_�f�=�d�ydĺ#t�Ҫ�$G�@�Z�/�{$�q��i� f��CͶ�<B�<�O��3n5��lPXk��t�h�8@�.#�4�|\%T�]�h1�5�q	f�12K�܋��I�㧟"}hý����-��b�o�6� ���z��&Bn]�f�67�;����G�^?^]��;�i�|6��_1M_����`#^o�͐Cl\�αf�2��TM���)#UD���<r��},�UO��'\[~��9�����(FV�W[]��B���uZ\=Pj�&6��_[+Z�zr|&���)�W�� ��q"J	Mu���AS<*��h�0��Ej���k���B�Q1r�u E
/S�w�&��yu86�j�KX7�Xy�P:d���2*�
;^�2��ie۽П�L �p�+hQl�w��ݮ����k-9@-�����|p��/�G���9�	��zP�E6���i�O�
w�� y>�u�	�%�
bsDcWY
gg��>F�8�RԒ��Ծ��[&b$�na<�|e�W�S3�����j\@9���5	��\r�&�<��֟����]|~Z-����n��Iзa`�ޞy�a��,�x��`t�{��O����YKDb�^:����x���\T������-]´K^�fX6�,�o!氞���x��19}: ���e��^;G��V�8����?@���+�՟����Lf-t�7`%��_}_P]�t�mAz�ڡ�~Xm`+�:Ⱦ8%_����AhH��A����^
K�V��n�@��@X,�ٶ�-ț�oa��_�cyvт��*�4�����Z������'p*29�,�sf�F1A���(5~��p����"yx��)st{�h6�dT�[S��e��ڃ��"��k���5��/��ǌwL������|//�E�u�@�E�҅��l��hC5%��e�p~�.����;��<f�3nٜ��IG��i)g9�v���N��(��
��AJ
pnp9Z�^~?���3�8�zI,�9b_8���%U��Q0�Jღ�iv�/gČˌ�,�6R����M���,�6�h�cE�Y2�7�Oʾ�/�ʓ��g�W*�Y���ӏ�8`f�E��Tm��K�/��aHXugpa�mZ���g(�/6A�A�j;�/Ҵt�S����4�?ڒB�7�$����f��-�A�t�$�$��R��zY���J��0�����	�{L�Ik|�"�K��r�.��!��WA����T|$ J��>�j��������ͻ��'X�ﵒ|���
���ե2^�_�M/�p�^^X`���#s$-�l�F=���t��|P��B��W�mqa��8P�M�j �-�U��N����Bگ4���~�dxBn��do&�ū��f�ww	��d�"c�D�ݳ?��-Ll��#��\�\H<��Ym�]��]fÒ��4슖v`˺$bD ��0�v�h9�K4�w�-�S:(�Y���1#k �䢷�U�l� Q���մ��R�B�e��׈�n�:*�қ�L[��v��J���Jk#ݒ%�4׌���������5t�дX��0ޣJ �P��e��HX��K��t��>+�B�	�`�bz����;s|G�
�g����P�����R'LV�?����25 eW]�×� Pq�ʞ�Qb�Y1�O�:��tL,0�
`��)`��N��?�{`\�Nk\q���w^N���:�]I��󢦰���	�;�M�L��/\#��a$N����l�!\s[��#�Άޯ�'��s�a%�\�5Dg&�[�W�i�	���x�<���bK���FΔ�����>��R��Ǩߙp��:d���a����bJ�KyKMuX����l���t���3l�GB�-XRd�P�V�"Tqh��ȷ�6��=�!)L}��8Z�x����	����Zg�3/�n"<��)ZU�\�8�$p��uR�ey&F3>�6��!T�����m�X*�9qEY:�g����5��6�Ķ1�u��|=&�T�H[���� \��4R��l�����P�2��j�i�9
[wŉ���+��;����r�p�R,�Cb��Q{� ��\z������9???�9�M~��L�(%��>x+�l��υt�����\�*<����p(�U�S��ͷ�����~�����^���n��`�T�y�c�,Ɖ��ꬨ�[h/]��s@!����D�4���p]�8Q�K��P"���/h�����LN"��)$�eF3<��ZR=$ӝODAI['��P7K�A�D��	�Y߿��d^���������T�7�.����L�)z$����Y��̍FeF��Ɠf�
-�hP���f�Z�BE���>�S��&&F)�,J�,��qh����@��䯄���0\�4t��52��@�.�w��o:�y ��Z��~?[�.CԳ�������յ� �u�Gj��O�%^qa)�g��a޷oX�N���$V.�����7����P�
�������2����y]Z�������aO�r��.^�����.c�ǌb�q�hU��,Q�{�6yѹ�^x�x��VSDwg�dm=��t���"�>�ؿ.~7OK(��S����j����Y:o��2U1�Sݎ6�3脍sv9w�"���E`��� ;8ƌ�y�<��<�+�L�Eܡ�0
�N����&l9������9��w�׏ݧ�J6ޙ<�]�c�i�F��>����Sc9�;0���5?e��?qB|����������g3�W--��-fk4��������X?�w��OR5f/�2r�^!��O���!������9�T�Œ�./��_5*���<�0��{Ff�s%��"� y�99��ul�|^d�y��{����b%��Z܎
R�^��G:��&�D{����q�����\���ٝj�IoGRD]yKr��[���K����Ñ���������3�%�y~�:,˪������G�U��M�uㆡ�2�m�m��)m��8�B��KS��'E�pg@�-�
�y��*`7x4Y�ܑ
�*'�Y�!pi���R��
M��{$MM�&#|�i?�����?`�=�%���fG�-1���u���>b�=�'��g�L��K@@{�r�Cĭ��Ͱ76 �x&{�A���՝N4���ur�I�,f���Q�-<R\A�r�
K6���+��9�V�s�ޕJn4���j�9ql�$׿DF��)�����&�p��O�]�H\��/�c�J���+8sr�6K$��{�~�9�OJܞ��RG�Rwp�ΕB�	;�C)	���mWPð��I���H�X�/�Bn�,�|��@+�Ӡ~�_�j�Œ-�N���?�*� ��poL]�{�<��UhV$p�\ߠ�FL��C@7FE2���cT����tl���W�4��=�a�Tϓ���BR8���L��;�Ô`��md,l���wtĥ\<�(i���ڊ�hF�Tg�����Â�X��+� @gY|�eK�k���`���f{�"��h���P-��p������<}��p�z4[*Z�]A��ϫ����B��?D���O��2K����M��Dv�]�p�z&Z-���1��[Z�M6�	?��oNh2`�W���9Q�}G�(�l�c�����*�L��[��T\AЄ��[G89�����?%�pV�E�/x�5���9��/�H�>ܥ����@����2��bn;	�%_e���8�{��4^�E��qqYܱG͔���n�S�B�|!��
�a���à�?�#���'G>?,5�.�rӵq�h��DYp���G/�|^�t6�Єs�����v��(��ǓΌ[*c29���<K'T�La�.13w8���K�&�R���=�@!�V�(�Oٳ�����b~F.�H�Y1߱7�Xm�:G3Q�!U
$C8T{K?!�=Hł޺MSeϴ��N�w��'��W�~�H�ɴ�=�_�*�ٹI��"�2����)c��Y����JD{�Ɖ[��ߺ��׷
PsN����XM��Qf�&g1CJӭ�6#ں,���@��������PV�*���Mh�+Y���B����R�S2w�U�v�g$V�B�,&�b�+���ORl��i�|�o����g5;����`Bln�!���NbL��,�ė�A�B���1�� _va����b�a�ʜp݅��M8�M����t�.����h��7�Ε��b�uX��i�(���0�������s��-X����K g)��\���tvB�U���:����?�^��!M��NpQD�TK7W��(U�4ciɦ|�Xw%����8�oT�y�̰�y$K�h���ܡfJ���2����9k�ث2��������F8��l���O2�"lɒ�/H�� y0�j��U9�/ V�Pm�-�f��!�z9�`1���~q�R��w��@s�x5�Ĝ?���ShKj���P\��� ��]���0�5UпQ�B\�9�����	����M֜TRwXG�l#�O���1|���e��;F����$Q����Kޮ/��}�z%	����RT4u���WMO�}��#�74�?�,�	,��A�W"�>ER�e��WZ��d%����W��rՌ�j�W �Uͪ����Mg��v�Ʋպ�M�&�v�~,����V6 '��8�g�S�~a%�B�A߾Sn����:�A��0^Ts�;��o� ^d0g� v[�z���:��g�އ{�*�0K�J1����l�H.�+HE�1�;`���ʳ�P�E[]� O�4-�b��KַuU?<(���kLc���%Dlf:	=� �t�jv���j�г-'<��\��#�p`�tl|�҂�B�6׍���Vh���G�Ab	�B�v�`�
��֨b��?�\6�B���J��'lh՛�%�N�v$�0�IԒ�7����?���`��9����d~�
��>��	�F��PMK�s��!�)#��)��/~S*�F�r(��=��S[Rk�Y��}��|�g���y����Nȡ������s<��i��$v�B��}�n��7/��%M��wyh8��!f��&p�/�Xg?��?eRd�"��f����Gp�	��w}P�e��)i!��'-O��>m�5�n�,Z饷�T�y�H-���E3tc�-�th��S�:O�u�#%։�]�~��L���~d�^Lc+̞���-�SY#>���戀l��V) 0���4�jQֶ�2л,��Y��a�:���&���ȡu:���^'F�ʬ_����n�ˢn`ߒF��h��Q$�\X�E��7�#�e?�xkj�Zs��!���|D]&(�������	O�
�Ax����JI1Tn�`6@��j��z�G×^��)H����	(J���U��{z-f#ߦz��.+�����%��X���x����\F���*/����"�Cm�d�����%����ܢ�r4M�g�����������֒J%���NJ�����j��{N�ё���I��`5���?2����"xLLF�E�� S'{hh]����w�[�>���W�������4�t����,�>�U����R���V+]1�f#��i�#!��:8��I�6�ǞA@yZ�`��3���ˉ5�#�嵮�-́�u�f�#".�@�*�-.���^�9�A���XG�L8$����Q�v�#�>`�e��v��U��P�wN�-Y%�]�s�}b>�L��`����x�j*�M]��W�����V�����FO���Cd	�>�&f/"@ɉ|w�������cۦ��B��l�?���+oW_$�EUD�<;(��\~������<�#VA$i{��Bd="+��ק��f	Ӥbj��x/i��'�6���Cϐ�&�񷝎��G�X�y���B���5��K�-R ���DA.@��(��-e�˫�p�YlB��R�H~`�n�W
D/`�H�b%�r�V���ii��
�����8M.���	ef%�^��|���p]��Ǭ^G$��˗��"X�%�²�u�����G�ՠ; 8��DZ�+\�;��������cm%�w/�u�%�hX��At��h�����)��a�e�GL���Pb:��OW,&��iK6��z��M'�GE$�;'�U�!�a�s����Fc0�����`�XRl�P:c�0ԌV@���?�a^й�e��2�i���å1:���P<����"m��)����ϙ�g�h�qظ�a� !1��+�yX���pU��il�A�-QR�l"d��w����}Q�3�K�j!+�ހJ�on��Z̝eK&���v�L�Z}����[u�:��U�EEa�]���ǔ��=��PD�٩B�f�<�����O���H�XI���-[.i�O_�Rw1]g��ij�{��D����ڃ�$�7�bI��d4e�e���v�33�������&Iv��9��Ni����`��z�y�lg��*�)_<�<x���k�N૭&��pN4iNN]V��Q:�ZG�`B�x?!ԌL;$�c�Jk7Ei��@ձ4g
���o�y�ÇVʥ�5����)QhM�0J�b����or���L؜�資g,b@�M�+1WY�"2�:�ײ�~)���6n+: �>6y�	�ڈ�Xb8U3#}y�փ��3Ǎ��Z�O�xg�e|�:E:�߶�ͷ�(U�4(�N��U�bQiW�v�נ߬m�{v?�C��UT�sǼ�Hy�(���p��P*��ʚ�r�0��ޘ�K�e��45�ղ�vk�Կ޷�]M&��n!;�:WXV���sr�W�e0���U-?�Mή|��O�l�Ӧ_��WVUV��	�PQia��(��~��E�4m��i�<�=j�!�^��<=���N�(g�pQAKR"2�?�'����Q;R�<����Ѓ�ßރ�o&�oC���M��¥�T���yA~��~Z��0a7���#�Ķ��խ�	'�a�MQA�@.$nY�h��KI���.�O��;qܝ����̚�᪆B���J.��0���f�rHGR�t�l���O����S��BR�&�/U� �p�/zxf����4pE}����\��\YA����?4ǘ�9�����O�ĳ��f�'�Os�_�R�$;��J��H?�l����d���H��N4g;N�C�S��EŔ6Jl1���x��e}�m\yjZ/Q8��� M����zԲ߁k7$��#,k���2���ٹw{Y�w����X���FRX<@>ӄ��+a(����V*��5� ��~U� �l�B��1������F��sW������Н�Ÿ�`���2�A�K\�ڐ�~�e���%8�R$�O��XVeb�Q��՝B�`wO�1J#�R�T�O�A NMnqxYz6�{x�¯�u@��nO��Qz	=��Cc��u��3��2p-@y�*�u6,��.o��'���������}�>,t�!B"7�݄Eq�Ɖ��F�ms2��87=�\|JY���81�՗z�M�'�T`Ȋo��z��>p3;/Q��4���gOUk��!b��\�w��Udm����e�rӜ��8��J;2��ӥ�-.�㰐�o� 3�*ɚ�@�*=ya��[?<������\��Q����C{OlA<������=�<f�]�z:V^�؁�p��+��Jݬ���S΅tp���{�0��*�Ak��x�'��$�]n�5��ޠ��#SlE�(^e��t�r��7u8pU��RbP*&y�)k�~�HM t�4	��0s�d0�ӻ�ܞ�b`}����%4s�`Z�L�����R:@z%��86m_�(p����T��}i�z�wӉ"�ICwF�Ľ�LZ�_��I��D�v��w3Uk���y��a�h�惻��hs*�/��ѽ��V��2�ɕ�=�L����a+�c����B."��QV�~<Yi��]�%�dj0�!c����'���0�aG��A������
&J��"���|^([�7Pc�?�O��7jQ�\$E�8'a.-�42#-ː}�7�J�s/omذ��v���l!M��J�{Rٯ��(� !a@��y���k�2`xK�*�J"��U��ء�^���&?0Ft>J�;��8&l��K�
�m|�,�����Y���lM6��0�^�]��b/㭝�ޭR#o����U��w�0�g;��X��r֬�@���= �Kپ�%���Z7�ҕ<��|���,��3	%M�3|}�I��U��"-;����	-'4٪��G'�9lۆ������n8HSp�3<~�o@1���G-���\.�~���������X�3}.j�7�UQ�P��+34�a� Ҽ������\�C���/���M%K	08�EQ�8ȑt�q��!JnP`a��ۯ�Gr`I��r-�ŉ�yn�L�ϥ�$�zM[`�Γ^^��x��HW�������s�Z0Bj�a�l��m�3 �˵W<r���_%��6���;�/��~.�j�q�έ<�S3Tj���	ͨKְ#q�?%-�(�j���R����!m�H`:f˧���\�KD����x�/H�쌵�Ԁ�4���ؤ�������5yN�=*pd�	S4�(���t@��{�� -@��ù�dc2L�\�5%�N�%����@�E�W�z�뾲\��^��@�AR�A�~M�%��	1��R�H�v֣� �cf��U45�#s�֖-)tniOcj�������\1�����0�m,@ w�&Z�������R�7��=�l֚}��:�@Y�⯴�4�X�'�����?t� ���.aЯN�� �:�$u�%֫\�COႪ�4����ˢ�-��&H��}�(gx����R���D�J���5��{���.��y�c'�@Rk�!1�	����*�����.�;P���QoP�x��s���LT��u��Ki�W1���` ��Dz��Af`����6�齎�� 8R�-b��%&�w�y�4�a�Z6��k3X� MMXܱ`,��"<˕D��:t�7��(;�q�X5�L���V:(em���4��S���lH%��	nk3�i���N�#Im�D%��{���葛�4x��f�c�@��!��HJf�,1��0��Z���#HK���,��C��C��7�+�K9��Et���F��3�g�ح�aW�͊2mqT�����Q�mY�D�c�$���M�'FCi�0Hk5|�h�T:j▌N�����fl�*�T�:
)=H*���(���[^��kG��P�2���mI^ap{װ�����v��@��
��ЧL����8:��:�]������}�wy����P���~��V�HF��
�����fCҭg(��k��}�>�P{���2'Df�����͇Q���(� f��&���E�#��pr� 5��{���[���q�n��vFN�7�a=Y�Y�����'�I�r-+']�ׇ��������2��Bx>�Rh�A,[`��=O4��J��O�g�E�Ϋ��?=٭1$�ё�^<�j 	�Kz�O���&���qIn�ʍrq��gg�l�s��4U6���m���HP���N�����L�,�'9��E�&��&�օ0�MoR}o�~���Ee��(��Ǳhr��]Ȟ�B�#��mk �C%vX���EO't�`���8�1{�����S�}�tw�~*�M�<$ijp��+m�H4��"�ќ�h�׶�f0����R�SFc*8=��ؐ#�we�N�D�L��M������s`W�{5$�PL��W�g��,��hu��;��cN_M���qdC�7���x��vm3�ȧ�V��ȼ�~����l#ItC �ڷ�B���-Nn��RK�2�uv��gU4���x��:t���(�-	��sf�{]B�����Nmf�&�`K//��'1Q�G��yd=锔�J�0z#����d�ZNDP�XĿ����'H�𖤕h�ڌ!ܝ�|�?������m[����^�\�����iۇ���\�cN�kر�4�D_�t@�En��d'�%%{,�ܻk����T�N�������V���[�ҵsN���e��|�R�˰�miڠ��!<��DL���l2Bfu��?1b�6קП�U˲;}6��X`_^ΓG���@$��OO[x���+���Ů
cd�E�����4�5f-D���D ��9 �ącH��x^j�(�B�go�9E�C��U�!��
������v5-ř���dD��R��J��kz�!�~>[RD7a���o�W�^����|��C�y��q
��Z�M��;=~%�CЅ�LB��*{�zz	�
�O1�p���#s�I.��r�5iL��)�j���xo��$r@��s��2�Qꕹ1;�E)�'������x�o�?m��ɏR\�~M�4?6	�B>~�o�cMP�p�_�>a�ȋ�7����~���+��$� {��>��
����k�R�5��ױ}
t�\��96z3�ǳ�ދ�՟Ek��LH�n0R����Z�0`�[I[}ɖ���o�d3a�K����0�`XZ6�$����Z�w�z���ox��f6@�E+%�����y���,�_�-��ƃ�U䆣W�!���[H>��*f���ʡ��-�+��s��ԁK̧��������ʝ���p�NH/�� ��Z��ɧu�E;��?�-c�|����wu��.M�Q��9�F1�+잊��f�����V�NI7��
*����靱�~�ou��x�+���jK'��8I����+���6_b]�g����8�~VШ�Ϩ�D����v����/�pVҟ�ˍ�G��"�}�2��s��?0u>���ڰP�I2�aq�L����9^7~�}6�=E2k������Ga��ɹ�p�4r c?�]ߴ[�+R|˲
��>�Y��� )|uŐ�#���ڳ�8��f��W��J]����o(�{#~�L�(Ie�֐?q|6H��9�f\�3����c�#�&+@"�?����=�ImkTZ�
( �Ǝ:�z;�䀚�r�}�=���|�/������Q'$wjK����>�W�w��[X���P��Wφ~O�x��m�~�K�R�Y3?1�w:��m�=�c2&)_��u�A�� Y0B7q��K�����'�hX��t�����C\��u���w�m����<�^��!eS��[r�^�֙����$���������l�����z}C�_.ƀ#��KT������X9�4�+����)5N��n^$@��s�>�N��	w *h��xw�-s�} "b�(;ry��BiIL�M���m )~m��ϊcz��M'"T	�"����U�$��8@l�r:���I5��[����-��/���I#�����=�� _8~�.տH�A������?�+i�u��<s���{��F�� 9�p�I8m��k��dK����gm�O#���8�F�P,{;z��c'`����x.��63o��6�r
�L_ʇe��M����f}:�K�
9!�8X$����0��L_"ᓷ�=�,x�X�u[�s1ih���l��t"a�.;�Ϯʫ�Hi:��u�����ć|�M^�լB{��.�R~g�q���a��Od�!a��v�q[��D	z��y9��a#E$��8О�?�'j��oj6R�ۈ�C5�*��y�x���q�����\�2��#�Y�3{o��f��-�{IEC��^ #v�#�_�pd����b�������v9�ן�D
XD^�4M,�xt������ڕ\T:��T
Ū�g��YV�x'ֆl+��V�A�D�'��h�?l3�ĄJn}�CԸ"V5@�D^���AL�����Op5�ą�
�A+�6 8�Ԁ��@�b��f
�1��z�8
���|�x���B��Y��>R`[�a�o�rn9&�hc0�ɓ��3
�L�VI-
}ly�æ��CBVD������ �k�Z�[�3�����]�^���s���$9�͙����S��;]�����}�+��@F��=��y=��h��9�í�:��4\ͅ�AE�_������ pиaN�& i�G�BM�q���ssh'
 H�(������9��=��5���]�~j�B�=��I���ۄ Y�� DU&�^���}�>/EH/�����⅝��J�Q�'7����*����;�G��M'v	4�Fh���Kܠ��n��G{��	N��9��o�X��Bރׯ4���θ�л�������q�	W�n"Ŵ�o����Y�3.Zle�;iĠ6��ۇ8:M�]B�����ZT�jV�(,�DQ��_1��EN�jyZ�U�	?��x1��0pm�S���AR�=��}t������Aȼ��JΎ�j�hb�rò �A�"�Ǹp��@�D�=W�P��������(��~Z�G��� ��E�0r�`YF-������4�!51a��cF-1� �'EI�dq��ù�L�v�N��i�.;|�e����[
l�I��h����q�7�ேL�;�}�b>x�7��چ/����wZJ��G�,y6�v}��=�a���#����{w0��1�5��E�@��-]�[�����|1��K�qĆ�9s5�ڝY����Bn�V��ҰI	��A֤6��� OA>���G���܉��g��."�/�}g�q���=樐Sv����57?�NSƨ:,�ʦw���т�� ��� ��H�� %�$u���-g�e�n8�쥄_��q/���̒�㴾�:�Mj4��s~ ���b�[J��m"�&,e��i�ɛ�99�;uQ0��O���3~�OS�\y���8�i>8�T��
���˹(NE.Y�DK���M+����n2Ǜ
��+�3�ʮP=�\�'M�[�������"q�u��PhhЊ�0�m<dl1|�v2�>=��S�����,����q��}$�/�Ӕ��f�xpʩnD��
q���;��+n�?��*@S�ȉ,�9-@{�2;g����(��+h�t��ES����M{o��SK��0��)��k�a��ц�M��2�
E��ĩd�Y��"��5j�\t����,Δ�Լ�w�7�ۙ=�fuTOY����<	3'��]��k���(�z��I�ԴӰ��߉�8���:�Y*�`�=�������X6Ne~)�%,Z ]NU�v.���ر��ms��6�.T��t�����ٔ�h�!0�C�~�>����s��d�.��I�o��Ԋ��:�Oe�Ąe��X2���PA��񂆡����Z�0k.�����.�C@��$&�J�P�+y��g�K���!gD-������S�$FU��¬#�|
�����W�����q�������F:h*@��ڪ���X��û\H�j��cu<S�,��z.%Y��"�n*� �\�McK<R�(u���D���$[����1��=[)�����e��zwŠ�q`���&��*����SUN�s������8�e���3<r�*������d�����G�R�0 ��]�&%I�?�U�����y���ʸz�-&K߃g�m �ƛ�'��D� FסQrk��*@�F�`8�ep�5@�̵�����HR$��P�҃���R|\֥�d��<*?���S�\�r�n����<��1�ѕz.�1���z^ɇ�`^:en��/.�Mj��3�2d����#c< ���� ��(�2�+-HSzvUz�a"�$���� n�>��Е��m.% t�au��O���W����س+�2>��0U�GW���q�l��t����@	�W�d��h�?�iJ�L<�����?���NT+��?�#��Ϧ��c����8˽Ӟ�}��b-Z��0�'��_�.��<��V�E7�S\�2й�q��VP�ߛ�#]�fWA����B��d �2�0����f��6�2�m��OM��2@ �L���3i_M�d�-I�?,�Zc5v���~!l��5�L��t+t	A]������� �%����(��D���W���yܪ"�}�q5N!�Up��B.��>]y�y0��]TPI�=���=j]�K4�ԍyo���h�շ*m�z�p���Iw�[0խU����Hb%'h"Ut��k��@�XV$�j��?�ؿ�����;���|"\־e�c��Qq�1���m����PAC��	w�N�&�����1�  spf�Cu(���&��0��J����}5��ݞ��0��*n�d��di�(���l���1�r30P�d#��g� ��a�,s1���c���h ;�_Dz�d��Y��b���#�Vn,�<�t��*����o��C���������b����VL'���/� �4�[��ֹ�wk���w�_�ЄQ8\U y+�3L'��18�k��Y��ƍe��a07�b�0^���˸�0,F6)$&�`3D�$L������{y_�!RH�&N���7
�#�O�|.:z�T��DcS�8z�|3�J�0�i&ma��z[�q��wpL_m���<}�?x|Y?�bpV���b�?|��A���KH(�w��0ZՋ@�G+ ��%��t|^}_χ��A�4j����m�}iQV uhTyp�B(N���%�����2d��jrޥ3����P��?$��͢�W�,E}�Dp�2�94������N�l����27R�̢k��ۣxC6,ݜ�X���j=����� $�z-�H��:*����y=.x�G��j��h�����c��o�(d��b��/���~%����Pϊ��q�D�%C|�u$$��cdS-��V��d1C�9E�������VV߭8Bԁl�Q=�2�<}����I��^O�������9��bH�.炸`d��3X����Fej p�vݤ�Ćr�~|Z����4��$���m�^������[���.bp��\�"��X�~B���d7����gL��E�A�����!ޔI_].J^�{��LU��"�eU~���G��� ��F %�	gI7�Q���V�%���q�:\�1b�;?�<,��?:�X���������q��sT�^a�֢=!|��91`eJ"�tz]�pV0��O�,��sEl�m�OȞ5��М��H��zd���zv8`<o��#��\(�6�7�l�7i��1�*�dQ\lO]V����6�죓�E��@��lW��B��('���j^���.ݯf�-�S�Q\iw�t�z�s��M�tԉ�����vd�A�T��s����j�f�i1NЋRQ��QT�!���Lu B�{�����u����㐖_d7�2�lT��l�@f�+�͔�����YuV># ��J�i瞇ߪO�qtI|���z��{��,�'��1���ʉܪ�ϧ3\�����^m?4�)Q���lIeF��9?��|9��b�C��x<�K%��ڔ��]w6H���$otbhG������C3�(�B+�0o�)�p!�/i ���v�ӗ�A����; �!S/M����N�
�g1�V��ެ}�`�Y�K9k���.�<�Ŵ�iQ_m5=�m ��\02,F�UL39_:��4��h�x���K���&�Z%+��CC�h�}���c��#b;�b������#�_�!�Zg�0���3�n�����4>�V�r��hOqX��9�����HWO.�M.�%�/�NZm�( � ���<]����>YKq4�+grE�궳@GD(g����3���h�d#��z�x��+G_�����R���uv�,`�-'ؚ��=��u#J�@ǖ8����P���	h�Pu�?��(���W���d� ��ɘ��I��u�k�ӓ �fy��M���Q1cUt�O�@��}�e�]ϼ�_�,�+����"	G[88���&0�G�l=���C.b���m;CeR��i�ӥɿD�=�Ϝ6����)X�ľRf)O=�=��?����zv�����ݖ8q��y��&i��V�Z`����yG9`�{ӏ���G��ӂ��N�nn}�2Py;��������B2%�g�
�V֞�=�����H�:@@��a(��礨`E�PL�u��ī�6� �T)V��s�.���0n������π�����k2�M��ֽ����:���w��������ڦYg����
c���%�G�8d�n]xg�����j��m䅖M1X��7�����"�d��wx]�?l���N�O>�����r���]�7�L���)1�ƺ;�+���dH�J}ƥK���9hQ�hϠ�Kyi�	�oU01���Plh7��S�".��p���Vav|��\�v��4)?�<2����`�\|6W�e�de�
��4x+�����Ը�}d���k�c��v\/��z2���N��%�KN�FPC���yn
��sW!�]_ܬ=F�|G�+�컇�X�J�"�C�6�5J>��x�af1_y�i�s9�_-������H�it�׾tۨ�^��r�8��"�7eg�Re:'<���Υ�mט��X�H6���WSSe�z@�aS����2uZe������M�e4�4^*��-=�Y��ڥ�خ��v
�wc,�OX�����&�҆��yރ�]w�z>���F2;A�o$�V��A����p��O���(��T��U�	K�Uģ*�4��=*ɚe�V��'�9y9ZW'H&b�R,�˥j?̮#�}�r$^LA�.y��1,�+0�e}1$(�mxdf������%m���Ջ\#�6��T�fwJe!�`�?]��Ɂ��p� �
�<�
a���y#o��L�	�T7a+�Y|�:\ќ�ػ�f�O f���b8)�*@kC�2�����;%���e��у�H���͕K�Zh
������p3�U��''@�ɼ/F~%�Z��V<CjRC���!�E:����IK!ڈ?.��5դ(N�8���e6���<F؞�B��r�r�Ze�����!0� ����D %d�c�,ݸ������8^��R�]��9�ɞ��1zf����FoM���g��eԚ@�u6�%~e��u��k�S��j.q��fz�����I���Q>~�����g<�s��9������Ǆ�Ew��@>�q�.�=3��5�Btm��
�}�i������]�~* ��0�8q��qr����H1Y��F�>RWđ�v�͆���*�b}0���t�,LDD0@z)G�m�=!�U�@�Ǯ��q��s�j�{��Hqc�[�u����$-���v����e�x�k��e���n��=���|�]�|S�L�y6�V�ԅ�)���ֱ&�-�#.VjM���h*��C F�{n՚�ĝ��8R,G�:���r�T�K~KL`�j��]���b ^Ž�s(Q�пľi�*��;j��m�-���8ב���]��K������x%�-������˒-t���+'a�'mh������!���y�7̈��uacZ7@����p�j2��i� p�@�t�/s
��F3�m.�'���|u�����0�z${��7�/����T�����&Xx��������n
ě%�jf}e��wݻ��C�J}t�]-7�"<����͉[�	;+<N�Dy�Kwc�нBjþ�J<�܂gc�e?��P\�����L�����3�u�����K|��\E�`'8Cx�XQ��c���LH��h�����7eL.�݆���	��&$?Ʊ�����_�e�a�3�$ɯ��=�@�����`�t��I'|�}~��{y�#j��_?�L�_��I"D�����@�h�m3�P�`�����}�e|��y
��Cw����Bu�����1;j*�^}R�
ඞW�%6�~73�Ya�W���z��'��4�M�.6����9�~��z�$�yC��%ݘ^���K�^ۓ]c���^sz^	�$�ٮ�I�ԅvKz���ײ1��a~�5�*{NV�
4��a�$4͂����sI	�v���4��
�]�;�r&�&��2o�Q���@���Md�Z�ݨ��jނGu��9�~x��7<�$���W�!X�$ڇ�E���(Z�u!:E���`cT��⾏��aK�*Y☳N;���!��2^�*�^U%IșV�\������4q���ɪJ��k�-�Z�s@�ɘ:��g�\�Nz,H���$i�O�?��%"�=Q�'�hڜ�5��)P�iT��M�~p���c��l�'h�l��䓰~"���)�ݤ�cH>���Rg�Ju0j��6�Z�O���kQO/��N���u����c�#��Ȭ�ֶ ��@�j��?AW��I[�ORyR��ek��]~�3��v*Ξ�/.�+���=��H�(:{�Z���BIw�kf�Έ�I��|}@�Im����]�9z�1V��b�c.����[7ԇ;�Xp�u �0]�e��5cj��>`,�;�:�i��ؐ�k^��۸WaD@tݐ��V3�k���;҉��Џ8� ,����3=���׽:?
U��r�I��.9��y#C���#ETɵR�������d����~��h�o��n�f�����������့Z҉�i'+ {,N.�����+V���t�����2(�=\��|�-�n�4�e����t@����^}��$�t���?�<]��I�������8鎙�;������%�uz
>���H�R<��bv��]6�Y8��*�h�E%���oq]��i���a�Jq���6|*uP����9/�=�hj�OyD��o��k�u�}G%N�p���u��\���~�z�v_F[��\j��X+`Ž���)@z��56�6I��-�M������^�!z������+R2MBc�Đo�lj�LQ�'^�%�V\�W�h�do㏎�4��|��8���!�\��/��Nm��7���kwe�^��p���#�Wv��s{P�}��a��RL�g4W2���7y �ö�0����+���z�bQ	��D4j����td&���)�r��!�c��^��S��y8-j���"������~�D������v��A:��e/M�֬��@p޾y		g�P�j��|u�� V��
6�6*>N l���>��aX�s�ه��t߽�����I�5�(�7��١��:��Ԍ�_���
�j�����i��L��^3+�r�|��_ȴ#���F{�j~��☓�N09��r�;?����٠;3��'t�G+�R�D���dx7^ �m�Y�����'_j����~�����w��~��������>�8��lP�=uli)���t�I�����-X�k�+�'͢�=��tB���&߽iܑ�>�S`9L�
J٥#��?��)Au���Q�8�����*�v|B�������=�16����ak@<;��
���t�N�9�iv��@@Բ=��.���nй�7�~8;�ކ�����7g���DY��>ב�F�-G�C�v�d..��T�RqK�^Z��ɟ�=����񠈼6u&[�-(�3[)��]�Ln�i��9@J‚�"ʀ߀��JvF��=�$���'{�:� �ZX�=�|4$�D�}X�$�m�(s#����
�v�E%��p����d+�����hꏱ�3�`����6�%*�o��[�0i���!�Eq��s$y��0��Z&�j������N 1�|��Z�NN�Tp]d��g�$%f�ե��{٪N��9��s��*]9΃1�G�tF��M�g�w���w?�GZY����/��|�8�3-�|zj�E� �+�0V���1��zuT')�)�';��	tz;�H�j�O�7�n���������oP�ל|��o�UY���D�YJo 'G�O���<��0�p�C�lz��S�D&x7_E�d�Ǵ�AI"�S�cz8_*'b�����ww�qa���oґQޑ�P����D��&Sʏ�(ʥ_�`�=�r��xց�n2�u3G��.u��D�� Y�*NTeY�Nچy|�	�Z�E���Rs�-��e>ZC�ʌ�	������ ����	��oy~$�=�-�Rݒ�o��Y���r�cZ��!0�a<��%�n��ڋeGZ�	BǬ�ُc�b=�0G�y��Q��*���Wh���x&�3&���'Z��`3R�������U&�è�c҃h5`2-�r��נ��"�$!�?o���n��Mk��h��^O��P�Dvi_6o��d �6���U�)�b&|����V>I�B� t���9��DF��Fd�- �wj���e�s� ��PJH+ԝ^�*��-�6ؘ���:�8���z,�^����Kƹt�j�rc?�#�x��1A�����8��g�+��`�����(Ϻ�ya�N���2���&�N�J�V5>>�J~�M�dǕ81�;��=\��t�nӶ39��6s�v]y���U���$���a���5�%����)�����^(�]�}nkl�U���	���G�Q�i�,�#�ο���c��]�^+�s�siLJ��Q0r�ț���̧�=r�l '�c�lB\���~2.w��`Lu�yq]��)3�7� ��݇@���]Tp�2<�8��9BT�]ȱ�8�V�2?2�X@N���\�5�y���cmJ%�s>�厜ߡ��ܻ��,�KGqv��r,�d�K����f�R1����p�+zP(S�z�j�ܺ�B�WH�Wb�{H�R�����ۆ~��&�4���)�Y.�1>����ʓ7W�1z1��5i�	״S|�~��|~���@E�
��G#��_,�ٰSE��ֿ;�UJ���g�H&�~��?KG�4hIQX4.�dɽ=����H)������W���QpcD1SP�;��i��kn���u;���Ygz�����3�ܡ��wS�;j�Of��ó�6���U�PV��9/�� �T �oQ���� Za;�K?6��"�Q]�ч�G��Q֥��M��t(h���#.}��w��5#�Qv��iC�rg�BKUS���Qtӽ�t8/^hWB��큔��/}c6#_�z���Xx�,��۪띣e�J�8��M%���&t��<�m��k���w��l_���&���r��Q��|�P����?)"3.Q��X��Xh;������i:7HOJ�0�CD+қ0u�e���㵌s��<���?���GO!嘘���)� i�����H=&쒄�"H�uo�*U�!��G���ܵ��~�4) "\����Z�hM̔آW���P��t��Y�a��d)�܈i���� ���$�Ib	��'�X�K��/�ʥ��gS<��)GMv[zr���7�J(�X�A��φą=����)���u@9}#,�~txa���mZZ�&�:>��>ק�5 ����ؙ͆
�=*�ǖ�'�����`o��r�)<���*e�}��?�qc���0�������Z��0���n���*�/�E��S%۷��St���Uxn�����b~4t�?�7�`�e�W����ᯯؓn�a��N�b���y/=� 2�*,��JSx7Q:���q� ���x>���j�"�&l`ѹ	�ݤ��
�9����Nw���Ջ? l��c6�O��I��/6ɥ�/WmO��яFK
�g�<�Z/�Υ��2EM��Ήz*Y�d�+�'�>)��\�X��^	�I���ཧy�
���*1���-�	�9 F�"����0��p�$pٲ7���}YH��ԃ��\��A����̸S?����*��uݖ�k���B\���%��������t�EZ(#�*��r��C|~ZRjvM�|)�� �QsAt�J��2��nz ���Wq�Ⱦ��Z���B�w�`����z!�~�SI��|?8nB��3��� X*?�%�Q�-����y�/#ꋀ����X��|||�r���1��2�٣��I�:�p ��0OS|�$���@���p#p����d�Ǯi�߅������|^�������@8��b[Hm�K>D�f�[ߌU�L�gW��$ˋ�����c1�)};�\�+�9}�ğ�~u�+n𙇚7鎣��a	�W�~jy:�Ϳ�6%�HWg�R��w���p��&��	L��~�e��7���pc�
���pV(�k��V��@�=޿���Ӥ�	��O�{��T̮���Y׉��t����B�Ҋ"M��DEa�9��d=8�P1-j����P�w~�wH˯�^�C-����e-��B�_�2i���?�'�
~�'����1�Z�@dC�S���=�4	�i��]Uj�39�Ѧ��[���'��bئ�ʞM��������|�
��)X�9XQsGy{_�K�h�D`(p��������|�Hj��J�-,�d��p��P<�*�������l�����1Ȑ��2G`�Xz�b��B��{0���[��i�Ani��^:� �E=#�n�5U~Fz�S&|�P�u$���
#/x����-�qi�`��f���7���Y�2'�c_],V^��[pZ��1�b����W��t8VCG��X؆��ó��x&���`k@n���/Tw�3АB��U6=�yt>��#8��)�@���)@�D�]�+f�a@b� �똬���S�4��`D �+(�6V�z.���Ae��z�9y�?����_�E���옗�2逌��\���^�(�)>�lI��&@��\eS��wx}A,����{����akhl����������KTe�03�ɔ(�|�+c��Dh�m }T�}�����nE����P���(
_k!cD�#f�0%�������qq���\��jN�O]6OS `����_+>JW�MfH@����.ċ�,hs�`1�gz7�$E�썲w�Y�׻�u
��,��L�Дx�q,����Q?^>�N��l�j	$�ɹ��~<%eq>���{YV����񸓐�;�28Tt�-�#J@gU��"�`�_s�Wo���t�w��
ʍOC�;<hj�\� �H�0A�;��;n��AkR�A�Vg���|CM��0U�,*g\�9)>t����Fi|��(?�<�-�c��C��6�:*r�l
�	`v^�̐��DP/�ܵDb	��9X� `��T��GI$~R���C鰑�$Q��j���_�ҟ�JryZ��y��4e���n��`V[��G�aB�QR��`�xe�  ����	���zU2WL��:����}���2����Pv�����`kق�x��K7����"d˛�_����Vl�ck{S�"�|�a���0]�(�H�D�����t���Rw �t[�"�$�Zz��U�[T�z9�.@p�E�)zV^�멿�y��蹽H�qӤDF���k�9./Q��S"=�iD�p�$A�)�3sy�i���o���Z����`�Ά��#%af/~�s�WZ����C �&eQ}�A�D�@�د^Eۘ\5a7��p��nL"�+��A�ăU#��.��pU�(N���	�Ǿ �1�%Ӓ��M(�@W�W�q�����%�^l�z�B'��)�63����/E�A=���h\J���԰���8�t%�:}��e-��TKa4���  ��� ������D;+0��\�c���6#X�U����^�p������a'��k�3��K�U#v���&����qkI�V���|�ۆ˄��q�p�ʓu+V�T
ŧ�M&�(�r@7��t�����j�Զ�Xi�6`�uӴg��g�c��N̮�/��%��%�|2�$~C^��17�E���z�k�ύ���oTmE;e�t�;5�f4����4?ڂ�G����.[o�U\2F$�bb��pD�+�ϒ2�n5lêĹ�Kgк�4p�8'�u��G�wȊ޿w��<+� T`*lʓ_k�7��5Y��mY��4v��0RP���UVgy�c��/IE���l��L;)�j����ȫ@@��,��j-��ᰇ�6{�z��0���:,#� �M$�NNz�S��G�7�=�4�����yz`���]4z��jNۢ��v(�F�=
����'P?f�rIU]n(Uqx+";*dP"kg�0ؐ�LF;�g�%��ך����������K*�Pf|R��/R��EH7|��53��|7�2��Ȝ�8��&�aWu
�Ǎ�$����4��3P�yԵ>����yT��=���p����YPEς�+<�>�D��+��RF��ⶰ(���Z�&���8���0�2ğ/�)
j����Z�Y�Z#W�	�zgA�_�@>{�7�Zi7aT��
(���F�Ź��=�}��(��Ǻ��2�H�&2�r�5F�޷%�F���W�D���,���.T��"=�!P�q�Ä���K2s�Z������0�ž�L���Vdl"�'�스��a��.�*K�9漏�1��,�O@c31�Mom���; =�ERbsP�f�9:e��n1(;x�S���`� �B�'�V=��z3�X�a�Ҭ�ůt���� ��f\�������ϱ�؀��dB��5$:�v��wub ,��vB�
�A�E�-"�3R�*<�l�F��8��=�:J�����+���%�bO�'�Xø�ӍѬO�
�x_q����{�`��6��2�'m�X\?Ŷ��ރUo�U&̮ ���H����E�L���q�DE�ɡ�'[���3�MwZ�I�#7+1��O_�ґއ�^4���~���B���/݇�zIJA��@Ϣf4��p	���X݊����t���ְT*H��1�����,��8�!�M�	J���O�Ѐ����ү6��/AC���������<T��촋Jрv��C�=�O�
i�j�J�Q����KnQ��8��q�����قP���َ�8(�7w1`A(����k�Q�#HW��x���\���~�p���5B#���_�P�֭��K��V��e$?�b)N�V�B���P hϼ�g���W��*��u��6���X��pUى��_G�Oj'�؅^Z��6�Ju��vi(H���JiY��	8�Z� Ȁ���ԯ*|x	hmdG@�2�5����|���n��1TzC��<�����v�	�wy�֙�*�pZ���a}�(˓D&)D���O|U�إpyk�ys�f�>ЭS:��uzC����x��aװ���0��{��?0M��7�:�.53��L)&��ۑ�����xڴ%�Ռ'Gy~3*)E�P�i!��~+���&���~�өy�l~N��
��.� �Xgť��㖒�ؚ@��[��W��R'{���T�(>7p4E&�g���ވ� ��Zi;�m[�%�f������ęT�H)��V�z��s� 4X�7��ar�����]};e���%E0#����|�b�w
�G-'�99+�5*r'��0�<#~#,�W��';>�d3PJ��WځD�,4�� 3l~5 =���-n��n��պg�k|�]�⻨��_)��̪xLx�mg{�4ʫq��r�n��O�N
�{� ��'�ʗ
vF���������;C"q���熓���K�����?Ih[� ���b�Q{%7�p.R�#�K��Mr��Ä~�W^�f�n�zZ��D���/����.��'�v�c�O��d^~!��~(������x�斫���i��Gv0_bQ%�H\�P%�5��v����Zo|�A9z�b:-]tОX>���+��۩j�z|Q8�I<���k�py����>҈rx�h���_f�5�F�4^�Da�'����Vj�lWMz��R�8�$C�� #�P(k��e}}�jf���BxL*��#���E���k�ͺ:<��^�0<�4���ii^��!�|�d�t�[�X�fD}�m4^kW��V]�#c�p_h��p�?�92+�;�`�n:7܋fMvP.OH0�-�� nҬ�j.��O��U{�{B8Ї��ثqd����g�4�AO_�&���&��c1qnwN>`��* �U���5,Ң0 �]�!��:�x0!\��gŤ����h�Q5wFB"W�5��/��Lы
p�D>w��C���s/����5ƽ���B&���Q��c|�k{VQ%~�z�[� �� [�8س'���a������W�k��^�Ľ�9��45aIg���C��h��Z�Z�p�j37��O!�p�"^���}Я�ė���"lu	5c�ޣ��g, ��(�6��/X�_}.1�ɠ�����ۅyϕeϛ���i���$H�囒���/kѢ�ĝO�@�o�-g��|'�N�z�n&1�ۚ�m�r�CT��Q�[e+"�dl����Yp�#jhy��r����m%�G���L�����Y��\*r�� �������nX��.�P�6�7��*[,��b�ݱ�萆�|TZ��K	�QR�BΓ���ԗ������L͠�[�ݥ!a��u6PIDmS����"��.��7��(+�#��  5R1-���(:` 2ڃAXl��|��Kf�-��\ '�,0I��|ܭ�:sv���*�y��� ��;7�P���he=�^��H�R��}Q�5�кS�3!�� �y�+C��V d�u��b��<i[�5c�o��)JsҔ'���4vއ��3?qeY��Ȋ�Ȱh��RW�?�[�"tC�`����C�;�>r��D�98M�[�v��q�*����@���]���&���8�_e��tN	���{f^
�h&��R�XЫFQp^LÆ=�*���E+�\����c�g�C�ϓ]���@��%x`�vwx o�KS/�-[��$�6�u�z}���gC�mH&��?���x���@mGN�q���X�QEf��jނL������F���hM�>�����=�Jxc�V��}�i���dӬ�:���.�g����dUR������G�af}-�3a��{\z���5EQ�C��w�!0�)ѨVgz0��[l�A^���,��-�� ����{mُ,!a����"$!L[.�][�Z5�Č)�
�w��N�M'b��oզ-��{���br8!�j�$�G;a.�R��/m�:�g@a�ZG�����d�A_�`3C(�")��X�)����[�d�>��.I�5s�M������ήj�\��(�.�Ti� ���M��C��Q�l��Y���]��H�Ŀzq{2|�o�[K*��{��0�D�'��z� (!��#��_�1��݄�$�F�I�O�|pN�e�W�ޱv��û����1�U�!��B�Y�`���Ӥ�B��a��+h\w-�o�	����&�9��>2����f<[��ڪ�bB9������M��h8��se�@A��Ћ������
�g���{�r�����6��/��q��sJ��$���R�W�m�yw�5�h�4�I��H^S�0ئ��ɋ�{�{��]AA8V����E��D�bѿ�i�IEq�
����L׌1͇�.�ZE%�'Ьm[�?�Zل�!�+��}�p��r��o���;yK��k���-zl���V�wl�*^{�0J���	�[Bdƫ(y��6�"�}�y*a�FB�����Ŧ�|l�1.���ў�^�l~XZ��w9D2ڤ���5[H�`��k"/�2@�a��a�;�X�˭�@Ixvu~�±�,��5�뾸X}rP~
�I��da�#:����J2ݷp��2�Ted�ڨg�`v�wI��5�A��S�'Љx@�5w��p��aQ���u��qj�&��^�gW���t���b|i �ԕ	Pje�M�M)d�i8��b�p�=�߃5|0ʉ=ȩ}0~YV�e�+`�\jW�)ܫ� �����<1L	�����<�XuT��0;3��'�v�2����X�[�ϱ���ԥ���jH��L!�F�A�A������E�)_�-�Z�4���{�ˣ ᦿ�D��na~H}�;�=�\3FzS4���I��_��N3.6e�o2L	�%%K�q�?EC-==N��}��n���bzf���-ح2��M�q�.;��Ȗ���&?z��_\mu�Ǚ���ŀ$�x��� ��>;��bE�.��{�}�{�{l�պ�T}��G�iV8a+cP��h�`]�U�Dͤ_9Z�j{�d����^Kb��n� �>4��%\3��;��%�d�ݼ�{q���#}GB"j�D$p�{��a5�5���.)��B�=:���W:��"��%�r��  []d���,_�3�'e~c_I�f����'F�G�y/=�L������{\e�U:a�$��1,������0I0�c$Ǆ�$��G��ᱎ:����¦��?d�l�����{*�r-�����eZ�Z���rъV��w�`�K6>I����{�p�f'�rZzy|�S��
�~�,�`V�ثP#]R��zd�;~��Մ���R4{�93�oDPM�8��r&���ofk�w���Fw�R���Z���İ6e�.�*�^Џ��H�� �-+Z���	��o�c���X������u��6�`қ�ֽ�I^+0�� [��6�q�k3�s��J�A�+57l�Qv`٩2�{8DkEn��ں�3A����΂�l�:�#g�B�Qc&990����v��b0�uN�7tу�I��/]�A-�@���4Q�O�Wmo���U{��mI������vN�_�2H��J=�6�v�.?i�|Ǽ*����������Č�t�+�$�(�q�O Լ�v�Qց$����:��r�v�`��		&�S�3O��}������m��w��7������h�/���/��x�xx�y�ʧ�c�yaV����ȀK�x�l�����M,���C���N���34�Xݼ��+��d��J��##8�h�֤���˧}��`�v������ͬ(�~��O�>[���1S�xW��&6����*(�I�=�sl����xh�ǻ��mR��We�`�Ϭ@\�ߩ��)2az+"Ĳ��$;������S�x���?��	l;���xb�sM8��EL_��zaT-��qF�o�h������b���	�[X�>9����@�:
���������Ӻ��b �'�>-��/�bܲ>J���s���@1*����I�����T�2�Aj�Q�}OP5`�6��ZI��������PL�����a�!_�cQ�P1~ko�6@
��tL{��,
�5�g����П����O�FB�0lnKsaG�~	^��y��!.Ev���F��WVC�̲NG%�5�7���iWl,0aQi�çޜU]�i�YH9��u���ٯ-�����M���gJc�Q� Ч>1�Jg���no�9{��R�6��{-�+����D��I�3e2F�m�!��j>��Va�g-�2����$ �� ����5z8F�5�B��S�;wzΙ��TTi�N��@3�d�)��/�j�U���޾h�%:��ߝ?�<
Z�@�u1��^Ihᎉ���:%�.G�r?��~~kj�7Ck��� Ŕ��ϵ=��m��^�ll���N0k�Cxb��Φ�&�����l������.�O��O�R�	�(����x�����Qw��u�f2	ɛ�/n��3C���w��]l�C[�lW�2���_���R�VP[/��xq~$}��]��U�d@��}��:��l��ED��[w�OC{l4��|?�c�5X��q�ƾ����ǀ������P�U�6!�  W��̴�-`��O]��[��=HWd/��L�/���[rj^��a�,��ހxo�$�����e�Z��ɡ#4��Kt���<x4�5�29l`��r��.�b._�<PC;5	0A��	jTru��l�}Y�{�ts��O��yS����GL,��V�
�gq�3�J���^��H��� 'È�4O���2�䃔�^�V3�H�����^)�ߧ�q���u�X18�ͦn��a��S�=��W��'��+Β�R�Ӟ�Nn��Fħ�����M���E7����Jp�g��QZ�
�{)H��}��-�PP��z�]�L$�Y���>�l,��)iT�X��R���2R4��7lJ_#k���Qx?�����U�l&�Mq��Z&>�=py�Õ��J��bɋ��*^����ɽ���`�{���g���:)���):Ȍ����:q�:	l�/�����D+��M��uqg��ۚU��83�`���`y<DhGt���)+�<���>�$��`!�T,}N�^b��}�E����tS����ӊiٱfoT�{���L�glk�� �� ���tx4Z}�35��P�Z�ӳ� ^�T��$���>q�c����g�=�M�~��㐤	G�.S��4�n����%�I"M�i�ւ���Â$C���b8ZS}%��z���p	�� �Ӵ)2��9���������5+��H�ٰ�T��`���N���y�^')���:���6����~-D��~�-�r��S�Ƃ,Eb*o[�CFIL��=Ӕ��`{�}S8�R�̟<��a�= ,���s�=5R<����T]����4�M7�vS99s��q�#�B�t���[���](�Bڪ���[L�7�>�2P�Ď'���PҺ��wE�'XT1܇��;D��e�f�-)�;�.t�<(r-b5ܖI��G���S��DM��*�q0�|��N�{�R6�EA����7G�H\� ��۱��h�CN��ijм�E���/�g�l����R����4�:s݉�6$D�g*خ �TR��F3��� O��^��֦���R�+&��	�t�:�5��f�M��R'�Ϸ�x5�o��}͍�|`�a��3U[�>���>Ṡ塓'm���$����4Ķxu�|�Ēc�Z���F�ck7z���#���S�Y�3ErpH=Di���8�EV�3i�p�Vc��vt��h���U����������:#�5�7E[�h��p�)Q�i(�V=�F���p�~��K�5�c�f�^��$��0I@|�<��]s,I7�@��d$��Vf�_K,s??�2HO��?�w[Ī8.�M���ZMvίC$���f�$?g��O��w��m�lV~Z���-��t�2z����YJ�"������ƃTyE�Ġ`w��x������}��im�'�:�4�aWՍ���r<L3���s�Tf/ L��y�{+��J[!��R��I�$tƇۏj�}�TzzvAwN�:ڎO=\���t�}�P��7�x�9��K��n8t����A�������"�)]q�P���q#�{��&5�E8�AT��$��AbZK�&�b��x�?�UM���h����W$T��B�����Y���K�*}	Wr�"]N,�ɫ5d���m���;/�Ɏ������X5W�� I#.�l7�O8�� "�N���fߺ�
*�e�Ԡt�9z=}�Z8��3EN>5-X6�cyr�Tp�:Z{E�w���v���/�Gc�2�/�����g$�����=�0ߚ������=��ኴ��Ā:�AmPB	�/($뎺O�я�{s�tU��u8_.Z�}Ҽ:
�H����ئ����3�k���O����)��b�f|��Q]'��̝?�IA����eV/���i�[�?�?�IDQO�i5��p���J�G�����c��ЀR��İ�e7p��	���i�ejMLۙ��n��Ό�}E���C�����/e\��.�4�C�>
ޙjgA`�[nX:�F�B�"y���/vt`�U>G�&�z�vNЃ��t��u)���~�^Zd�����M�6�S�}��~�� ~��P<�ʗ�t�U��K�פ�]ܴz�a<c��¤�/���F�������_�Dq�Ty�p[Vl�~�kk>�#"�v����<�H��T����F>�Wp�9�����_3���5��!ѱ!�qBƈ蟶o����(Y��_h;������Ci��6���~��b#��qN�ظ|���a,ЀU�SnAv+��9�|���!��L�&�2è��[�jd0}d�]�M��Y0h{����6��.:��1P�+����<�%��3LPqO����0V#P-~���S��r�+ᣮ��i�~��n\�,���w�)��.��DG�}[�k�a�n�3�Vv멺�=�� �07Ӓ�qّ_9�����;�Jk%8�8��&���f1jʜ�g���O�~mW�`VۂX��J!v W�@���؃Ň�`j(������	@�׫-��t�u���Z-n�?ڦ�N�'���Y����	i�k8$/k�j�*R���8b�� �8��f������~��cD��>@�N-�xfEz�	��k��АXM����7|9ʆ��d܆��v��0ac�NZ+��W��d�6�|�Rʋ f[N��Nن��P L&�I�Ԓ�n\eN���m#����`��-��>p>)`��U��h�'���� �/4E��1x�v;����M�E�m���%ڧ��}���&[H{q�_L��ސj��Q�n�F�5\R�qvfD�:)-���l��%��Z�6��|�Lt8~|2�D���$'Ok5�hF@��J���!y#�gR['���{�Q�]>��zr�
$��8��C!,e05���<�tM�|y>��Y��g/ �P7�OTd����#��p�2��NǦ��1�*�ۈ�?�{�V�V	��^����uw��t��;L�_>R�?�z�.g��Ǻ��+g�ׁ��Gk_5�;5��eU�\8�#�."��]+sVC�@�`��+���8~����hH��Gky����X�����Ȥ�W\��������/:+VX�!����a���W@O��=ĊJ #Y� ���(+�5��r�\/���l'Û�䅉�T�.^�3�}��|heȤ�)^э��$��<��h��W-u��ƴ�)i�k��3z��j��S��Z�(wʘ��6��!���Ҵ�,��O{i����&]H���N�~�.�fO�t�I`@�f?K}�����" ��5o�^�f[�Cv�*UhD�cq��9�~�?:�O�Qâ*"��~��t�si�t&oB���U�<N9�H�DVք&��r��]c�Y�9���,F��]f�ѷ�9�4�a�)����J<�<(��I��$6�-�S�����2pNYH�x��p}R;E��V�
��
�*S�7�Ө�}wS��l�R�d>���*^6��|ѝ�#-0�`DH���GWS$��{��PQ]����n$����i�^A�8�s%�V�L��Y!+<�uiI~�dO�Q���C"C˴�0����]���h�Y��L��7���N�ė���-���5�1J�xg��7���s�h����"���%g��5��_+t.x����*�\Q��ڲim��pE�'Ƕ�Y4��C�.��T���|��!����'F�]�+��u�����R���0S���r;�t�P~U�L�;ë��N���J��a�E�Y��UCI~/��|S^6b�K%����I^����+����L��V�h���zI౟vQ}JV�f����������X5��g�ƈV3�q4YP�t����x��5�Z�U�hw����*�}"L���X|J^�D��^�O��Ad�-W$syU܇z?�mb��$�즚�q���;ZX#���(�h�#�����E�[7�g���Ū����[<&�V'��
���p��M�t��0Lk9�2�7T�c�!�1����7�<:��>�e
|���%�)�s���tS@�J�9�hh��u����M]1�Q�Э(�K���=��b��އ0����0s0��d� ���ta(���~]fa�S�M޵L17gu��q���d�-7�}GQE^(X8^�k.Q��g�3�k�v, t��2"�ȭi�⟚�/�t!3Y�ʩ4@�b�ߍ���Q/�_q5_e��{F%������-�LmY>E�y���J�P�Ç@�d������|��H6��^��=@��c~"/oq@���7L����e�}�iג=�Z����-��&g9	�|�1�P����5���l�'�Cp��l������e�ڛ�[�"�S��u8_D�ۻ8�6d>���!("tl��o�5���Kхz��aG]��ȾΪd�;��Ƚ}r��$��V}ge�)��A��}���7=��ș�U�'�6iϝ��'��}G��ԃ�Ϙ��mQ�錵	9�����JZL�&o_rˆ�t��*����!�@߰���DFlP����;��)D�#`�(�J`��A���+>-x[#��u"�㐷s_��^�n;� ���>����o�-ۜd�2�~����(�Ȭ�K�> �Jٽ �5k�gd��ĕ��}�1���������~d�y��$p�?]�U���/�w��x� E��~�DZB��׳�Y�;�5����|]�&��l���P����>�eo�P�T����)�k� ��ÿ��aᛀ"���z��D����ޟrl�<Q<=G0�H�>,��s�D�K�*�o:�inQ=�B`45��e�<��gI��b�c��BU��>��+�HV�g��@:g�OzI��|Z�K��r~^��-����@�RW:�r�Y�ؕy�,E�@oi��Z�|p܉$�!M�7٥PI���&������`%�`>�{�rj�����l�hW�jl���%Ksլx��V_o�1��LW�zJY0w��ɠ��8���+P�V���EΙ�vE`��̦�����oF*�e�Ǌ��6ـ&�Yޝلt���Ю��.ۃ�r��Q�p<F<�p
�q�_q�%��
����Gbtz^b|c������澇�d'@������6���7P�V��D"�=�F�V�@B+SV�)����'[5����j�t��Ww#=�~�9ڝ�[� ���ˊy%gEΈǿ��=!�  �h��2�vHZ-�L;>xY�G/'ĨI��r:Ni�)p�N)[W�ǫ��,�H��"yș�Z
�c���Xo�3�nw��D\�ؾq��	h(��8�d�xv��'�9:��֙��?:@�TK<62>�E�u7I��5\�� E��`�o��7����;@<4S�T�(y{��.�p��<��7��,nbp �g���h��ڽ�tx��?r	! ;��8�6qn�u4��^���Dw�Q��_�-Gp	��4�K�!uL� .c7	�?��k�Uم1S8�{���rB�]��%b��Z�0]�}@NB0�&);�]��D:b0�?�P@��.@���n�$�l�dph|j&_��1���ڒ�, yo��w�^��]�ҀBl��L�:3�TL��]��[o�T6�"�C
r���A`2%dIh���>0-r��1�¾I�&A*Х�%�;���B�~��*6"V��� �7˩l��u%v'�N�A~H=g/u�|^J��YJҧ�0j������z<rfy�qPU����.ӸwLvB�C
�cv)�C�-�C����n�s<3��1`Y�.#�h�oR��F^�/"�a�������nRf`0(��2t�i"Q8��Z\�.?��$Jc0o�[���P�+�l�S}���0�LUyO�.�ێȓd�H����A9)e��We+�(�`�>�n�w\6���i
��".�g��C��jR�4��~>,Ɠ�� ���������Ŏ��ŵt_7>�+D��E�Dx[�w���򜯌��I�k͹'�~b��j��ji�1���M�Ւ#�]����<�2�E�?��+ ��d�K&q�D�zT�"r�G��@A�v[�V��b�/.�O�i;G�qk�ʯe��/�چR3N�2��ʟyI����?��r�u��ME�g-ReHG�-��/��pq�q�FH�a&)��R��6k?YE�E��*U͋Ë �Z�FD�Eք�R�Wq��u���r.)Q��;�[ �#�EL�[P�t�[���O����<�]�ǂ{S�mX�Q����<)_k(-q.�+�����.�N%�n��9z�	�� ���'��C�E����1�ts}��p�9�[ZakP�,� Y�#�V��HĠ�����Jwgx�^&2e=[{t	�fS�l�v�x!i�.z��I���P��Srm���/��:ܗW(���+ ���ȓ^�?~��,�
�E�`]l��0x�V��f�w�-���C�9B�X)!�6
Ǹ�"�NOZi���'�O��+#�./�' �R�w����+\��|���@V�G�l�<��C��);�c�E��%��5� �"4�w7�ʛ�`���ic⻈�I��q[�W��[���0y<�yTB��N��*��	T�x0K֮�Q�<��o��Ŋ-Wv8=�[\�%vJĸ�kR�ZkD"F�OKT���=�NH�2���j0�cT2�G.�/NC�<�iD�GH�d^ȯ�VG}x��;��?�@u9ZF�"��vmӛu����'��y午�D�}�d'>BF]R��D(�gӦ�G�B>�y�&�z��*wґ\�����J���Sy�t�k�]w��RY-�ƴI �	�4������i�J�%��&qi�-��I� 	������e#X"z�Z+�����S����1�='+o��+���*Yȗ��u��6����z�k������{���tQ({b���n�����.�]�H��]�4�'��-9&?ũ��w�˳?/� ğ�>�]������ШUa
P��NwMX�{uU������:� O�6n���6������I�P?�:v�pv5���g�����bL��oL��!3�O��/�{�~;�Oͭ�r�J�%Y��Fq"�i�,��w
`ԑL:␛�	�'U��j���Q��*ݖ)MUٞ�6O8@u_�
�*;�@x؁��F�8=��I�`����[���/�fmmH�v �ix�!���/�`�-��j�P�n�e���h�E6��HoťHu�_P�7��=�gf��a�мӉ]/JL�:	'K��[ϙ�@L�z�MӤ�Y���'�w%Gn�Y��������� �T<J�2�+��@���,�i��s�m�@������	o�4��Q��<���^hO�=�]wQ�NPs	]G���~��W/艪�>>X����~d�t�b�9(��B��&�h}u���{����kY��!9}j����� ���D�J����P#�a0�T���D����کM�����v�U5Pd���hG�|UL���;�oy���������\>�%tEʇ��笮���G��kcD����}x��j�9[�7Yכ�pd�3�ޤQ^♎�I�x���(&vQ7�)ǣ�y��[,Cr�l�`���v�F��l����=���\�^�6�k.� �X�s�p&�xGY�d��Tsy�z�
��`5L�A VR'�F�>�M���Y��f`
뀇��� �����<_.x納Y��\[WJ�m�ӏ�O��/E����cݠ���Z���E颦�3�U�_��#oۀ��ِ]��Ǐ��:�"���YL}�@�GNȾ�v��CN��T�����	�l�Ԉ[y�����lT�Р`��6i�������0I>�r��s�&��r���}�}>�Q��s��Ҫ���_���T�1�g�29���"��9NO5U2f�ov���ռLf!�J{��%��R�|�,X���Rj�!Z=��+cUȝ��B|��D�,����^'P���e��M�B���-K���K������7Ԑd��R�Ŭ��;pT5�e¹�ʅ�V<��o|�lH؄N�`(-l�S��;o���C���s�����v��D���M���b�.* r�&Hp?&�uT��'��}M7�#��4���֪�/�(�偿��SW�+�㡉}!�R�6m��Ǫ�l��\Lq�`��͇�����qP[`�),)�>#eΌAo�!e���:��}�$[Ry��g�������>�t����b>�rힴ���_��l��1+�59����ت5�OiF�'`��q���	�/�O�ٯ����� ]���ʟ.�tՄ����d���#��{�<ve����/��Z�/p�O�=�XD�P�ez��J0����Sf`���l�Ǯ=ׂԐ���x�5@��I�@~�w����/I�����Q;�vP)��ͥ��~�ݖ�rQ���_IXO�+@��˛�@0��\
T^̀��ܪ�v~�y�M"p֋�o����r����>��/J��Z�W#��Q'Z�G(��)m��zЕ5,1�m�N�8l�=�W.����YM�;�Ŝr�JS��EYQ�+�C3�}�N�.&��E������f�g���oU�"�[��R#���M��:1�`ް��Fy)��L��.���5�̎�Tu�c��b$�^H�A���1�k��g��O|>�.��o���IwƦ���6��v�ʶ%3n�{�~��D5&�#\3�,�g=ٲ�=V�YRl��t���2��A����w��4��R��Gd�o"C�̯��nC�;̡��D�Q� ~�X����Đ����>_������5�Y��WY ~�B��.@')z��Wn���J��}zX~�1.����M��� ^ ,��O�Kf��bZ�T[�����ZfB(�C�\�g�&��T{QL�Pi�.>M�[�G�*�p����1�AELk3B
�>P�B��m�?�S���-Bg?�Յk�J`Qo����T2_&�e��Gy�C�
lJ�� K5�qf��T�hmLn�o~�4�I}#��(��Y��,���M�;\z��MV���=�e̓��>������G��p�ț��J�c^K �Q����jh}���݆�Kq�V�voǺ�n>zK'A�El�������z�٨��w$d���6���U��'=�О����0�sٓ��sR)������8�\A� 0q��E','Ol�Z.E������J5wD_U�b��5IK�7���%�/��� �$�ـy�Sօ,�������t�)�-�p�Jwa��K�:'�^th�.� �jvM���Bf��Ym�[H��P���g����%w��N�Ӝέ���Kf� �N��p;v���LD.�.��Ʃ���?}��Ί"�2��l�˽t87z�I�n�
���T����@f< S�>�p+i�5K�I�����îл;������K�0�D�]�ъ,�}�����X���/;PJ�;�H3�yEJ"i$�b�懶���$_�� ex-�����"�-{G��Ѐ�9^��P� �!.ݕ7.yl��?q�7-z�� Wz���{ǀ�rC�>�O���K��]L�@+]׾�R!U���r�`����f��%�H���qj���� �8�_R���d)��p�_��DĬ둝�øz,Y�,^n�_�i.X�Ta��|<#�_�ʎIݜ�wN��<ZWنs�ӝ��%�9����l�w�Ȁ�)�ߦjpU�<�^J/��넽�H"���̿���9�a"�^2.OD�����)�Y�1������-��GT�p��M+�`|M8�4���*��:GcI�˫����(�n�:RN�E�1���&�KT��S������3���m��<��(� ��l��4v�C�]=�k�D پ#�D{�qC@I8��
EL�?�GP��P�G��A6��4z�wc�w�v�fB�D�Ï��.�'��������g�Ժ��| �����ɐ>����kK]LmIw�}��Y`߇f���@��f����<{0�dZȭt�랕[HTef}�p�e����Xue$�HOy���`���`K#b�.Ԁ���X��w�=�mu����Q����G�Z~i6����
��tS:yKy��X�6�Ɠ�<[+��9;����eqc2�y~��n���bSwY)��������`�:���|��E�� 1�/�Ѽ�*������j�V��&v����|����L5�#-�Op$�Yr���{��?;��e!V��]��#�`&Hi��E�_�����Qx�uᡤ�UC2�"�kRg��|�����b"\;�����R����(A+���K�,Y"v@��)��]��F�2щ�U!i��`U�o`D����w��HZ(;c����ʹvC�*@��`jQ�ۑ=ڵ���ܔ��V	��U~��׮���l�=һ��'FFu˻�~�ü��S=�6�� ��Nb�ѭ|�/�_������x��g�<����3km<���|��^��P�r�K<����m�#I���uɂ�>%�R<�g��ϪnP�ߝ������a߶��vGЇD��XW�O�s���6�V�f�þP�K��X�3�ʖ�S$	|�R=bW��ϐs��"|*4�zެ�.��̸ĳ�(8��1��HZw �^Y��|��=^�`��7`e֬�׶�x��1��wn;Lz��P�C���	&��L��⏈���'dY^�T��ԣ1�0�Ƨc����v�-�95��0!��i�!{���=~�B?ە�˛�a�9��}Y��엺R��c��TPk�q�"Q,t�Ҿ�v��´�eY�{�oŕ8Ɂ��BpS�)(\˩ �X�T�_�I�(��'^�OoA��� y��E����u���A���f�Gz�5&&�cw�*�nN`y̓�fԪ�'��Ls7��O�����݂�Wm���$���b-���V�d�Jlܭ(��]� ̷?�|�2	��e�>К���*N#\��;�Ju��E�v�B��gU֝�[�O��i�Q����5g+@�Nll?ߘ���;f�"�\[��Fu�F� ��:q�����NI=c�b�p~N�����[M=cJeᶄ�3T�������1��e���o��:�\k�ԝ�ErAj9��@�-"��"I5V�fl	��z��q�5���N�Lv9ݛ��CmY9
�L���oR�y���	�Wp!I|�ن9�W�5IJU�YH`�]8��ߔ<!
�������%G��)�rm.�Æ����K��"M�� ��7�G����WNgv�iV�̑���n�B��q;��}�����l����M)/�P�BB��+�L�`��<L��Q߽���G^�f3�ɕ�QDq�9Z�@�ZZ��j�J�;.+&��SV�rB��q�ױ�-qy��Ղ(2�[ܤ�60�[9��o�0v���˹�&���9��cM;�^lomOc{>I2� ߌ�s�D��}����M&�� ��YJp���-������E�6�2zL����cS�6����d��9V�E��\�������{ĉ#�=�Z��%l<4�i�V��jh̦3Z��@�O�~pԷ&���{(A��wb�O�h����`hLm�4k��_L�r�k���zbj¼4gZ����}�W>��F��l���Z�]�5�mj}�-0�̇ujz�FuC\d���u�"�=ĸ��k��$>�IO�oN���
{�N0N3�VC��Y�"7�8Ô���zr֚�8d��	�aB2��4�>i��Ob����M����9�_#ߣ����gAmv�����P;g	.�;�˜��.'����o��6��0��L��&�������ƬTR����j����Fi+ �GrZgS��Y.F`��vv���:��ݥ��J^��r�-��>	��_:�p���F0�� �4�՛���a=|e��q�PQA�`�O��ǓVq��d1�c�<�KT lBJv���%��wII6�$7��8�z��*����:�:�~!��e3Tݘ���Ť�%�)�T5?��KǱKѶ�s/;��=�����LݺGu��-�"@y���䭢0L���b�q�,��������:y��V1鴙��1L0j�1ג�=���V��s�9�W�DH�ӹ��.qy�	[Hݙ7�u�K�F�EU���멕����	�B ݂0��l|�`OZ��z?v/����2����Q���eh��f=��WT�n�����!V#I]�,|op���Zl�,�dBZ��O�j��.Ep�Nq��oU�)��"lK�q�9��쓸�Cn��C#Y�ʨ����$�,m��p4���<
�F���]w\C��Q��.Q�E�a5����=tz�s��U�w\ �Q>��,������Mѓٯ��#�<h`f:���?;󁪁����x3�{�D����SBr��	�Bp�����w����V;#�
=�[�h��G��J�|�7ر�~8+��KD����VR�[g�|��%m�4;,3�ԉ�;>e6��٠�iG���˗!=رs&��䷚�!e��$�����Z���7��s�+�kh���v_�����EX�AǣT��T�:c����'r�7z|�T�9ϻ㛫�����X* V�̯W�9�a���;5_sN�x�_���8TjF�iJ�c�dщ��X��������qp���%��e��]�i'W�."K�����2/�*5pc�"�D$��v:tf-��m}��֫=ꇈ.�q#�1y8۹��G_ҍ�r�l��Y[�?��/�
R����4 l<�*%����c`�pnu��:t��J����k��*����H�$�utG��=���܌l̢�%�+�y|w!k]��M���W�Y��������g=�r�RA�b0Ut�x�9eV�7"��w �k�s����áB�P5(��Ǻk�$�ג�g�3=�@�??�8����.���g.�:�T���� w8CmOWH&��x"9��m붉��Ye�ݾ:t��ȣ�^�!wŮ�Y�ٞ��G�p�b��p��9B���t���ï�dP�N��(��l��\y$k{
S)�nR�����p��	���v���w]a]V�>Y"3��� U2{��j(Lv/?}i���s�Ȋ ��IWI_�u����>�h&���bM{MKik߾�qkț���$�
A%SsS��"�Y�������8/^����	���pP�=0w9j[J�vO+�e�	��
�4�I�$���	�&~�N�˒$�ܕ���:���������g
5����䲔3\���KO-�O����$�����.#�o}�E��MP�L ��B�?�����z+�W(Z���$�?q��nq0i�#!�	%��j�ga�7�?j3g%	�Q�>��5{��(��w�Ge������D@pL�Km�yH���8��}<E#?6�)��U+�w�~!-Tj1�T��n��T!�I�@�z�=��pe�L�x�Q�<��e���c�4�����r�2ՑJZv��K��e�[3�ƈE�}x��q�Mw�����$�q��������߄�~B�4{��WϦA�wl��="��J�n+���0i�[�un�c� x��CC�Z�+㗉������
5��w2^
A7�R��}��Ps�z�=&����H)�[A�}�@8h'��J�b-!�&���{�~�f�N3`݄ڕ��#Ͱ���� �,��/��~�cx���P��s��2^r��eO�%�d���R$$4_��̆Im�3P�~	}^�$|��N�o�G�$��T6j�8;� �t<�ޚ�j�����"�Z�6(3O�m����PF���u���f�	���ԩngyt<	�/��+z��"t��� C5��5����J @�Z�[�ت?�0�R�E ������[��yk���w��)6�)�D�F�W]��0
ƃ����0C�!d��͂.�C�FX�Snw3�xQY
k���o��M*d�$'�%��c.��p�^��k���^d�̦������Ynͼ���Z}ؕb��	:�2&�	p����	�� b`����HF��x>�2q���v��e�U�o��!&(�=t&�0V���ñ맃r�-�n��Ct�b6XE ��<��Wa�o�_]s���v���y%�̉��U��i�H����9a.�W.mS?�|s^ܖ�e���`D�ǣH �FĐ��b�SǑ�?�32E����̪�![oXM�q"���\ɗY��-����V�wEjˆ���_��������7�ru<�橺L�w���;���g>V���0�MK;�p*��ie�(2���Q|�o��z�\���l�W3EN���<����Z�}m�B���&'�S�����e��E���t���M�0	�.R�.��hz����M�nAB�<A ~N��C��>��Z��n���Jd9�
�,��?g�������hj�'3��f���*�%,��t��Χ�:�|���~�2詨��B�>�F%����,B�xt�I��� �
�ۿY�O��_^��)��ڳ��NބA�4-��'�Ʋ��Ak(@����l/[!l�C_;倓l��Oxron��5a�8dPR�������@�6-�w�
i��q�D	��o���a����U����?�`u9�@Ze�rL`��:q'}5n�c:���Y<�tq��j�S�����v��vyJ���6_��
�`XZ��,�b���aD���@��p�w
tmtU��lh"��F��2 �����)�r@ ��2K��8d����}�{�J�����K�ފ{�y�R<�R����Jj�������m�&���Lt�P6�sH��M����U�*�J�".�a�xY��Ε�b�֠PiI��&��-��2/��K��n�0�j�L�DK��w��O+k�O �U�r>��Co/h����A�S6�����b^�m*�S��5T�3�;�o�|ͱ���o����>욚<WPƏ�i�~@�<FCϳm��2�- [�l�ޑ��uEp�]�%�a:�u�3�f9���C�~�<�6ϳ�N�W$dt}'�{>_�.��Ş403�8�(�+�_$v�4��#PкU@��`c��A\���uw���M�{d��葒o��5ï���n��o=z�<��� �ݥ�G�H3Y�a�-�y<����Hoѕ��^�6;}����/��d�s�^<��1K��ͺ<F\D��A��]~&�C��K)%�Bۄ���㴭�����M���*ԃ��{�^�U@VY�x٫�P1��֌�Iz�ۼ|Den�6�0x�qLW�W\��~O��K���<�4��Y1'W�.1��I�����w B���V�]b^��P뷾�!6ww�R���.̞]���!"O��(��qM&H.D͏(� (�Z��r6WЙ,��KWoˡ��a��r����
�m��^�@)�}��P��n���~aEOր��Oy#=ނ�7��#?2���T#�.}�P�ޣW?8�}<]��x���ǿQ~�wM���/ 1���[��X����X�[�I�Z.�_#`m��qݐe��{N���e��{�W�JP�9�3W_"��|,vB�G� ����~�2���zE�o���g�]�������5���:[�8���I�B��Qo�ʘ�>�Bgf�5rW�#���U[di$F�k_�2��AD�3qCz�s���آr�d}�O��s�t���Ԗ��|:,o�=Xo��| � �뜹J
��^}`0[h�+�d�W��v�ER�D����8w?<���Q�Jl ����Aÿ�6����1|ңO���`B����(�8��k�)�jL
�/R_+G����¾r~�����Z
Ɩ/�w�f�*��-L�ǷT�t���J���������Qw6�m��a�#���l�M l�;:#�����~$��(b�B#�醌�]�{Sk�W���P>��Ss]�;bTu�=�jҋ�a�|�����k4'T(�U�yf!mF���í�;���I�U9��_�Vi
�]��&k<�7�Z/d���y�`��a��9��|kV���^/���|"�Wޑ3G�>TZm̊�`>�0	T��w���L\�/��rZ9�%�R�GaM_�$�y�S�hFg@,�N����Q	ה�|o��D8Q���6�&�+
�Z�Rf�5�F�;&�s���m���PR���� 򩴤�4����ѓ�9�6� r�*�vf�AagX��]$�ի��a0N/�>�6,
Ɲm�lϏ�S�d)�?	R�1IY`&���l��#���ڜ!&���Ճ�l4��a�m��b������]菟�_j���?��Уc�𛞍�)7K�$2��r��Z`��[���D�V �1�Ҋ������ʚ��ۢ�s7�
ǹ,nD׀V��=;�h`i���
��1B�,�A!�-EQ*w�D>��u]�b��S�����%��E!/�ˈ�bm���G[y'��J�ȞS��&�2pM����Q��4���&�ʾ��,6���^i�dw�`����~l�E����P|�/h�>���6��v�.�t��gS�Hy�M	^���ǔ�RJ�}����+: ��+ɴ@�aDhT����3�!�����@8�_g���B��dP�/����i����?6���r�K��ElK�9t� \y����ź���2���e�fW��_XvA:%��b�j��2�>���^]�ć&�WE��t�Q����()��8�9f5�

�&(M�`4���)c۸���K!�$fd����\w�^ޫ��_�u�8[��dh� ��{0����\�;�3�<�~6���%��9�7G�tdH�\�Y��ı^����%�ђ��\͇6�����.�_�N�q;�XM(��s�Veݎ>a��[A��."u�(�(qZ��cAQ��K�*�2nc�G�eG��Q� ���Ln�Ȓn�a�E_p�@�����D�Y�L9�	(���M�Y�f�F�P:��n����7;�Զɱp�$��HJո�[�P�.�	ˁ��$\U�	��#1���$k���$��B�fў�z5A� c��Ұ$��'Gz"�R�*����f2}D��Z߁q�|��ɘ�4���ϵ�!��:��<��'A��~Y`����c���h.�׏���8�/��l����焧�����;�M���} >sBP��v�0z�ӣ���TK�f�uYz<T��Ծ�2,8���<�G�Ɯ�Q�>�2ƟДՒmL8vj�p�#���K����Vf�B��E�`���8�������R�)ъI����=�I���0�/�R�nZ���Ԣ��\qj��Vnתּj<_�çM_C�y�=ր[�R5�v���|�`�q�m�BsI7�J��\�c�إ �1��Y��6�z�!��E~�%l��r>��Y_�
Ŕ�
���)!n�-%D�L�pf��n��m��uy9�^u���qT]�.��HB����/�z��l��G,��3�^�7�	Ǭ�5h�_vr$��g!��]u���o	�F��Q\s<J���W�M����1jf�l���4[tь��R@H�\&�f�,r�� �S��<7�������dX�:���|�g9�T�}�\�s� +L�1k��"/8�\�.Y��U��v�^R��̆��x���sML��Xx��RF�ꂛO��H�����jJ��˾���4��[��(*���_ǥ �?M�~?���3$�2J�+Nv7���igR���=���]���uF��^�1�N]�������F��Ћ}�T�P�t޽;*��h�5�@R�$H�L��c��[G7�H5`F'��I:D>�K{N��=	Fe�\��j�H-��.G��K]����v�����I��	��Z���f6PEʃxX*]�� 7V��ѻ�V����7gq���w�";*����[&�*�V�����/ؖ��~#���\O Б�³��w�ȃ 06Q����7���y`�|��a�+��ӣ�H,�ct�0P��n�^')�t�:�{j�?����FᩎH�a��W�H!��d"Q�ow�|SY��:���.�[�O��/�4q��f�G�UECtj� ��H}�|��qLW��@��l��G�al�I��Zje�5�_%�I͹O���#�ۢ'zZ�{��b�y�]�C��=�����>%O������ǹ%#(z��h�z���	H\x�:yG6��]cpa�����M��(���3��ܷTW��`���p����uI��Zs)^�H�5Ӣ�a�Jwo��Һ|1�߃�i�ZU���V6�H9Z>����J�pg�#�"ć��]觡�8#~��n񶋾z��{#Yi�9�"��${I���D��Ҿ��"z���sX8*�b\)ț=�P"��]7��p�A:0Y��@�4p���z����/�-�d��I{�������_�֬�_|:���c	��67�t��s�)f:]��\���5����2��WŒ̿ap&nt���H�A��r��u�>�dg�y"����"�)�͍��^���M�Rg�#r������c�ߣ�P�	�t
��Cئ����ޯ�[󫚔R������1[�t=SB��H
�d�i��Jؾ
 ;�3�Z���ƃ�1����	�H#������p�M �h����`���B�����4Ce��������I�>Klms݁7}�\���Y3J\$
�/
\]B�pL㪀"Vi�2�w ��/��A�N�i7$���Pf9\�s��vbuK�E���q�-p�_+%� B"�1�qE�I-�u%xډ��@��AZگ�]�m��{T�x��SE5��[��QH5ւ�Ã�!�$�{�&|�o���ߙPmwk��2TCy�.�F��JX-�A�,���#;�3W�Ў�DH!���5�T�jبG�sf�'8�4�v�V;D��%q��dx5��S�h�D����CE��E�:���(�uJ��?�"mS����#슟e�A�w�x���_��W\~� s�����>��G��f�.��8���}ӏJ��Gk�}ؔ�oLƓX��{�������a��S���9�^��}���Un 
dRp���Ǆ�ܱ�h�Iq��s�U���o�tw��'���4x�ĀY��!?��@���ͻA����d�Q�_������%e�����57F爘����;z�9�J?�oPc V��F�O��N����㯮�� 	�R�H���#�E���<QZ�~�r����pz�X�T����fQ�w`q��$ Eod3Q���|��VKُ� ������$%�����_�;�����#"8A�^�H��Ff�p��?�*i�����b�8%�F{������ۈ/K��1����P�ᫎT����mr��z�������J��,.��C�D�陽����a$
>���5`\i�J��%Ϸ©�(}���L�� ��ͱ��_���s�t�y<�ވ�.m��P�P�>ܐӺ��
��tIN�{��PIE�l/IR5{��Ty��OJ [��}��1/=%����<S�Mj�k��yN:\�'v�-�FȖ��a��}�Ke�ٚ9F��ב���bn�`jd��!|�B+�S����UY�)�O� ��k��ӧ���y�ι�҉1�I�͜�$�̳W7Tv�C���Y���Ȃ/�`5*���_������[�YԾ�cHr�F�X}cʹ���=l��#n�C����3с.��~[�2���f>�'.jL,~g��;y��GYOZL�2��^�����0�==��Y�8<��,�f�<��k}��5���5a<�p�?: ���B%���x�8P1LI��������g�+4��P�����t����=���=J:���F�>�j�M�������װ��,ۭg�ˏ��͌���d�G��E_?��y��n�����d�rE\]��aH����|�E�^:a�~u7y	S�*�ޞ]��G�m�Z�T�������'��Q%w�C��M��LF����G��~�D2b�yG�ԧ�#�i�n�����
�{�r�T�S��?��3Ş�B쯛
�j_�������+�F���R�l��*x[`�0�a��|���1q>K���w����F��͉��ا���
l���i��@��J�fʒ�4� xA�����Z�P)�a5�}�nIQ�3'FCaĆ� TSvW�&�-�%�ms�%�oq���y�� UV*�#�9�2V������G��I��~b2?����O����!j"��6�&�鷮������(H|<0F�Oͳ��؟�E�	!_�rBZ�g���<C�A��nx��ZDpq@ �	O��g8����Ǌ���A��òP��K����)�%�u��S:�c���$&"�Ɂ�8Ɂ�����[*;�X��
K�p�b�T��u;C��4�H��L1�����%,�15��3��������2�4�Jnu��w���1J���+��#�/>2s�<DIS�<.Kik�BG۳k�soV�e/:aW42~JX��JLK#�5��q�7����_�A8�0A����\��p�lĨ�`	����ذ=b��ލ�	�q����uU���z4�yܠh@7j/v��D���*MVI!�0�������d��7_PR�޽�D�iG4��
2�j[����D��V�|�Օ��&��i� ��>Q������S4���bx�d �#!g�--2앀��r҂@�s�§�\╄���wp��}�����Ǎ�7/�n��ߔG��� 	lWb�mlԓFTK_N�wݓ^���U�5�-#Έ��pM1���@��c�D���^�@v�{r�T�P�"v�1��]_��z�0h*�@��pS��7���j_���X>,ef��,�z��Cx2ճ|-�Ad�787&p��M�dU�+�� ���t�?�o��M�0~�.�\v�"� ��Y.��Cz����M��G-S^�w����|
<k�-=yH�.�ع�K�3�.�Of���R����+�1ǣ8*��&p��;k��*�ܢt� \�]k�s)�M"A�z��<�(��w�����ɭ5�'���gu:�O�p�<�7�4��b]E0�EX�j����ׅ�F�H��4*��n���y=YX#cU�m�/��V��D���U�'��]�(��Obj)QV6�l�x@1J�����Hvt� w��6�N
����)�3g� #�e`���v�X��y�ŋ�����{��r��{o���e��>	�������|iQy��$�������\��-ur�SI���-�J��-3&�\��*i��.�4�7��.���g6
	�� ��0�DT�Aa��o�f��5ƚ�G-��z�}u�%^w+4���,��7��=�L+�u�A�>� �g1bE�{�F3fX[������N���F}I�X� ��ж{H��Ģ��S0zQ�؅�L� º�Xx�kT�y��|k�4t�[�&�����k���>�1�4)'쉆�}���q&��]#���#����囻�^�H�a'>T6��:�s`�d�"�qfFK
ة����߭��]�5(p�����*f$YkLS�a�b�M��ߓʲ���yI���Q���, �[��i9��/���Guʻ�^.C���֎V�C[��pJbًQ���BSV�	DZcO�������;��9V�e�bk헺�p�0�m0#�	��Fۢly����9dH1i#˩��k6�x���Z:����ʖH�l����Wg�z����4��O��C��➇ab���{�k�Wj���Eꛨ%������:;�0r�����5VNҔ�F�B�M�O������ae>JF�&LE^s�����z$�k�C��𞊀� �e�:	��}���á3���G3��6�@wq�҈��K0٨B�kN��I�z.�"�v��t�ḏ�Ch�K�~�Tgby����kj�o�q#̓2��2�N|혂ˇ-4[&��R�Cw�>o�n�av$<�W���^ջ�R*���x�C�mL�-Gs�N��>�vAl���l6= �s�$d^��h�[!GP�Xw�T�h�p�F��!�'(���J���e� �����7��Y��^6�ЛIk������*��B_Ka����ȑ�/;q���A#�G7B��S�;����'�H>u����f����]�kd�z�:�V�0���o[#�$�_���@�o����WD�=��S��eˌ��vԽ5��(6k?�����v���m�ƾǐ
Jl+~(��/v&�C��OC=�bרK���%`W{5�3�~J�$P9)@J馌N���9��z@��r;
��\/��ధ�~��q~�pJ
�%ԋ#�1u��Ʃ�*���>�<5��n_ϟ�_LX���k�DJi�T=���d+�����Ţ�_�����W��F:��*s{�q�|E#�HX���K�(�����O�/X6%V;�F�Y��1����7^u���N���w�t�{e�|?�����cjaho�1�{.�4L��ⶓ�*h/I��B��A��y,I��1]��'��(tI⩪	����ڞU�0r2�������R��i�'t�U����RZ����휻�\�?i�O�Q�9���Ә'��j��&�wo%F8�L"ô���WL��p%~=�vJъ��U��A�z�qt��2xJw�h����3���;êbXɾ9�t��zYnI�L1h���Ņ��E����I,򕽗M*|����K�Acg�뿣B�>���&bg��2$-�:�<�m�[Ƌ���I�(P8���tPo%?���ͳ�նN�8���Zy
<á�1Uzp��Kh���p=�}� ^e[O~%�cfmH(�Lʅ�T�O(c�@�,��wJ��}�_;����E�XR��@ķ��B�D+S��t��8S2&�z~n�j:j����y)����٠�4�ZT�B��lY週�������%�8�������b:��}j9SK��}O��l����5�|@�0�F��f�e��²�[�#(H��X�����?�5��MI�'���F��v
c^�[;��N+��xx��|6_q����Ң�Ѭ��`1�I�����e���l�E����F4�Tj�=�>�5��Gr�KNo��5�KG�{�b������كJܿn�	e�C�;+`-?)0��I�(Ђrƞ��M�J��\��?�u���3�ɉ���1�ԯ����]��6[��#r�Md�׊����JE�8����1s�Idi�v)jD�'/�}�������4�}'-�PT���VT�p�^���|MQ+d��W[1G�~��H0*5ӕ_�\�h(`::r���y�!�+��m2��_TC[n���}������VJ��*mXJ���P�Ή�a�D͙��֟���~.�@CA\G��Rv)*�`V]ſ��=	x���iѿ�@����(ٚ�����ӄh�M�إ�!��4hň�f9H��ܦ�Lw�7���j�MVX������Lޱ� ��B�4��J���qu�{��p��\���r��e`�lH㚲%|x?�2%��B��[x�?Jg-�A�M��&����xU�V�8�Z��g��r��[�9̲�Ejj��ahƢ�4/��TB3�G���T�pt���g>"Y2bj��p@Q �
��lغ���(v9W���@Y�u����K{��@�д�0A���ҳk�B>ěW�� l�d�E��f�X��%��h�������
�.�H��|�i9�Q�9_:i�b�� �mԭ2	�7��d!L���9������oO���/�]L�ߩ��Bdm{��	<?wA���l
���A��Ps�.�6@�����q>��m��w�0� d��`�U��q����Gy-�xO���"Z��]��PVms_��"6�Mþ�����g�J�rׇ7�8m7P�k;�����������/p�3�c��Z�q�}O"���4"R4mϓ�.Qg>�_�������4�J�	��)Cr�|��1ڈv[�Q�r(����Ɩ:k�~���R��¦a��VH��&��BXo�郊L�h�<�d�Mǭ�W���BiI����ԎO1L��%m6K�G�y+�G]��8̒��-����
Ȁ߷i컼̩�m�"KZ�{c"/��PG��Iv������dAJ���~��<���S�ȣv<|��"H�E�9������!�^q|�����O�r[�J;���kn�)��hb��*0=���!Zmpy��sA!$��ӡ���o��%9W4��%���[���z����jT��I�.��۳��ѽJS� A[��n��z��9�yn� �,��#�I}R�e��n!ƶ)�+��b��2��9 �&u����Z��Vٯ]�z��;?ώ?L���,UY�2Pv�m	UH�,47���)Hˣ�hV����$�xwk6{<��пt�����6�$L�[������v�d&ug)�%�ѭ�ŖD���c�����]	��e9���V��:��uk�+�/n�iW'a��f�3�.k�.�Nz�yf,Y�Ρ���|k&4�Y��lƀ�6t��)�"���i��{�����@������Џ6�"��d�~��K��c����(|�a��C����OA�3��ci#RvRp �^���)��'�:z�+Vl!0J!\7R��\Z���t"�P��2��fS#�dnzv��Q�랒(��Իq�l� ���,p�8g|�x)7&ʿ4��Ta�*�^��SR���ĥ{�a]���/��L_.��7:���M�4�s(;Ee�.�P7�8�(���\s��ya��
���ԏY.�H('4Њ��b�"|mf����tD���tLاJ�l0���zS s���
׉���������)�a��~�I�t��QԠ@�O����zh)��L�WD��*�m��[=?��K�
xn[�-���X��H�3�II79o1`s��]P�>Q���iQ"�u���ݸ�r�YuV�n'�yQ��^�Y�PˎRED�z���uxr��}T�W�e�}Kny��U�͑
��n �R+�n{������y>c������� �)�9)�Yw4N'�crvyP��1j�f������1�K����yu8"�nr�fp�bo�'�t^���:��*���}�QQ�;��j������U�IV����Z/_]�;
�r)5����`�@-�V��1��B�T$Ts�4o���b%��bQ���:R�尉8*���i��@ZH�����`EKh�d}���������F@|�(��G_�^�}K0B���������ޏ�v�5 �|��� �l&$J'��@�N��PGh���s�P;5���*Q�9<1���YY�v�t�GYq�ss�pVP(���R+�0ғ����N�n~9UqbE�,��t����~��a�,f0��.63��������/52v�q�F���UT���n����bo�R�BDoA�%U��E\1p�����Ǟ��n��}W��:,�陃)z��`o����#���ww���1��o�V�����2iU_#��!��N�bK^Id/��\�#/��@]�r2�@��X���^&ou"4.���M]���_��O��zm	V�5o��G�}} �S�J�N��B}c_������c-|~�p������I��ԇ^2�@?ܞ\9��$�Lyڏf��~�%��`J��XR��2N��(��S� �~(}�����S�4���A�4��������2��f?�V�F��.Ú�a1�5��Ց�p�8,�A3��_z|���(�ԱE�ʶm�����M'.DP�ͱ�Qڋ��������*��L�Qh3�x�1�ᩘ|�#8m �K^غ�/-ߔL�= Ma#�c�x(atpf��xzɁ,$�6J{~_���t"x(��d�%�,��ԿʄSܐ 3l�Cg�uP���+'�')�E%<��+libT�VY�t�Z��q�Q�-j4:�c�_��,�	x���*��Qa2n�0E��J¸�"���{�} egYp:ķZ��qr%8
U��=Ҍ�8m��މ�}���M�%Frnx�� 1�ڲh�Od�{�`�[v{#�\����ONNi�G@(Az�7�Z�$~�Q��t�`�; Z2��,`�u�X�OD�ׅ�!jlS۴��B$�����h",o�s䗤 �a��t�,N�@P��;�b4`�2�ӝ������AMSg�bd(�����P-w^Z	p ��ݓy�i��Cį<Ad�Eu�|-�<���X7�uWw\��yj�Q_��2��0��<ȗT��S�Ν���c`�6+l�$��,6�Cz� 1o#��+,���1x��p��pc�8�=EýA�2�p�����cռ�Ro)M��9��<eJ�����=�¸���/g��V���Б�L(����J���(�Z#LdIp#�5��&��_y��&��ئx��:��u,�o�n�+�1���i_���u�38��ǩ<�
��ѡ�+��G�n6=�·�\T;��PN&�o0ە��^���}9#�])v���e����),�v�1���h�!��K]N��������� ��!�g"&���o�y���Ѱ��E��OZT
�K�+��T�=�+�tn^�z�Z��l���y�i����	�	���v/u�U���Aof�R`�k�����%�P.�bh�9�Zgj�MA�ZKI�^��"��Ƞ��xN��`���ӬP��++�
\ጹ��B�ʎ"(z`�9�K�_�58��k�v&J$�k��д-E�g�6�뽿��9��7r���Z&9w$�a�w�P5�Ktm�e����1�  5n�W�-����02O (t[����t]!��#��O��}��A���k��X�g����`���҂�g2��~UE���Df�Je�������!�m�|u�Y:k: 6;�ޥƧT��^_9�z�����xY�*:Rϗ��B��[�dV�ϔ��a�ؐ��LaL����SA'C޿avJ2!��wA�޵�%���M��x�#��Li�ϊ�I�����)�A����A@9���h�^�=��A��{��kF����Σ��㟀���*���J���+�{vP�IY�3�uY�D��m��Sq��lt����ո�����O��`J؉��<��Y7T�B|�@fj�RQ�d���S1��U>��O-� �Ju���� Y��e��c�Z��S%�B��k9ܖf��5yuv��h�=��Ką9JZ��	˶Vl�n9>�$�K�`��
ϕı�F�4���I�	;6�I�Z �1P ����%��,{;@����NPI���<y8;���^[o�2Y���v��$K;��#��#O����z�`��wLb�T��
�'���+
�.J���e8&-r�V8�2��]�!�]���g�<]��P�ǝ6��#
��|2wK�>Sxj�0Z�����t��!��䓔O�$��c,޷�}���
"�l{�вy�G�҃bj��k=g�NP�X᫡�SZ�����j0�fC���?bJ�Z{�
�"�yTDڀ��!+;���3�������i�_��^��Q-��.����S/Ѻ�9�f�dg�P�H���;�,^*G/m��e�7�ڎ?������^�-��:�o��`�N��J�UR�}�N�幌h���+��2Fh�)��Z0�O�_ExY��Ԕ�!�{��Gp�-76&���.�Rh�K��܆�'�$VH��aztke6�4�T�T�	�g�����e�O�I��3�ki�4R�dy N��6/��i��׶7=���?׫�4Zc/mB��pu6/1���ѳ�[`�݀	��Z�����@�Pj\yH!͂��gF�7�N�J����M?lM7�b|�i{qz_�D��HAz�h�0���_�;�u���葆bS�9
��o�aW@�"�Fi����n���_��$AZ����6hǪw}��׈���w��<�7|��-�
�9�Q!qY�f��K�a�Y���2:����K@k�L��,����/F����e5�st$�;�<���z��5�P=ϷZj4�<����Kgl�~s�.f�)gm��?��-�<`/Z����7�t�Ry\���Q�R��[C�Cu�Z���HYϫ��ve�/�s��i�m�A���r����CV}���^d)��s�HP(�l���"���mO�kV�05��%
�3��]A-��_\�`��u�>ZO:BY\��P����z��+ѱRrw0�#@^�&1$�>?=�%p�l)hN�U|{��8e4�����244�C^��L�WNؚ��ܨց�|�lի��:�0��|�1.�Z˹�n��`�A���D���h��G��2�0H����U�Hq�CUo���RS`Z�vE��Gr��m�*�>��6\6��<�:�U�ےXVE�%��"f*h�d��������d p'�3g�6D���/eƊ澉nX�灸�z��LAY:��d������;�u��:5�'��m����H��P���cYz�o��>'�FO}�ʾo�|YAw�Yި�{��O�JRC/��(�u���v��t��V��O��#	����=H0AR��T�[��<#Ĭ���M��`��/Chݶ1��v�$��S�<��1-=�+�v�������j��WL�Oe��`��V��:�l�ա8�y�U�O�Үq�J;�H2n_�6u#l*� `�Ɓ��Ù��έ�>��+Tu6��c��=����<1MY~"�� �<�f�|_��ڶi���vv���]�FC�I}�E�(���]� �:��%��
����=kC�B�E�V����{���q@�[���<�ks�I��H&Ó,�!�����V�8:�.�$������cać ���� }���u$	�K���9��R�j�Es%���#�0T�F�fЩ`J�M_�hZ�����,.�gf6;��y~���x�Oa��%b�}+�
!'�����\Nxp8}�y�ڏ����ZF��B�C�)y�Dy�}#���*/3��~���K�*�ΖB�6:��$#R�Q�qC4�[���Zge�]�3g���!����Q|�I��wiY�UӜ��Ŷ�>EUV�=�� ˛T��=�#���u��\�>�z��]	-�c�v�}��';5i,�lpbUt�����oN����}i3)�� ��+�FI�2��۴h;k�A�����|�"��XټD�hx.��)�v�a���Z�.�5Ns��i���.��xÿS�v�3ǰ���hie����Hɽ��%�pSƫ���r#����x����>�	G�������q�i*���ɰ����Ͳ�[�o�o/N�%\�종Z-V��+4���܊�^��bX �O��Bm�����^�vz��:n`�T_ry��VJ\�|�y��T�m�� T��WԜy�\QM�����SR8�o��j�Nw��5/�a1\= �J�N����PBn*M՟W}�pm��Յ}a�?a�hb�v!��8	�\!Ǉ�$�3��_�d��7�`�Ɓ�\�|�홸��,��q8俶d��m]�-�*Z��|z��et6]QqC�[&�)2q����m_�S)cn�����D��ENdB�^��h[�£����~�63��n�U�ʡD���{���eH��Kd-jOT����L*�77��t����ϝX�ߺ�zl�W�~6V` �L��eGJ��V�b��>bK�F&n1J�� Y�x��5plq����'���XKԱ�#F�>q�����O�*-�O���UH���X���#]�O�sCIթ7�Έԩ��P�n(�l{�g�-��'e�Ubtk{6?kg�x&6P��T^C�Ԡƞu��D3�8�.`��S.b�� mq��?4�1��;g�2�� �?�Ǟk�rMn���\�o��@��z ȴ����a��v\=:-��_V��N5��=>3��`q���=��]Y�n9.H�w;D9P�ŤA���៴�X��� ��/���s���/P�� ����O��^�(��9��i�#x��3�t��C��f���o���W��K��cը��.*�xY��[�U�p$@����P��\�DI���J$��~�
#�����4� �U�8Ÿ�ߒ\�S�{X*�=��<��$��Dp�_s�W����Q�
�X�x9��m�N��o�yFD�>�"z1�⁘窜>=��v駻aJ�>�]����Z����̳��9�%2�'�&��r~��_@2>n���W2ɝ�����f����u�1˔r����W��o�"��`~~e#!l�c�B��35W�n��ğ f���;���� �\A��?����H�S;M��^�-0�f���[��H1��ƌ���\U�~S k�m�"ӥ}6��;Yӭ�)kG-�\e	� #�|�
���x]�-%���_���(�s�Sp�۬F
An:<�:�7'ȁ��)���6@�U�.ҝ�t�C>�N�S�rU�)/q�ȷ�.<����'O�c�97B�.�<^&u����GN|�ї� n�Yu�Z�ڮ�j����w�����F/פ�ĺ9��g#�wD\��
������������ ��b`���T�E��ޏ�g�L��ڌ,1��0�Q���ɉN���i�Pi��6���ȋȍ�t{���h��q�OE�[Ji��-��\�0����i��U�Z��+a
�
�Z;�1�K�N�,�驇��Pr�	d2�o��{�s ^�៾��4sh��"��1��>������q�|�0>[����G�,2�����O͍��P�`%{������ʍ27�Ǩ]���Я����.bg�h=�7���0ca�Bg����.�t���L��Ĭ0�����]z���EQ��	M�F���$��	��^�1��� n������g%=ߺP4:�_�w�<�w��h��)�{v6��iX{7/Ef��}�3ߏ J�
��8.�:���7O���'�B�Lj�̵�`�O�v����!�*\��$&�)��]|&]���z��8/Z�� TΉ�4(|��6���E;`oiپ�ڲ^���a��j��ۧ�k�׆nl�s���b����b�g��	8���o�� �:ý#p�p-&D����y�5y!	�G(���i��p.z�g]�p�����w��v�(ʯv$=3E�*Q�>�h/�������NW4.��
C�{��]���������߳��N~��svˬ����oWW0f��,���<�a�}��Ĳ��9�,� 9�7��C�����ߊ���.Ε4���[�K���� T/���]"�^~�r��~|�N,`�V�k�~�>��h ��B	�Av]�	����g��02���gY�A�!�O� 1nW�(��T�_���G��F��Z1&����g5m%䃲��:�,h��/��0@\�ӹ#��.m�ʄ�{<�3qqޮ��k�C� �$�m{��?U��M�:�ʌ�L5�\���Qɰ��o�}g� K��%WURH4����G`Th���)s c��Bˋ�w�`��A����ط���o��<���ur�w$ES47�&�;�d)CI�F�`����,�@�}�Õ�u>f�Cı��edn�^��M
�M�'�%�
`��cp�
M,h	R��7�:f�W�D�*������h�#;�-s#��IY_�5���� �jR�ž����	�����3�eP��<Ȝ]V�Y��'ḷ6&�gz��a�A
�,����՜�����&���t�:|h=��%�H�	��#̦7ϭ�Е�������/z͕�b�����b���5���&'/�D��|�/ ���V�8�%��'�c��{�s���:|ڵ6=i�ܙ`Ik����݉�x՝/`z�Vjb�V��p��o)wv�ݹ��h�}r��gG�#�6�z�z4%gk�12C�sw�%�����I��N��N�����Y#�tA*�q�+�s�!���nD�`��c�P�}uM�ʹ]�cxq|�I��8��RF�ъ��*�5�]�����+���&b�*<��d�oo�ٵ�M\ɼ�th�"�b�<C0s�H4�yz�o�=���)KfL��(<���4�(/�K�&�X>ٲ��<Ä�4�-�#�f�-�D�-��:D�Y���25�5̪b����omvn'��궈�N0<���8�
��_��&�.v� ���s�.�|,EbA|�M����J	x�:+�vЫ��@;����I�|�]���`k�fc+�4gɂ���tXLk"�p����a�D���4nYq�A-��F�ۭ�b�4��@�w��mJ&�s)�S���'�F.��U�*9ɯ��y���'E�)ĵ9ᙢ7�b�&����m��/�,�cݩ��+��b��Y�\&���\F#jL��vMќ��XH��ξ(b�����(����4�E��_~�T�QQ�=6���;nh{�a��SA<���2*C
�{�t�@��R��F�}�L깊�B��i��d�~F���g�8�xM�]%�W�ȝ��ݓ,�%/��=O0Uc�|�]{$}��	]�s��.�I��_�S�}���Hb|�wC�zש�Qt��9G��N�^��W����*�Y2�8Dmz[%+B���q~}�`\X��*�!��f�Ӿv\(i�7(�eP��<+g$V�yEkM���\��3ϰ�.OQ���i�،~�;��0[�O��ᡲx�O�zz��L+��)�w�,� ��X��% ��W���9v�A�xG�k�t�������RI����nd�e�����!��c�b�y	���NI���"��\�'e�i� *�	j�r	�{��H_���$@��e�6��`��<��7.���pٔI azm��;w/��*�����.��S�g��e�5�A�'�Q���%��&�gŖ��G�#ӯ_j񩕳y�;I�d{	^��1�RH�{��<{=Ai�O�#Iz_Op_u�5'꺻�`��O2�5�!�E?�z�A�����1<�i
�9��?� ��]��@���)T	�o�͞TI�æ�ُ����Pc?0e�����1�g%TV��1����9q?�~Υ��3�I洆Ex+r��S� �/�R�9��=2�zJX�*7Z'mo4z�yI���z�jԶ{J���*�EO���a*�M���nh�&��2j�A7~��Ő�!ïABk�t�f �@&��t����,� ����ѹtF�}y8�E#��up(`5�K��g��?���a����Al��X�R3*J={GFz�5�����=�^��o�����_�L��]�v�k����r]5��)sS��UU�9�SY9��(�̴,S��hv9m6IP=ɗu�C N0�o v���m��g��%�<�N��|�J� ������}��&u���;�]��$�Ԩ1#:�Pj�zA�(�?�ڗ��A�K
��_1�Q�� ����tu�����DS��#�:��t���D&�Hh�!`h�F��O��@K�����-���QO�5"�j�5��8-:vQ�@J��6�̲����(c�Q�f�mן���K��"����^TB�5�r��:��GB�����cӯ�
�X���Q���x�γg��E�A\ aZׅO8��\8�Yr���
7��/K���!����z�I@�DOc#�=����("Y�Nvm�&p2)����]�{�J~���ζ�߲���
���*�FgR�7��W��s�Yd����/� �-��݇2�-&��~㠅$ފ'�=2�z�'aǂ��j�����n~�s :c����@��i�,8�M��z�&��"�S�.�J{Ok������$�%$Wߖ��[�T��C�S0�*\:W��:i�&Z�_5:��CYK����?����B���y0�P��J��j���|�_l��DMMϺ^(DPn.�.J��@�fd�׺����dҋ��W_+��p��K1a<{��W9��d��,Gyac+
���#�`�5I��?D$PB�Z�H�ZZ��F�������6�K=2�_CϿ�k#�ׂtU=��U��F�Z��by��@��K��6Pz�K��w�V��׽�y /� 7o���@�(�.���R��֙��>>˴?yV����"�j៲Gj�/�!���1�"����.\�>O�Q��t���e[+��-':�:{��@we�R$!ĭ&K���}Y-/�`AR�����)%Ց��5�I��&�G�D��˃&��"S������,�$��°�$B�v�E(n��������þ0�ܨ+S����@®S���7�j�Kc�/y�:�S�,��_,�3j(�4,+� ��f>��e��R��y�u�������i�|�,y�qtH��kgi4��8�Fp��d��>�@����HE ��
Q��E��mD^�j)���PC��Ě��|#���k� \�x�?5�J+���Zb����-��v�#U�c$YNX�ZZL���-�Pln��y�:?��c#qċ�3,�L�a;o���5�n�R�=1I���v���	M��6vi�=�Щ� q)��E5LF�?u3.s�P+dԋM(��a��S[�'.Ã� ��v&���E�`ŐV#�����Q���@~�_k~%/����va5�5�j`�D�T9�+Zhq5���HpO_�<e�>u��İګy��v�����J4��F��g�\E���d�V\U]0%#��E���D�ћ����ΐ��[DN:wv�Hnpb��\�6����.�y���|����_�D�q3��KJ��ҎM.�P��}]��� �==���l ����T %�g%��+��w�'J`���,�#o�F�O!/)�'3��C��>�Y�D�
�ٗ��^@��h6��J�hX� 0�@��W��}�E�����H&/hc�:��PN$��!���
7?P!���=l|5��8�;�v�'�e]%ɧ�p�i��G�++x��Y~V`��1@1~〆\��S��-9�/򕫈��@p��mL]�3��O�6<tA��gh�al�DI���{Kx��ЩwX�J������+����N�izU7�M+/CJگ�f߀�Mc��{��1��.�k��2�/��5���b�N�l0��RP����C�ق��z }�q,jԿ1�iD�z����43��;qPB�l�h�<rwWf�����4���%mM���w��L6��>�������v4d�Ǉ:�Pq�f ���cҍ�=�g����o��{N�o2�V�X�<V,���s�6S+��l�̰�}}�����n_�g�E��{�׀ڪ1@�i~¦Δ���I0:,EșE�,���J|�̌DCV,Ӑ� ��v������p�Z��. 4<V'z��T��sk�c�gn\"˞��q ��e�ݗ؍
ĄH�nQ�B�2e�O+�t��ڲ��F.V�Aӕ>��H������eK�����'��B�F�L��F�DУ��Xh�\nL:÷�Qbo�,��Lڦe������pw�ӻ w��F�j�\5C�m~{M�]dvs�q�t(.⣺�O�t�`�3YfbL�7[�z�z(L�Ddq&����׉ V�b�E���x� ��`
���a��͋>3�\�kѻ��|��݉I���<j̱X���	=���,��7PBk�LIU�F��!� 9����Ԡ[��^��S��$'[���;<�nZGI>�"�u��m0�l�r�4�d`@�YMH:HҘ�o��	�%.>��"t�3wV��8�g�q
�����S�?��k��8���ޱ~�V]��k�� g�:�.�(�6`�������*��K��/p��b�����y
pTQ�t����^����"{���<y�%������j�͈��t5Dxغ�����)M#�r�`�RK��*��2�凡y3�lFu���a��._���q<�k��a�Or6VH�Q2��}�'׷�2l��y�пɔv���._T+[�4ct��ޯG/c�(�VEs�_�xz����� �z����!�`Ҷ��s��ɟ=�u@��#�`�vE޹�M�zsj��J��KU=^���S��N�i����_��Ӕ*/�F-h-�m/�Y&c_��k a�>a��f���>��l"����r���!I=81;3����lK??������j�i[m��8��@@�i
��8��q�R��6_��Ța��^��D�*ڎu�죠T8X�ͪ`ϲ�F�b���W�~�p,K=I���s��&?n�9Juk��YQNLr����B���k��
yP�<��Ecν��\��m؟ȳ-�ǻ˓Ӥ��b�L�u93��\P���'��ٵ`'m!�Gv�#CT_Ë>����!�H�0$��ɏ3�K]�3E�	Za���AZ�ܝ�:��W�w�˼�G�w����A=\}�J�cO���!�'p����cR[q?���Z}����~�]C�as5e�(p%,��w��h#���"z2�Ϥ�"�}��Ͷ�)�$�j��tԍ�!����r�Qħ�z��BF<�b�h��i	z[���g�[ؕ�Ƕ���`��%d��E��q}C���0�I��Dг>��/ϰ��5��R�P���*/����OI0��-��|/����-�ϞA�A�F�,WWn����_̜S�R�N�R����_ŕr�A7�b=S�kMHH���?F$�	{׷a�L���l�?�������qnY�e�!�{������Z�hޝ�U��P���G�}Śu��2πrM�Azt�4S� 4h�\��w��|�[q�F���	󫜨�@Ì=����Л�ӗR�)�S ��݋�3�x��R5;$��u�kI:�Gesf�r�(0O9�(.$A��o��7֫)媇G��L�m�@}�v�|s��ǖI�`��:@D���{�|�Blhf��zX���y�XE.E��&�)g��d�������܉	8D�q<)\((Σ�ɴ�ȫs�*z���dGk��GT���菲��9�2�'��{5'RTC�QCǉ����e#�o�?5�tJ2F��,Dǵ��vʣ��-9o�[R�%�c⠳/E8n�/�U����e7��'� �4m33�/�� ��2&�o��y%�*�T�/"QY�R�.�G�f�V��	�F��VO2�2O��V�-Jb�0�I��G7�S&�G�?Iz��z�r%���J��]��Ļ>۳�����wVCǭ�ћ�C�n��rk�B�|�x���+5c�Bp�����z��´�Ĝ*�� $Q]:��Ts֫+m�ܮ���5�z</��<o�X�B�]N���h���{vXA0��,�l�#R�q% ���J�\4��*/<1:|tSz�ro(ϸ��p�UA�V�~���
���!W�sB0	wrU!�"��'؋������a����F��uBe�O�	3�ûM�A V@G{⻃9�<G݉���2L(5/tP�6��~�zl  �旃��@�_[��3m�Xݴ8m(ʖXea��l@���Ȭ�l�>��=@��QD�Y9!j�R���{�����P8տG��dS��j���h���g�.�`�Ͼs|2+Z����J�A�5�>?e��ZD�@m^���>%��J����};T}����/����R�^�a4i��A��wB��f�dN6�c����N���z�'���sTrg/��oD8qWc�˱E�;k��y���7��+C�=A��E��5q�!C����J�2I�[�+��,"������})�o�h1e �������/�)��+�4��})(X�]]���*�������=�5���x֊���$9g9��{�����
A����tɀ�bP�&��MIX4���p�0ܮ/(��1�q����#яUm5|i�X���A���j�ڠ/��G�mX���a2Ot$�cd.C/w%��G�����5o=�A� ��5�����0�O�n�N7��:"ʶ���� �&�fS+� j��E~��p;�B�ש�-�|{m�f%ir�άPTXv�k\z����^\G!i�-�Vu喜�H�4<�f\G)��wI�.�{��6��,K�4>��%9Q�l�y싲��"�ꃻDӿΙ���D!�o�I��d�.�Z,���mm9�&�����࿅t��}4-e��5�{X��+�����QͪX�,i���Gu���L��#�!� Ի*�u �54s�Ѝ����2�;Ru�%�_�Z��vzϐ5�����xۊ�ERǐ�S�|ngb )5����8�����\����X�b+�� ���Ǭ��Ny������x�]�6,� �W(�	
?�cq�����G�'��(-�P^ԟH�װ􋴱�z1J��YK҅x�%o��I�t�$����=	#�O5dZ�YK���OH��F�h�k�˱��7�(�������� ;x���QX��-��a�Vl�,�$��!Tx��K���na	o}3Z��0;ڌ��o�aR��i�uV��l��J38�����wH��6�[��6Y`�	�
U�&�����(;��O��l	�ptY��p�na�4X��~�"��J�G�<V �e$R&\^�}^6�čU4���tQ�.eL���0 ��l��C�t�a�c�$�v���أS6A}Ń,�2k̑�(�L.���<����������Y�9���'��Q_���9�h��$�	�Aw7��<����FXZ��?7T�J��S�;���<��1�\/Y$އ��拉�3a<�y^,&�+4�1���c�\��1\M^�ߖ(Yto�FH�������c���#�I|1|��S�=�.I�����۪X�Vo�H�U<��9��H�	����+����i�@������Zm�G��W�W�2C��;5��H~t]����h���2��{n]�D~�_d#o��ȵ��Y���:��L�QM$�����3�D��T��4 ���,gU��0'�,"�_d��'��)�B�:����;?L��]��?�Z�;� ���V7%����}p�OC��?��g/�ul�@M�0}R?{��T�Pj�Ip�+��v� �Vi|�֨*N����a-���g&Ȏ��	n������D�J����[n�yAhh9�H/�Y��7��#��\s����r;��S�l�����g
4����X��{���Z�_ol��"T���]�����#�]L����>����D�{���v�?��*{l�ڕ��>��C����D�c��0��[�0��i��P���w�����b}a"�����Uw^y!�Pg/��TR����Q@�	������W+rđ��Be�z�Ұ�����7�=[Q�6�$B�|R�����M��D�(/��7�e���d�8xro�ʐ�&Վ����(EgC�Z�̞%bM?l����dO��`bd��w���?⯧�:��ˤ^���j+�|<��5S&G*4�6-�j�8 j�D���8���K5Fj�z�hⱋqP]�l9��\!q��6=��4����d��|��Y���9�)<�d]��P.��b	3�=o�	��ZS@���),�=� �� 	���rН`�rL(�q��qëp��_j�0[^�i��bm�H��od�*E0�/�Υ�+��1?.�T|b�0٨�L�׃WMsN	E$��,�ÿ5�ӏ@6P����=)�-�@`V��%��?]�t4Y'�Ft-JI4_4����M��\)�0�#��X���*�'֎Ֆ�κ�b�h:�z&:�G��nI�M�2��>�M�J>A���U��~JQޤAV�v���3�W�S���зW*zM����
7i�#��5�lD�j�?���Ӟ��e�E�,��b�W����v�`N�ۂ�%��F�?�t����K'��)���x؍L�,�ƶ��6uxD�ٚU;-j؝�XS��b߫w��z��}o��@ҁ���E�����ρW�B%gn�?���*q���w���p���,ِ�wȿ7.���4����#��a�8:�z�z��^����)"���H��Ft.4K�cpu�\��-T��
sb3��9Z�7Yx����"�������)D����u֋��[dXe�L���䋄�/ǆ�Ty��dJ4	�2���'���b`�W3P��z�x�s�/ٳ%���.n9D5,�ɛ5Ȟ#OH��Og=O|�li,Ap�y��%ɣz�\?9�vT"G�''<�ԷٔR���/�wg��4�4V85���c��V���{^�7�]"R��c��)�r� =®��㟻�$�15֤I������Y��_{NZ �H�ͅ��r"����d2�������]�O����&IՏ�f�TJ�L$��*��GF��,�ߞAɓ���`Z��U����A���k���2��P|H�%=�b2Ѷ#��A�̽L\��rq������� �/"�;&�ʿ	�_F��j��kSq;w��"ZN�ӌ�Α��N������H�7�؅2������_"(?��(����rT�����՟�ޮ�_zD��+��f�{���3�n�y���;�5_5���P=��#�H�s{Ep=�%7�z��~*��F$LDz�]�I����1��ǔ��TH$equ��\O�N7�\�jf#%+�&wⴁ���CL,�]Z��u�zrYD��5��"��4H�a����W |� \���xT1(�;�r'pCof�L� ��Ta�+�e���f ��&~,9w�B�#f!wHv;��հ�e.�?%-lq,U�������7���"X�,�F�>�Mqָ7m��=zx�p��!xEr@6��Ӻ��p$� E���#3��9y��KW̿	���nc��9��2w,&A�����vh�i���Ʌ.9�N?���;>]�4�Ac�2~G�w�6r)��K��C�hE�M�	ǔd���G�C��vX��5�J]�k髢#TK�༦6�6R��j����� S�y�󗿐��%�אJ�v,ٽ ����'B;�����e�u�,g"��E91��R]�����C?��baf4���ʚ׈m& �B	��*6���Jy�6 Q�K�W��d/��7�J�8����� A֑Eɻ���d��8_��$��zoM��0N���\=�㌓ ]ᔷ4��n�L^�Au����IE6ˬ�8�A� B��b���+��R;���p��l\e�sG���w\�#��-�&2�E]�AE V�g����y�%��F�`H�� 9��,	z8����txy�$����Kղ�+X��"].mPT)O\��*���Lp�����/4h�n`'�d@���s�0��F�͜�N���V(��H��q!m�'�r;�O�řU/@V�L�xJ��s������7st�1�JΡbs�/aJx;ܡD���,4�.{UP��K�\b0_�]�$�����V���i&-��,�����������1P��9N��H�7����m����؋ϗ<�9���-a�6s�:7�i!P�5p���"� c�`�^Ӽ�±���0���5�_p�f�W���\�D1k��T[�f/:�P0��
�g�=��=1�0�ǌ<ﲋ!�&HY��(��&�w�RuvL��(�늯��#�a�'����\�8l�E�5S?�e@�V�y��39���9�Fk0�0�e����t"�k��t�k:�4%�m�Įk�m����h��z{M�*&��b�͸L�o��53� �0nŴ��!���Ȓ*i;P�K�u���_U:�����0j�hI)i��b���.�:ڣ#�W�q�L��$_.Sg&��=�ZZ�e���W��P�l�>ds��V:�v�7MLk����Cu��DQ�����Oޅ�b�Hrw^���#��o+up����mB.�� ��H�︴2Wl�������kd�ZȤ�t(�Ԭ;�1z���f>�u���A|�#粙���)=�=F�N{��ؗ)�@��v%TҎb|��	r,���7�دȎ���V�Y��w8��D>m�����nn�O�����cF�uF��-0�C?�M���.�qhg�n��J�z��~�	�S�g6&E�YVi�.J�c��x�O�8z��ł+j�b����s%��![�����l'C`7ޗ{��,J�����8��%���&�����|� iah���z�er軎���E�˫�r�	����=G��oF����+cbN�]]=p�ظĩτ��G�Oͽ�WaA��zXM	�������Oq�5��[���~�q�g��j��i'�;l+v&Qo�{Ü�ܜ.���|6���o��U��;��4�RA�G^pZ�G'���Y(j÷� �i�V����	��c�B������!"�8�\ݒ���"�}����R5<k���j��m�ǃ���Ie��� ���c��z2�bĉ�M��J����B'�:A��I��G�N-к3������$�M�����
g4�l]�v��۱ӄ���`�|�R-	]���y5��o��!=�[W���s��g*n9�r���]8������V^bQ�b�C�M6q�"g@\�>��ߥ�K��:A��/�g�̓�4�����16���G@��7�ר�/�?2�ԝ�FF��ۓ���m��j�"�˔�X{%�gغqb6��l�P�����e x@H�}��hf�t��p�ZS�k?�'Eh�p�u~(�m<�
����1i�o�up�SHs�V�ϖ�f��l"�J&Լ{^9�sٹ�RHn&�Ѷ6�|b�,�k�y���.��s�HF�>1�^
^�fh����|(�3�ޑ�x�@��
)RZJS>�d�Fۧ^����K�͓��A�cKp�CZ�%S�����ۚ���U�v�b�do��?�������t�����c��_ko~j.�t�U
F�*��3�`�&ڮ���AK�.<Hl�����<�4���Ǳ��uZZJ�ˍ	�W�~���Z�#�`��[�ŶJ��s��YG��ǜ����leA}�v����Γh٭���{gG�z�&�s�B W�󺖾�Yxq6�s�3.�6֛��~dL��?�"�Z>���?�܆=�>Wʘ��=�۽ZA����l����K��ES��!MH����xj�>�Mi	��ָ*�e�BEM��'�8�[��s9���zw� ����^�,��[��7i��햬-��N)��(lmͩ
G��B|�\U]� ��^C�����=vY,��q+��N39��j�w��SH�]��������q��G�c`k���S	6�6���('����"�u#U����R���r���(�t�}ԧ����`��Ƿ�y �g��V\��P����0��]u��9C����:�!IS�DE�<!�,�q��\|1���	�����M����C{��$�����Ppy"�� ~�?4\"N�6���$�d�j�HZ�"z���V�2��C
�Yӛ������PD���-x�*yA���i��l�]
�dߔ=�hpYb`��i�(,>���"��;^h���Ұ��ֵD���Ӷ����n�Sr�����e(��PF��g����^��tH��"���V�~>��{�`�B�<�@���QP!�G>�o�_W�e�P�����ʥ~���Pգo�i�\�������d�:%��M�$�0QoI|ʽ��4a�cs�tT�M�]�θ �_�������X5�&&d�YH-�Ī���I��mm`\��Lo��2�������.Ǻ���6�ۑch8�,	5����o� ЈJ�=�ʇo�f���Ξe�H��*��$H�ԕ3n�<���='��jTK���fb�Ӥ� ��L�5N^�Ae1G�C��Z���eՁ=g�����Wo���-#k���� ��<�Ɠ���_�> v��NQm3%Y���9�z=+��6n���kqZ���5u^*��'f�y��ϐ�~b�g�/���O��9�7��~( ĽM#��R�ծ�-�|�8��l+xX�F�K�ʒw��F���J��H=�C5�T�J��ԉj
ٳ@�~؅�;�AS m?����W��8�܄�%^]ꓗ����]���#*|r[�Ƈ��Q?��u�	���<�"�B�K�c�>�m�bb=�ޤ�LY*n�^��(��D�2�LH�kI���گ�ET�:��9��;! ��	A`�B�A������&m�a����Տܳ������QT;�%
�*#<�q�y�d:|Z�t���YSh_} ���03���ܸ�A�N��V�y�~�O2$u�Z Hذ���#O*;!V�r�J0����TP�
�Qx2򟍯W�Ji8}!l>dMA�*XG��pGA�
�����Մ1����)�5���B	�ǟL���.PhW�#������W FE�s-O��/�����y�Ҍ�h��ɭx��s���'����QQ�{���{ꡃv%Q��cf�k;�ꈹ쒔�<�(���().�-zlr��.�-��N��I��,N�hA�q���^V�[�]�N!	*���s��#F�Ԑ�<���_ǅ�D�1-�="�eF���L$�[������6LE�gC��2��#_u�'5Oe�3�Y{̌/�#�t��#��wd�LlN���lz.m�}Ѳf����|G&jL[�����@��oq��ȯ`߻�4/�[�m}^�|bf��@�prz���OG��F��2��q�4j��W�w�Û/�0g��G8�Ԯ&�t
ޓv���Ԛ���l���Nh���P�ϒ>����d�5&�7M�(��� EX���K��7ؤ���Y�w^���t�"@3���3�?����҂��ׄ�z\hS�(~����ʺ=�a�gY,�,�\i�b�쎨g����=�G�-�Qz ��_���\����C7Ǻ��L�w������
[�a���㣶j�+I����񋴘�)��zGF���c[1�E¯I��/b9?�'p2JQg�E~h !4��2���K�UG�Ȑ#;)�}C�H��vlN>t2h.���S�9n���3"f�� - �J�5��b���q.%���b�q�P:���$���4OB��կ?�G��a���\��C>�(_��$E��n�vz{�����Ep�I��-TT�@�?�
�ŰYU!ٗ" �@2Rl_ߟ��W��8ã����$���-��wR�����K��l�!��J��I��u|/VrN&�]>YF�0c��,�@F��I��0:.ܺ���z�\)�jt\/�������W]W����w/l���"F|J}k@&g�f���'s������c̪��� Lm�,���h��dW#%W��{A���®���V�$щ0(��Sw�'�������M�U�zv�'[k^]p:N�u���x��i�{mZ�t�^�D��w��ib܋X{��Teb��|K)�^,����m�0�;��u����4�|�
��[���e��E��R]�h�d=C�7ՍP ��3c fHZ'��GL��Fa��Tg��dv�U�%�M����
�����XY� 'YB��`YG�0Ю��:K�:��^ƞ��3���KO�S��g�u��mhy/0���٥�����<�6q�/��y��)ԛ�*[�d.��Z�����>5:�5X{���n�j:���P�eE�Ώs��Rï��4�`B���|Z��A�,ԥN�74-��j��?���6� �Z}Q(l�sjs�g�8t��@D���E�݃���V��}�j|�������'��c��(�Bi�ݪ����+��\>[���?�"����po�)�Rh����Ʀj]%Y�C@{���t��K��७� ������ȡY�6�/G��	�ߢ�9�'��=E+Ⱦ�Dc"��>���B~LA�/Ԁ{ռ|@���e
1Ҧ�������	��&�$i��sFR�@�_�~�3#���b� |� g�M��_���ԉ^nj��Ah��`���_∁с�?ɽ<&|y�����"��NhK���M��UY��Lw9cz� �i���a�4�Ez0̑�ʢ��	M�7c&F~��$6ƅ����[����*�>�FƶE`4��[@��y����<�&חO���g�K�[AZo�>��H��|pl�B<|�e� �	�1 A�d��͞���9�R�5K�s*��^�`�b��2Ș�j������aK/`���8�<Ew�B_�\EOo�+�s��%}�4��:S3���ͯiL�+a�+ ǐ��#͋!�|Yg��_(��c��<2�+����H0���aĴ�{����i?�"_e2�3�1v�&�@{�u/F�%Nµ���ZL;�(��-K���%�j���~ �(әu���5�t �#Z��c���̰��׏2@��e���N�7�n��W��JfV���:�L�a��3�R<�n���^��c��2:�	Y8(� ����l+1匛�
�%�PE3���a]ө�j��Y�����n����N�b�u�de����N�E�xѳ10ˇ����.�[N�[�*5.=~vlN��"�%�,�������\9�_\:�A�	�c��.0��;�\���������(�V�U#w��ΐI�Y]�vvC�_�mT�64��f��J�K�Uc	(�x�1d�[�7�W��W��V '&{7�GǱ��1*m��}K��to ˗��@M=TVG✿¡�Jja�GrUz���,9!�h=|�w|�Z��-<�dѧ��/�IX�w�fB�q%���G�4CK�,䚂���� ���L��g� �+Ï�eD��	'��D�6:W]#u�֨T��G�6bi{�_=���4���Ut�:�y�F�����\%}�l( ���7|���,����.g��^I��Aa\�ב�#��Q}��.�+o�E\q��,m�N�b����dP!�ͤ;���'.&^� r��T���Bv���0K��௒W=�)�ۀ�h��"��'ЧyW�\�r�W6�5`���s�Ei�xl2g�@Н������c�;UG��ދkd����Q*��ꖈ{�����Dd�}:����_L��#mO����b�#!�
��n�x��.�]T{Ms>�(Ϫг�l�?ʐ��Z���>ql.�w�Λ�(:0�,\y��9t�ȥ��C�;�\u"V��.������"��J�&/�[�G6;\>�_��JL��G����M%��.bC��~Ս�a���H�^�<�r%��������s��D#!��ȡln�jT�ȥ�>���:X����`J��l��f��U����9��'"§s�����n�̽������9��L#~F#�Ц�2܅ݫR�^����qmK�Q�Ɵ�܈��4a�z f�DU�6�ۢ�k݄L�i�h^[u�7���5���mDR�+z��Ho���+��K���-��yb�ޥuvV�XyV��sb��pn���K��1�"Ӥ�B�n,sgH i�K�Zp)���kIhe��:�M��x��籨�Y2óL�s���;K3�ũ�^fT2�_����h�U<�����2���Sd8V�eԼ��Qe�j�Ж�ܜ+�fօЗ2���z�4Ё�䱠���x�WO܅����ry�>��o�oE
�b6��4�Lqh��#\U C�=!�X ��$�;�ĺ�½@��`��e6˂���y���I3ե %�c�ғ��u�2�A���㶁�뢃�5/���B)\��B�x�z�:�ĘF�����Ƞ��+��p�	sZ0��Ow?l���M�,��QEp���<��֥��'�lop.د��.G��7q�*L�F(_FBe|��{%���P}NE8��+�^wC�$������}����n������f�x�ۃ?�4��|B+�����E�7@?���M`R"�tæ��2��\����q_��16���\����w ��6>��X4�c7V��{ꗗDr�( ���jʉ�A�m]�<[�<r�=:����� [� �c9_�ʺ�4}֜�� ��f��:�k+dY��b r)���D4�<d!��XX�v����5��2z %�;�����󐝖��6�opߪT�^�~��&�P!�7J�=�m_�N3I6���A�އ:eͽ��Ρ:Z��$b��jd_�%�-�7���sm1 �b�Bޏ]�Kn��}��޻��u�ԣ��Zq��w�i�(�֫N�U$�ĉ��d Who���=�MC̱�ѐ��p����v�b8����o��<��X[p�@�/ђ�=2^tϘa�[�"7%(���k��H����Q���M:�FV��)����_��F���s�h2O�N!/�w2|z^H6A�����V���R��s�����jǑ��� � �Ë�� ǩb>�@�A�Ax����'��.
��̾.;o�˵�ỳ�8Y�i��C"^�q-��L�D�j�W����&`���W��l7��,�/:���ð��(�؜�+J�`o[H�1q��T�F�,�6	����g2�O�ݣ��lm�*�~NP�:���X��J���iO%��+�pb�q.o�1^��4���V\�6�è��E�{�����S�/"i���T	W�)d`8!�ѝ$UY�؝����a35=��s/�3�� u88d��h$�P�6z�w�n �%Oa����v���$�y�{a�d3�y#-!�6��1��E��*>������Cv��X��hFeaEYս��W߀p&	��B�/S։h�.9L̕�cf�_��?��� =�]�Fh�����a_(Wr	�k��;��R�	�n�:ʃ�J��u}y�˅���S�nU�/��@4�բ.�V����N�����4l��j;��ZO��J��pw�f�PK�<�ӎ��Ɋ7��Y���r�mBE�b��BQw_d�Y6qŅ�E�R<��B�R��J���R�S�7e�/��`�+��qzw�}K���U�!5QjI�p��X����=fZ�/��\�粼��U�)���r��^�ݻ�ևhI��p�c��m]�함Ρ%�1�	�]�N/wV�Hw
X��R+T4	G�*�����<���s��	�{S&Cv��=g�L1�w�?�V}=��@T�˞?	z��R�|��.��
f#e���M,��h�L�r�B-��X�����	��������1c��^0�iXqT����l	,��q���$�zU�m�v�2�/��_m �zܡ�`(�M xO��qM^����6|7Oj�]E���bZ�Eg[3���AK����A`�r���'&�#�=B���&�m���@�nî��e�����,��P�$Iǖ�ew�E���/��麽��3!��`�dq��e������T���J`��A^�����Q���\�"��e݌�"D�
�1��8y^�����,�g(��WԆouW8�f@�g��W<����"B�as��5j��t���9�>��݉���.�מ���BN�� �6�^��&˭Z�=��dN��ʢw�	P{����.��[�=����ol�o��ؑ�됯r]�J�\� ���2|�����~��@�h�9�)��3�hhi�L���Uaԟ�0�O����Kv�s��g�+�°�>�?B��w��8O�?ֳI�� �ͻB[Q󃶊k�Ȟ�_���R���`=$oƽ��y�q<�+*;���ejCy���6�R�ގ�*b��.!�}_����R�+Ct���#�����7p5�?p� ���R��8=��I!I5��[����E�)�HWE���˷�oi�w��A���Z�����w/%�1��x�2�S�9��W
z�m9I�R��~�ʺ�Y�K��]g��zy�Ƒ��M�f8��a;Vc$���z�Û
�_S� !(�ÿv�{֌�Aę�Yf��=����dtoҊHA��F�>��_q��R2�y.��u��)��X.y��Ewx� ������wG8�����ç1k����(�K1�H���TcLLY���Kc��/��c]��&��H��{��?E���kR�>پo��C�i�� ��j���ٳ�_ʜ�j��S���2��D�4;�?`_Z�c!ɲ���x���:H؉�$O-��n¸��/���4~C�F��� �h�U�a2�y����ИaP*�x�b�e9Nߊd��b,����<{
]�R	����j�����M��C�ڜ�b�5��j��<�]{p�B��/��
�(ܦ�R2�d��L��b��];q���G��|*r\V������ݼ(Z<����Z����AMn���%��qݔ�;��[Ц��d]�rKnU��L�A^}�k�ph��<�$}�W�!���	bۋ�f�)��9��� �@RTi�ə,hIZ?]�<���p�!r�W�6� u^|�`��_l���fS���I�0��]Rx�l�h2�p�������΀��X�CQ�ϽHşw&�Y�Y�t�����r�Fe��C�{N�����"��'z�#M����>Ֆ�F��2C%��2��:�KA�0/��S?����*���j&'�E�, Е�c}6[&�7�3[g$E����
Vy��i�ð��N��-/�KM�f�k�|sMWN����^�L����s�x�kn �t�$n����	W0 �S�k�)�ࢂ�(��'���5��K��ڴ�F�9Ae��n�`��`K�A�h�
8c�1����P���)�`�'��)�#��w�w|�i�ċ;�^�w���U�V�<�	_��y�q�z�{�nƚ�x,<���J��X�c��	쳖i92J-���*�J�͑]�j���hp��_<b_j<���r15zZz�a�73ň��%*	q�������5X�B��\lK�?��p^�_�逛-�_6HEx)��n�W��P�+L���`Ws�r��̿5a#�|�p?^Jy��s�=M�86YRc����)��!��TzJ�q��
`db�!Ҭv�%h;�}�(L���F��%���A6�n�+�S�q��N��~����uD+]��� �x�rbl�^��®� cU�ج؜S(�r��gI< �߀De����゜�&��'  0;yLMN��T��}}-�Ш�k�"d{d�dI�����f������ͷ�cu�uCw�l���qΰ������XJ���H�{�$�[��C1[�nG9߬����#(|35�0�ʹ�T3�HvE��x`9;��*�D���@�'�m�kv��覛.C?��u)��ڮ�vqA��i5�,�mw�����'�� ���o�b�*~r�$F��z٨��1<�R�*/�cz|��pP��p��,�쩘��Tc
4z���ԸR���rk�a� f�����=�^����r.��̧�᚟�~�P�_w�&�ē�Ѥ���'���yt_��͓$
���z AaD<T(]k=V�C���$k���m[�}*�P��N����t����d��_�@�S���o}��//n� � �sq>$�6�2�jJІ�b�����=t�'�K`��0��B\�ha�!*��UU����K���)���:�ә���tgPʖ#���Է�^'�yJ�(YX�T�[pfn.a18Y��Tk�Q��^���^~�3ml[����F����߿#|���X��/)�Q"�WkB�:M!�*�*����N��Ԑ
�ң�^�u��s����I����u�}��L��w�%�7o�E#"-���^2
��BD��O°���3��������Ȓc�����U��C������r���=�J�l�
A��q��Om`��3¨h���(���hcr�>Z�˂��ۃT\UT  �ا�I�)[�Ku�Z��~�Ê�����!����T�r��#o��%�	2D�t'����gl�J��!�����>�	��.��~AZ������'�QB)�n�UneJ�L}e)�[/� Ȱ�Vy"Ou9p�Y��JPY�K���P��r^���@����<T���^�u�Q�h�pb�@�Oʃ����ϱc6$p�v� �X��^٠
�S���~�[����r��W!����쉱Ճ�bڝ��v�R:#�qR�H�ow�6�ը�7b&�} C�l����r�%P���Օ�� ��g&/��5�~E�܊`�FȊ�]�-x)n�P)HA�B�Kv4*�1թ��ȳzʻ���{Fz�V������`M �R�}��s|���o/��ٱg�,W�*A�d���FY7jL��gk���I�zê�u"�n� 5��M��J���{1����O�y'�J�B6�c�%�6R�v�x��;9Y?5�z�����_S*������'o�ɲ�����r���/��9;��n�gдP��c�3�D^��a����AY�#�Y�t]��c �n#�lGc X!ؤ���ܑ���Y̛��6�3o��<k��փ��(by�RT`L��0#ԁl�w���}�L�7��%���{������Z�T\#8Q��P? ��6?h.�)��O���X����������^'����:;ys����G 7���s�b)XF��<'���B*eU�}K�_��pY�^�'y�0�2���@���}�?9��?��� uc�+D4p�Ŷ��	Sa8�vF�B�Az�7�|U��,�IL&�d� �c��cew�
q��[��@l��E���Zk��Ni>�����$�UPŸqJ�Q���Z�S�jU����Y�N�'��i�/���v�|P-&�Wn̕`@&��h!l��9��%7Iw����_ökk�Olh��3���
�6$��Ί��$�ŲQ]@�q\�B���< �H�/q�W���6$55�Oz��v�`X[���r���,�5[����G��������#m2�����C�bx���C��H��8�V��)��"l�Q�L��r�׵m������me��Uک/O(h�
�B��5��5&T�����`
Y�!�(��ƽ�J��o^��c W8�u�v�2���kD��8���Ն�m���R�}�6�g}�+S`!z��CHg^ڲ�y��N�]!Iz��1�����Q�x�0�d�*ް��H��}��6����k_�����AC����Z�L��'��i�7H>v�ᆣg-j-�$4�}�U��ّ�lV�֙�p{㪢� ���$�;�%P�k��T�0��bN�'��fm~�$^�
n�#f�2�i5�����)�R��T	%1�"1L�2X����z)��S��*o�N�ZWF~��6��c��eIJ�}�f@����Ѹ��%pK�=����_����C��5�t�7�pi:2�4;�Ă��&�Gѝc�N�{;�FU��:L�S> ^ZB��Jof��˫�h�W�%�;�����}�
��������;Ӑ����v4ηHJ�(N����@o��n�'<����d��X/��@�	�+o��d����X �a�x3]���_���.hBq̍�,G�J��q$�3�G��\��e�i����=� ���cߖ2�QE�Μ +��q����\�S��M�Z�3:n���M��+Y����Y"�C�t�!7�ie%x��� �#;ǙB��.|ڇ���c ]wNT���[�;FS�T{��.�E���Z�|2/wF�T�N��TS�Vs!�-�2V��$"B-u��?��lA�c�{��N���D���C�]��uM�N��HHL짠q�1��J���F/l��5X^emM���ᔼy�^8��e�-w]�'�Z^w�JӇy���@3f�+A��)��S����pf��?��)s�k�=2Sc {�岁��92f��x��/��s��O�.�l�6�	w�ڙ;-�`b��qͭJ#��1�Q"=��Xi��z_3�}�M��z���A��	ͯk��x�5ԙ@�t��+	VP��D�\�P��J/���X�ك?���Q����$'#Ix�ݽ��x�����@-���۠eWd�Vx%9'+0*�hd H��e��5��ps���Iaq	i�52j'�!мI�=��7��e����e�zP%{Q(4t_6�ћ>CO>x��I������ϕ�H���� 
��,OA�xn�`�����,y�-Y=k$��@����W�z{3�\��<�b&c�vY��j�),���D��#��+��'xZ�~7�"�32�"�)�x[{�3 ��͌\��o�"^�l:�>��Z�N���f%��u��%�*Z�i�nJz�|(w��h0��1�8�L�
��s�C:83h�����Ҿ�݌ލv/��\���8=�E�	s�b��1��\2O��XM�ي�D]�[��"�O�a�o��~�*5��B�H�U`��D	�E����ߺ��	9�i�?�?æ��5�Q Q�u��s�I�j.C����\/�b��;"3�D�rd���]�k����H�i��u�d\G[�o�U��5roQ�r�`Y�\��uS�\�=~�(,ޮ�����G��Q9%����}#���߶g�ѐ	rDt#Jv]�È�+Ƭ[���w��F�g��.�v�<4����)�@.�5���x�ˇ�2.���m��u4��n>-2)��ƒ��%ɍ�v*8"��͢=9�Ҷ�A�������5D�痩��+��D&s�C�{�_�`��	�g�����IJ��*6�NRr��vI�)�h����e~�Cɯ���Jԃ��:��ۋ�D,,�"�)����d�����za��j̨F�U-|'�ە*���$F��V��d�BL�9Z����ӋabQ�-o�Z2'ĽJ���jau"LS7X�!�M٠Ɏt����g�8���;!��(�X�����<@��z���U�\7����m�#)/�r��hV�	b޶��LZ_թA�C"��F��hM�3��b��a��cJD�3o�_�]G��]�G)/z5|*�i���9�nů����M���/����S��y��`�n%r�J��%������M�ާP�u����u��xy �i�+^�)�U􀻴G#�DTy;R� �VH��7�=�����y�e/Bňq҆ �J���:��G�d��	�?��0��8�e(���r��7��ӟ?޻޸�:1���}^G���/�!�[Lް�$�Ѕ���N�A�v�v+�r��c\Id.�e�,&���C_v�)N}��{j�A,-�Ч�x#��&�	��Fe%FdL���Ȧ��jq�@RL�˅��{�A�b-z`��%#��\fI'dS�R/n����?� ,����P�F�*`��ׅIdd���w��^���s���V�qA��w�%wW�Z�=;/6�4aC���W���B�����^�2��p�?=�ɹ/awb�H�E��I9��j�}�< =N�`jg�Z�a���{{���G胷�L(����ӥ�L!&��*�����p�����mN%h�2��G����]�P�ˇ���k������&
��ħYHNGjIz̿��u���3X��	H(R�������k�o�g:�z}��
w)W^��oB�G^���C��=��>���]�ob�6���cÄ�O��9"��'@_�3{Z�?T���{��	P�C5��A�:�r9������CQ7�ϥ�2��y�!`Vd�M��;���U����i�hFׁ��Pݧ�i���`��V���21������i㹵��{D42���W�Mh��m�������`�l�(����;�D�K�<S��?A�� ���:�p<�Y�3���V��(Mld��/?�^%����wwVR��7sd(4�����Z3礵��m[�SVL k*�x:���:����%w��^6�S����k�~��+_='�
y?׊R�D@o��k��9d�p����?����ƫ�*�_2��f��q�DJ����a��HR��\tj���XH���\U�03���%���q���#+ ����6z�$�̭xs��4=A�eI��D�+�cb�%_�w��kN^mvH
�p&�Y����̤ѐ�^d@iw@�<��'�a7I�jʕսH;�K��=�� �����AO$�xqo�$Sڌ���6�xr�Au!��K�4#a`o�j^:˕�� �_ЏĽ��R��p�T� ��ձ�*<������6M��V�֡i��I��B�G��h�4�S�[����D�#j;�؋�jOe
W�tB�qX�n+t�r�{î�B7��'c�R�^�=�3\�n��]� ��k��l��{�{R:��4&І\N�"�1�����Δ�4�"��c����K�Dh��μ�[H�|	U�ϸ^+62�/���>v��Y�@�{�� S�|�N�Per;vD�?���,��lC�̲�zm���J�	����������*�QCo�z$;�<�)�"��]W8�η�0f+�����5�o�v3ʽ�9:D�1�
D��_5�7�(gk�]���֠;�����+�r�W�I��v>�'��v ����O-�ˊ��wWZd��=l2a��׋�j�}�q)\ʋ� E�精��@!iV[%�}�_����:�7� 31��;k�U�
�Y@o�q�N ���O� ���Y��|z��D�?����}�Nʯ����u�ob�lηQ��N:*�7�4��ݲ�УW���U�f�=*�e�L���-��z�Z��/kS<��s?�>iX�BJ���^0�Uy𸀨�c�b�^6�X��5�[r������җ5��:%��A ��T�9���M��A�U��Њ��N��V�L9���^�w��e^nv�7����j4�s\�<���#>K�}���E���� �	7JCEU5�m�w��#{@ֆ"	I�xmBMN�KZݓml����N�ԋ��1*����,:!h�<X�ć?q\���gu.�"�w���%�X6>���*"iφ�0�}��L�.�]���0��Y���b=i���V�kSL���fq��.���j��=A3e�,|}��2�8�X����)��̂n&h�%���1�R������}~��^���V�)�3��:"Y-H_��}^R0)�l����$��M()�ra��WTqKs��]'v�i��5��>�,�>��|I]�������՚�����:�3�Vd��_a8���3s4qÜr�މ���r��>X�Ł�-:���AV�'�bg��B6��<҅�|������=åL�|����G�1:Vw����xOT�.��CY��Y���P1�M�����`
z�S��\�wu��!�m��s�Uej�u�
+��5�П��t�QOt�<a���%�	�s�Cx1�at����9hfL�g�N�J�x�X	E#�d�q��Vc�l8�_����Ē4z	�{��CV��*P�Po��H�H.��
:�-\@ W��[��2���%�T� ����3*r����-DmȘ���b-'��n�G��#4]#	�1_�N�_�F)��}�Ҳ�'r:St�z�t���*X���$�	�;��ulf6{�� ��'�j:�ז����Skl�����U���/��7cu�U��P:��l`h<�������P_N��a��NAX�E+���Xi�?%��G��C^^i0v�"��`��f҂hác:x�:�B�q�0m6�,OP�*��2Fժ�	"v½ӕ��L�>{o<6e� �D�[գ�������P2VC�.\v�H���%��k!�����#a��D��D�N"u<9��),l�`u��"y<Q0�D��y8خ�/��uϦ`�c�����p�$��L�t}W%��nՏ�4���㤝4l�Ӳp�8�'�J��������d*T�%�-qm�����e�\VZT�����4����B�xW�'���=l�C����+��97	���i����2��1��l\፜qRc+���'�q����X�E1��� 3��ʮ��2/AQ�3r�&tA�MF�o��c��.��z�4r��)HOk�Q,UY��3J�_726�g���c��">��P���I��GP�����7b���O���E��g����Y8b���������@.����Y+.�dJ'|�������su��A����;�kfV�����'(�Є�D[wgsm�Cq�Ö���[ ��,�+'���~��������9�{�ה���QFр]�WgC��M��L3�b���V��"].ε���>�boFɳ��~�
�#�EQXzX������wX����)��7Ÿm�dPd�f��W8m�֔�]��xX������L���>��J�7���MA�y/b�%�#J���+��� �j�T���a�^�#cȼm��:��ꬌ`/���HԸ��}sm�gd�"�ǿ`y������gl��/fVZf��S��B�(�X� Q5��N��ȥ(��0� L$����}@j��>�v��rXfR-r��#j~(��K����d@�:.������!�nl��h|Q �JZ7H���H�T*X`ט�a8��re�GK�����	6��R��_���o��L���	b�!� ��9^-R�9�h���Nx��-����B�4��a%���2@�0����iS�i��^��,%!��нZ)����W��Qni��?pV�.��=0O���d�
��ԛT��
!N� ��`���Iڑ��(!��c��g=7ӓ6|�L�6]r���D��*;�M��cܝ�}Y]��Θ�$�Z@ec�^���`����U�}3o�.z�O�Ҿ�o���JWZ�۴�B��/�,T�
�ۛy�Q�f?������b�X�%>^���m�*�{�V��̴Ԩ��3f�}&fp0��:�����?N'�zm�ϋ�3 �L)��ql����l?��u�5�
��߾L͒�:�P�]Kձbq��}��*���E��uJ��tq��ғ�����Χ�x������ݏ��a�,V��P~�)�#hA���AwW'�u��IJ����He}��:���I���χ,g5vԀ�P��%�?����� ~� ;���f^tFo5=�iA�Ffv4su��Fr��� Fy[%�}Gă�3�
�^�r�q}�XǬ��1��Q��`������4�o��Jn��)��kj�7�"����V��hYr���.ӿv�(�5*��M,N�:my5i�Üp}T4�*� �p���\X�YU��x�ٱJ_K5vz�:Ť��@8���IN�8�����7��SpV����jKe���pW�ŷ�a�/����1�a=�C�{�;�͘Բ�/������҉����Y���go╂�T�#�@��)�k���B�kO\S��<��(�^�P�T�^��j�^"=��$;�҉�+g!5p6�,�QޙTh��ߤ����g�z�g�L{o�o�nL�j�"A�67I?�����������YvN#�����g)��x��m�'�\V'��c���̪�u�t��}T�� `oi�qP���'��c� S+�o�Lb��v��7 ׋�X���×B�����4d�ip�4K? 	������H�b"%��*��6g@R�nlȂ&%V�π+��q��������+�J�����Ĳ�	��@3�O�ZO���xN2��	6]�~&��i�<f:�=�<>������(~�+T���[��U��8����c���DT<j ���+���z8]߶�gZ���ם.@���r��`1a��W�oU�f������E^_>I��v+����,�K0���֦'-KUX�>~]3(�}[�
�F
�ܧ��N?�l�V��1I���y�w�@B���R��B{�݋��*�U3d��rUfɆ�Ҩ��w�'R�a�	g��Ÿ~�i��Q��<�ŭU��+���G�^R�(~��0��U���N��,�yz�,0�q�)!�ct!(&u��F�-P��g����o`�WX4����+��ͣ������k�#��.�e�7���;r�X헧��8 ���3��ͳ}Y/�DNfb9�%g��Q�a��?��u��.�"@�|���9������I[�U�z�ik�;:!}�;�F_2���2ZL`��?���G9�u�ʛ+����ՎI�`�i�o��ڠ���\����)**$�|��b��r�\/֚GE�	ر�mTi��M�LS���Q� �m�*�i�R�x'��˅ƾ�nvX�g���mMTTi�|�,7�2>	��V$0�Y-�-�@�l�g�1��7Λv�^�u�,	��S���m��X��X�� �/�&��]t��!TFU��	���B�l��b.���)�=%-xÞ_彀&Ç��uI��&v��SNԒ�F|U��d�?��]X�U�T�1/B֧�n~R��
-I_	�v�/p-���_Ya���wH�?�̶ b��V(~yf +HƗ�d� .Z��1����ʽ�Ɋ�����ε^��|���j'+yU���؎p���̒�� ��w��M�j8S��6�|"���x��e��$ɼoό�+�����72�������hL�^Aί~x}HKq�b�zg��bp$r	9:'�Ro	����'{4�<a7��z�7V�W�C���d� m�V��@a5�җ��gИc�����z�'b��})�J`�N�3x��3@DȰ�+$P Wmt_�P$/��jړG���	�t����=|��A��	,�#����Qjv�A_F)��L�&/;��\;�`�7o��p���_�	��WL�}y����"ωM�Q�����N>��$�A�	$���I��x�j���h���(yE����h��{u�
�B2��NM�8%'���]��9��8�=�^O���?@+�$<1ej�=3�l�p����4�2����j�ǩH����?̷.�~(m �u��y�H�Li�E��o%�=��g�H:�;r��i���6e1���N-�/�_|I��N��(d.�q�T�U�DĪc�>F��N�3a�
�<���2�6�4^gm+��Od/W׽��Ya���{���W8��ta|yK��.՝am�U6�,�����SL� T������G*
���>�mǳ!yP���G����� �j�w@����$�75D=?��z��<wu��򙄔�di��SH��.G�P��Vf7)���4+#m\wl���H��"�mZ}�Ua楘ӹ
D�1sO�+������m�]�����{5��-�H�^Nb��\m�<(n�w��yOⱼ�.%����J'�s�Pe�b�)2�I�UQeT���Q{\�#��=/�v��z���E���W�BF�#C�������]q3���[	D9�P��r�g:�ق��wP_E_s(:�<�6�Y���x���W�r�W��X5����fb􍬑o�W�k�N�ڿ�ImR�J�Q����B�}������^�h�datē�4Q3�t�X0l�FQ�7�,��BV�u�`�군�pD\ϩIg��F\ΎE>���e�7�gr�
�/n����qGT��=�Ȃ�YP�=���X/�f�밻NrI��D�o�!(Y�V")����'�k�D|��ࢧ���~b��#6Q�i�����	�}1]sc�%º%��n)����s��d��*IlW��8P��[�1�!�fQ"/F��1��<�[Q�$-������	��R��6�B,����M��[Z�P��7���qH���q�f���M'�B�Y�KM��D������'T��Z�F��J
��Lw��&z�:�i�YϕR��|�K�i�M���r£�9i���k����6B�XF�66h���F�ev9�_�������!#0*�ʒ����\��4�Tק��{���S�������
��Z�TsRXt��2�M��,�.�z�d�:<���_�<.;5�������>8���	`�4pԨ��)y{x��D:%!j�� �N+(穅P(D,W�!Q䓉��{fȑmc��_d�Y]�r�/Ժp�g�"��x
Ԃ���(�Z}�X5��\��:��0�ܐ���y���6x�k%oY�l����,3���v�g7�J��b��G��{]����5;y @�tI��O�i���0߹@^�D�=�!�J7R��{���:S�F'{���2���q�b�>�ڕ�$UY�}��'P�EҮ��]M�)=A����-�P��]W��^��V��|qhƍ�-5B`B4�w�tgj�S������<X�r�yt�����1�0�B�	�G`F4K�,�t:�fR�2��{�G�NF�k�:��g��Ĥ�����X�$��3������Q2��H�@�?t�;UK�CY�j����bo��0�u���n��l�h8������J�ߑ��/V$/�e~��2�M��{��r���i�!$ �t����D� ���9��>���yp���1��	�l���*Ե,T���t�)�q�$���p��H��ŀ�������3�m|�
�}�IS=��i�"�wspx��Q���yR[�C����7���Пv���7�-�@VP�T�P��h��sq`�	��ԡ"^�&�韰�G�͇w��]�b�
y��H���H{N��H��t��-��4�ˍIµ�3+���V��F`�X&����+e�f̗�]x�%z�	��k#���	r�nP�#�g���6�d¤���H�"{��o*��}�p�ZL!��YU!F}����U$�ժ?:ю�,�\�Mr ����*[ZVHM+9�[�N�l�G�`~J�1y�m���B�oi�����N�����̅�*O*��S�aK�<�;�B02��,��j�W����b��ԑ07�_D�$�rSЛ��zY��
��3st�U9���+H�VW�8�sӕ��gاV�-i{z'H���?�I�u	+DOz�5��B�18o�F�z�Jy�
N��n����,���rīe��~�}�l���5~�sX�Ƀ�]m�ՠ���2����h/�w�q��ލ!���QU�������0��~�����li�0�$�Cѯr�4�>�(<o��ב�}��}Ue��to
6�dH�`X���q��T�&�3�Ԯo�
ʔ^�Ӂ�&�Ȥ�����"�>˦t��u"=�䴰�hz��R���Q=�����S��#؂Sٜ�9g�HPo�e�EU��#b3bJ˝H��(�|�WZD�oU�L�<�1L6��|�Ϟ�y���?���>͹�)NH�tA�Fc�꠶O6�V�d�)Uh4:��O8����6�v��q���T��(�!�I��pzI�E¾�>.0�p���(�G�:��s�}Ȝg3�\G�N��v�L�[�[#eP7��c=�k�=�h_z��KtTX���m��@��W{G�$\JG�����F�2����*k�.х���D����+eL6�,M��2�x�w�2�*ǫ5�O*;;W��g�Gu0PR���c��$��&���T�v%��vsV܃��\���E�i�K!~$� �V(�JO�T�w\�����n.	�I9_������H/�]w�����j���q?*X�?kK߁�ˀ8Ɏ��v��ت����&���U��ǒ����z$�fY=�x-7�lA�T-��,؝7���
��l�/ VLM���uU�BĶ��G�e{9���rg���gb`!���p꥽�ٚ�a�:��J��`���5�)Bq�A!���yN�3���Y@7�uzӖ���oa�5~��>W�A�*�$m�N��w�����	EҤ妠?6}����#�{��
����~/�~�s����&~+71��P ߿βUU(�ʄ]g�ϗ�M`���R�(O&&`�@o��[L�6�p�p/э�;��p�\����u����ZRdX�����>���b	(sHS������r��	.�1y�B�^)�ȡ�f3��~���O��x�>��g/h�'A��8��5r`���ۦyl�|�].���d��T�we��4-\�0pӿr	{/?1=���_����Ҹ[�B�J��Q����/���K�(�4��b�v�j��M��	a�;%1��^2#���fu�c!n^WO�.���7W%_������� �H���A뇶�g��+��OyI��U.�ty�y��9�Q��3u�������ܶT�s3�^�� �Ψ��0آ��t.M��K�-|�㯐��a�/�?Ӌ�ߴ0���owz��;��C��*����12P70$�^����a�O�"Q�Lg3�g'X8���h�J~^�F��eD^��OVuW��Zؖ�;[���[v���c�i��W2ϸ��Y�{?< $6�\�mW�m��+���Cǟ����TI��hsN����[���$ ��?e�}��"��<�dZ��8I9̸�B.����H���/�<?I�������`��g.M�|.#��05AX���MP-$B�%�x�z��4ө ��c$9�|���T&o
�̍�"�ֹy��Л�����R~H��U0���TdI;�>�-��Y�<�_ڴ�8�¾��LNT�tG�e6ݟ�6�E�\����0�^3�O�M�� N����K��aOE��M����s�0��p��K.�W(/�,�Ӂ��!��;n�j�
�(~:�R��wJX�b� �,��0:3�8y����f�*ls~�4���ϰ`-�e[`�y�J��؎+���?+�_��OnǄ��frF���P6)19�t2 �h���0��4ij;V
���( ��5�ނ�NВwU_���:����*��CT��q0$�-������	i����R:O�G'��OGi�P'�z�����~��	��M1�[ 仕�K�-""�f\��D@�J��F78-yp���Ţ�J���Q�O�:x�4^��~+�L ԏ��A��!pq�G�����&���@�铩�U��U�db�����;���F��O�eobT�I�W���ْ�"��2$�Z�R5�����=��ݨ5��@XGbF�^�%���DF,\��U/J���GO�a?��/'6�u�)��y�X�x3z��Ć�r�EΡ��>c�m O��WY���j���,�X�WH��-Z��=am"�4AĞ�N4B��x���j�؆W��:���ȥ��:ѻ4�U&Υ��f�PY��	bu����l$�����.�~����fA?�������S��1�r�!S�6�}<����U�����R�E��+u7�Bi���D�0Z�X8Nx�����F���ˁ���F9��Aq�Boǚg�ݧe�@�9",��	����r~��Va�~�m�q(��9Tx�K��$�^j+O?g��3��CRxڛ��d��.F��x�dS�6��Y�P x�R2	��;'��e�����{�}��J�9�+���B@���c�o���x��_����SK�Ѭ��;���X츥�2q<P����D%������AϒwtYd*";�cqɊ�ߋ��R5�[��Bx�A����9�Pܔ��㞍R�n80���f�����R��b �C���D�!����I�Ƿo)�-���u�W�2�u���e.�e�\vb�����d����:V�˙b��تp���X��5"����g��H��oysL�v��s����s����p��n��;U�±Ւu��*��3�f�s;�P�����}�ӥ��k���j��h��E�EDj�l.+����/D4̶����p:��ώ��3䥀��OwZ�N/vu)e����E�'C�@g~�'��9+$�z��ϙ���j���������;�nZ�Tw0d̉�tCN]���C���e+��_ ��۪�\��I6mn��>@���p��h8%�&RҎS^��:Tg�aצ��L�A��u>QY��u��Y�X���X7.�cj�3��y�>��pϲu
�M����2(��8jVFb�<ꧽ�B��
X�y�g��F?��t&_X�dfY8�x�R�!A���������֐�Ց��D�F����^(�l8�I󲖥���4�Dq�M�8�J�����e�Pk��Hm����Juk��G<���-u�r����B�i�\T_�u���zxc�ܓz�&>�ʌ��@u�M�0�����v�aqd�o���AC1n�$�=v�����#l�]�+��Gf�zƤ��Oy���;�U�=�Uˋ���+�}�<�.�����(�
r}$���)���`(3썪�⥒">��/��^�_�����]��pIr����q}^��ei��KPʅ��tvm��a�Dȁ'��<^����RDY�v3��X9�ő�.��7�g��c:��`	��~��o�i��� ��B� 	^Ȕ9'� �K���o����-Wx�Ɉ\�@��̠�i']�nRD�0���-��R��@���A�8�
@�qc-dæ5���3�����0)M��`+lc�L�d�`��;��v��H^I�͏ۧ�M2w��1�F��.�&naz�̅β*�7��� J#�r�N 0? ff2��蒴�)g�8E���}Q�`9�'��F���M6���59��zu�8L�u�ѲG7kQTӑIҏ5��C�}>�c	���܏F�J%��Đ�U~f?��һ���a���$��<�L{�U�"�ԡB}P&�  �w[]�i_��894���z[wu)*��Fr����V8�<�g�G��C�,���n�����p�a�9�uY�^��#w�|D�G*���$ֹY,a	)��_dp�4�y}��'�re'f ��}^`ڎi�jV�!ӝa	�&tءbүl3�w��^�T��wV��-\Wa�ɼD �P6�0k�I+D(aQnX��ɹ]���Bc���:��D_Uу�4aw"�R��y0zf�ݺ\�2o&Q�x��W�n,�����t��6A
���U��t��DWV��X�"��Ԇ2ju�3��x(�,I�����&��T�5�π�uj�J<t��~$�^
���t߳Xʯg�RM��^�����C�ud�h�[@0��bҍ?K'���N�X͔l�*�o�[(*���"?�������`Z�?�g�	�X���-�@Yx�N���������k�ʆVC
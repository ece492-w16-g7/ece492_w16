// niosII_system.v

// Generated using ACDS version 12.1sp1 243 at 2016.02.08.14:55:45

`timescale 1 ps / 1 ps
module niosII_system (
		output wire        video_vga_controller_0_external_interface_CLK,   // video_vga_controller_0_external_interface.CLK
		output wire        video_vga_controller_0_external_interface_HS,    //                                          .HS
		output wire        video_vga_controller_0_external_interface_VS,    //                                          .VS
		output wire        video_vga_controller_0_external_interface_BLANK, //                                          .BLANK
		output wire        video_vga_controller_0_external_interface_SYNC,  //                                          .SYNC
		output wire [9:0]  video_vga_controller_0_external_interface_R,     //                                          .R
		output wire [9:0]  video_vga_controller_0_external_interface_G,     //                                          .G
		output wire [9:0]  video_vga_controller_0_external_interface_B,     //                                          .B
		inout  wire [15:0] sram_controller_external_interface_DQ,           //        sram_controller_external_interface.DQ
		output wire [19:0] sram_controller_external_interface_ADDR,         //                                          .ADDR
		output wire        sram_controller_external_interface_LB_N,         //                                          .LB_N
		output wire        sram_controller_external_interface_UB_N,         //                                          .UB_N
		output wire        sram_controller_external_interface_CE_N,         //                                          .CE_N
		output wire        sram_controller_external_interface_OE_N,         //                                          .OE_N
		output wire        sram_controller_external_interface_WE_N,         //                                          .WE_N
		input  wire        reset_reset_n,                                   //                                     reset.reset_n
		input  wire        clk_clk,                                         //                                       clk.clk
		input  wire        video_decoder_external_interface_TD_CLK27,       //          video_decoder_external_interface.TD_CLK27
		input  wire [7:0]  video_decoder_external_interface_TD_DATA,        //                                          .TD_DATA
		input  wire        video_decoder_external_interface_TD_HS,          //                                          .TD_HS
		input  wire        video_decoder_external_interface_TD_VS,          //                                          .TD_VS
		output wire        video_decoder_external_interface_TD_RESET,       //                                          .TD_RESET
		output wire        video_decoder_external_interface_overflow_flag,  //                                          .overflow_flag
		inout  wire        audio_video_config_external_interface_SDAT,      //     audio_video_config_external_interface.SDAT
		output wire        audio_video_config_external_interface_SCLK       //                                          .SCLK
	);

	wire          clock_signals_sys_clk_clk;                                                                                      // Clock_Signals:sys_clk -> [Audio_Video_Config:clk, Audio_Video_Config_avalon_av_config_slave_translator:clk, Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:clk, Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, CPU:clk, CPU_data_master_translator:clk, CPU_data_master_translator_avalon_universal_master_0_agent:clk, CPU_instruction_master_translator:clk, CPU_instruction_master_translator_avalon_universal_master_0_agent:clk, CPU_jtag_debug_module_translator:clk, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Chroma_Resampler:clk, DMA_to_Memory:clk, DMA_to_Memory_avalon_dma_control_slave_translator:clk, DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:clk, DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, DMA_to_Memory_avalon_dma_master_translator:clk, DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:clk, DMA_to_Stream:clk, DMA_to_Stream_avalon_dma_control_slave_translator:clk, DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:clk, DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, DMA_to_Stream_avalon_dma_master_translator:clk, DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:clk, Dual_Clock_FIFO:clk_stream_in, Onchip_Memory:clk, Onchip_Memory_s1_translator:clk, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:clk, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, RGB_Resampler_1:clk, SRAM_Controller:clk, SRAM_Controller_avalon_sram_slave_translator:clk, SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Scaler_0:clk, Scaler_1:clk, Video_Clipper:clk, Video_Decoder:clk, YCrCb_to_RGB_2_0:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, burst_adapter:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_005:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, irq_mapper:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller_001:clk, width_adapter:clk, width_adapter_001:clk]
	wire          clock_signals_vga_clk_clk;                                                                                      // Clock_Signals:VGA_CLK -> [Dual_Clock_FIFO:clk_stream_out, VGA_Controller:clk, rst_controller_002:clk]
	wire          dual_clock_fifo_avalon_dc_buffer_source_endofpacket;                                                            // Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	wire          dual_clock_fifo_avalon_dc_buffer_source_valid;                                                                  // Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	wire          dual_clock_fifo_avalon_dc_buffer_source_startofpacket;                                                          // Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	wire   [29:0] dual_clock_fifo_avalon_dc_buffer_source_data;                                                                   // Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	wire          dual_clock_fifo_avalon_dc_buffer_source_ready;                                                                  // VGA_Controller:ready -> Dual_Clock_FIFO:stream_out_ready
	wire          rgb_resampler_1_avalon_rgb_source_endofpacket;                                                                  // RGB_Resampler_1:stream_out_endofpacket -> Scaler_1:stream_in_endofpacket
	wire          rgb_resampler_1_avalon_rgb_source_valid;                                                                        // RGB_Resampler_1:stream_out_valid -> Scaler_1:stream_in_valid
	wire          rgb_resampler_1_avalon_rgb_source_startofpacket;                                                                // RGB_Resampler_1:stream_out_startofpacket -> Scaler_1:stream_in_startofpacket
	wire   [29:0] rgb_resampler_1_avalon_rgb_source_data;                                                                         // RGB_Resampler_1:stream_out_data -> Scaler_1:stream_in_data
	wire          rgb_resampler_1_avalon_rgb_source_ready;                                                                        // Scaler_1:stream_in_ready -> RGB_Resampler_1:stream_out_ready
	wire          scaler_1_avalon_scaler_source_endofpacket;                                                                      // Scaler_1:stream_out_endofpacket -> Dual_Clock_FIFO:stream_in_endofpacket
	wire          scaler_1_avalon_scaler_source_valid;                                                                            // Scaler_1:stream_out_valid -> Dual_Clock_FIFO:stream_in_valid
	wire          scaler_1_avalon_scaler_source_startofpacket;                                                                    // Scaler_1:stream_out_startofpacket -> Dual_Clock_FIFO:stream_in_startofpacket
	wire   [29:0] scaler_1_avalon_scaler_source_data;                                                                             // Scaler_1:stream_out_data -> Dual_Clock_FIFO:stream_in_data
	wire          scaler_1_avalon_scaler_source_ready;                                                                            // Dual_Clock_FIFO:stream_in_ready -> Scaler_1:stream_out_ready
	wire          video_decoder_avalon_decoder_source_endofpacket;                                                                // Video_Decoder:stream_out_endofpacket -> Video_Clipper:stream_in_endofpacket
	wire          video_decoder_avalon_decoder_source_valid;                                                                      // Video_Decoder:stream_out_valid -> Video_Clipper:stream_in_valid
	wire          video_decoder_avalon_decoder_source_startofpacket;                                                              // Video_Decoder:stream_out_startofpacket -> Video_Clipper:stream_in_startofpacket
	wire   [15:0] video_decoder_avalon_decoder_source_data;                                                                       // Video_Decoder:stream_out_data -> Video_Clipper:stream_in_data
	wire          video_decoder_avalon_decoder_source_ready;                                                                      // Video_Clipper:stream_in_ready -> Video_Decoder:stream_out_ready
	wire          video_clipper_avalon_clipper_source_endofpacket;                                                                // Video_Clipper:stream_out_endofpacket -> Scaler_0:stream_in_endofpacket
	wire          video_clipper_avalon_clipper_source_valid;                                                                      // Video_Clipper:stream_out_valid -> Scaler_0:stream_in_valid
	wire          video_clipper_avalon_clipper_source_startofpacket;                                                              // Video_Clipper:stream_out_startofpacket -> Scaler_0:stream_in_startofpacket
	wire   [15:0] video_clipper_avalon_clipper_source_data;                                                                       // Video_Clipper:stream_out_data -> Scaler_0:stream_in_data
	wire          video_clipper_avalon_clipper_source_ready;                                                                      // Scaler_0:stream_in_ready -> Video_Clipper:stream_out_ready
	wire          scaler_0_avalon_scaler_source_endofpacket;                                                                      // Scaler_0:stream_out_endofpacket -> Chroma_Resampler:stream_in_endofpacket
	wire          scaler_0_avalon_scaler_source_valid;                                                                            // Scaler_0:stream_out_valid -> Chroma_Resampler:stream_in_valid
	wire          scaler_0_avalon_scaler_source_startofpacket;                                                                    // Scaler_0:stream_out_startofpacket -> Chroma_Resampler:stream_in_startofpacket
	wire   [15:0] scaler_0_avalon_scaler_source_data;                                                                             // Scaler_0:stream_out_data -> Chroma_Resampler:stream_in_data
	wire          scaler_0_avalon_scaler_source_ready;                                                                            // Chroma_Resampler:stream_in_ready -> Scaler_0:stream_out_ready
	wire          ycrcb_to_rgb_2_0_avalon_streaming_source_endofpacket;                                                           // YCrCb_to_RGB_2_0:stream_out_endofpacket -> DMA_to_Memory:stream_endofpacket
	wire          ycrcb_to_rgb_2_0_avalon_streaming_source_valid;                                                                 // YCrCb_to_RGB_2_0:stream_out_valid -> DMA_to_Memory:stream_valid
	wire          ycrcb_to_rgb_2_0_avalon_streaming_source_startofpacket;                                                         // YCrCb_to_RGB_2_0:stream_out_startofpacket -> DMA_to_Memory:stream_startofpacket
	wire   [23:0] ycrcb_to_rgb_2_0_avalon_streaming_source_data;                                                                  // YCrCb_to_RGB_2_0:stream_out_data -> DMA_to_Memory:stream_data
	wire          ycrcb_to_rgb_2_0_avalon_streaming_source_ready;                                                                 // DMA_to_Memory:stream_ready -> YCrCb_to_RGB_2_0:stream_out_ready
	wire          dma_to_stream_avalon_pixel_source_endofpacket;                                                                  // DMA_to_Stream:stream_endofpacket -> RGB_Resampler_1:stream_in_endofpacket
	wire          dma_to_stream_avalon_pixel_source_valid;                                                                        // DMA_to_Stream:stream_valid -> RGB_Resampler_1:stream_in_valid
	wire          dma_to_stream_avalon_pixel_source_startofpacket;                                                                // DMA_to_Stream:stream_startofpacket -> RGB_Resampler_1:stream_in_startofpacket
	wire   [23:0] dma_to_stream_avalon_pixel_source_data;                                                                         // DMA_to_Stream:stream_data -> RGB_Resampler_1:stream_in_data
	wire          dma_to_stream_avalon_pixel_source_ready;                                                                        // RGB_Resampler_1:stream_in_ready -> DMA_to_Stream:stream_ready
	wire          chroma_resampler_avalon_chroma_source_endofpacket;                                                              // Chroma_Resampler:stream_out_endofpacket -> YCrCb_to_RGB_2_0:stream_in_endofpacket
	wire          chroma_resampler_avalon_chroma_source_valid;                                                                    // Chroma_Resampler:stream_out_valid -> YCrCb_to_RGB_2_0:stream_in_valid
	wire          chroma_resampler_avalon_chroma_source_startofpacket;                                                            // Chroma_Resampler:stream_out_startofpacket -> YCrCb_to_RGB_2_0:stream_in_startofpacket
	wire   [23:0] chroma_resampler_avalon_chroma_source_data;                                                                     // Chroma_Resampler:stream_out_data -> YCrCb_to_RGB_2_0:stream_in_data
	wire          chroma_resampler_avalon_chroma_source_ready;                                                                    // YCrCb_to_RGB_2_0:stream_in_ready -> Chroma_Resampler:stream_out_ready
	wire          cpu_instruction_master_waitrequest;                                                                             // CPU_instruction_master_translator:av_waitrequest -> CPU:i_waitrequest
	wire   [15:0] cpu_instruction_master_address;                                                                                 // CPU:i_address -> CPU_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                                    // CPU:i_read -> CPU_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                                // CPU_instruction_master_translator:av_readdata -> CPU:i_readdata
	wire          cpu_data_master_waitrequest;                                                                                    // CPU_data_master_translator:av_waitrequest -> CPU:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                                      // CPU:d_writedata -> CPU_data_master_translator:av_writedata
	wire   [15:0] cpu_data_master_address;                                                                                        // CPU:d_address -> CPU_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                                          // CPU:d_write -> CPU_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                                           // CPU:d_read -> CPU_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                                       // CPU_data_master_translator:av_readdata -> CPU:d_readdata
	wire          cpu_data_master_debugaccess;                                                                                    // CPU:jtag_debug_module_debugaccess_to_roms -> CPU_data_master_translator:av_debugaccess
	wire    [3:0] cpu_data_master_byteenable;                                                                                     // CPU:d_byteenable -> CPU_data_master_translator:av_byteenable
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                                 // CPU_jtag_debug_module_translator:av_writedata -> CPU:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                                   // CPU_jtag_debug_module_translator:av_address -> CPU:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                                // CPU_jtag_debug_module_translator:av_chipselect -> CPU:jtag_debug_module_select
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                     // CPU_jtag_debug_module_translator:av_write -> CPU:jtag_debug_module_write
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                                  // CPU:jtag_debug_module_readdata -> CPU_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                             // CPU_jtag_debug_module_translator:av_begintransfer -> CPU:jtag_debug_module_begintransfer
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                               // CPU_jtag_debug_module_translator:av_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                                // CPU_jtag_debug_module_translator:av_byteenable -> CPU:jtag_debug_module_byteenable
	wire   [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_writedata;                                                      // Onchip_Memory_s1_translator:av_writedata -> Onchip_Memory:writedata
	wire   [11:0] onchip_memory_s1_translator_avalon_anti_slave_0_address;                                                        // Onchip_Memory_s1_translator:av_address -> Onchip_Memory:address
	wire          onchip_memory_s1_translator_avalon_anti_slave_0_chipselect;                                                     // Onchip_Memory_s1_translator:av_chipselect -> Onchip_Memory:chipselect
	wire          onchip_memory_s1_translator_avalon_anti_slave_0_clken;                                                          // Onchip_Memory_s1_translator:av_clken -> Onchip_Memory:clken
	wire          onchip_memory_s1_translator_avalon_anti_slave_0_write;                                                          // Onchip_Memory_s1_translator:av_write -> Onchip_Memory:write
	wire   [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_readdata;                                                       // Onchip_Memory:readdata -> Onchip_Memory_s1_translator:av_readdata
	wire    [3:0] onchip_memory_s1_translator_avalon_anti_slave_0_byteenable;                                                     // Onchip_Memory_s1_translator:av_byteenable -> Onchip_Memory:byteenable
	wire   [31:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata;                                // DMA_to_Memory_avalon_dma_control_slave_translator:av_writedata -> DMA_to_Memory:slave_writedata
	wire    [1:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_address;                                  // DMA_to_Memory_avalon_dma_control_slave_translator:av_address -> DMA_to_Memory:slave_address
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_write;                                    // DMA_to_Memory_avalon_dma_control_slave_translator:av_write -> DMA_to_Memory:slave_write
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_read;                                     // DMA_to_Memory_avalon_dma_control_slave_translator:av_read -> DMA_to_Memory:slave_read
	wire   [31:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata;                                 // DMA_to_Memory:slave_readdata -> DMA_to_Memory_avalon_dma_control_slave_translator:av_readdata
	wire    [3:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable;                               // DMA_to_Memory_avalon_dma_control_slave_translator:av_byteenable -> DMA_to_Memory:slave_byteenable
	wire   [31:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata;                                // DMA_to_Stream_avalon_dma_control_slave_translator:av_writedata -> DMA_to_Stream:slave_writedata
	wire    [1:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_address;                                  // DMA_to_Stream_avalon_dma_control_slave_translator:av_address -> DMA_to_Stream:slave_address
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_write;                                    // DMA_to_Stream_avalon_dma_control_slave_translator:av_write -> DMA_to_Stream:slave_write
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_read;                                     // DMA_to_Stream_avalon_dma_control_slave_translator:av_read -> DMA_to_Stream:slave_read
	wire   [31:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata;                                 // DMA_to_Stream:slave_readdata -> DMA_to_Stream_avalon_dma_control_slave_translator:av_readdata
	wire    [3:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable;                               // DMA_to_Stream_avalon_dma_control_slave_translator:av_byteenable -> DMA_to_Stream:slave_byteenable
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest;                           // Audio_Video_Config:waitrequest -> Audio_Video_Config_avalon_av_config_slave_translator:av_waitrequest
	wire   [31:0] audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata;                             // Audio_Video_Config_avalon_av_config_slave_translator:av_writedata -> Audio_Video_Config:writedata
	wire    [1:0] audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address;                               // Audio_Video_Config_avalon_av_config_slave_translator:av_address -> Audio_Video_Config:address
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write;                                 // Audio_Video_Config_avalon_av_config_slave_translator:av_write -> Audio_Video_Config:write
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read;                                  // Audio_Video_Config_avalon_av_config_slave_translator:av_read -> Audio_Video_Config:read
	wire   [31:0] audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata;                              // Audio_Video_Config:readdata -> Audio_Video_Config_avalon_av_config_slave_translator:av_readdata
	wire    [3:0] audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable;                            // Audio_Video_Config_avalon_av_config_slave_translator:av_byteenable -> Audio_Video_Config:byteenable
	wire          dma_to_memory_avalon_dma_master_waitrequest;                                                                    // DMA_to_Memory_avalon_dma_master_translator:av_waitrequest -> DMA_to_Memory:master_waitrequest
	wire   [31:0] dma_to_memory_avalon_dma_master_writedata;                                                                      // DMA_to_Memory:master_writedata -> DMA_to_Memory_avalon_dma_master_translator:av_writedata
	wire   [31:0] dma_to_memory_avalon_dma_master_address;                                                                        // DMA_to_Memory:master_address -> DMA_to_Memory_avalon_dma_master_translator:av_address
	wire          dma_to_memory_avalon_dma_master_write;                                                                          // DMA_to_Memory:master_write -> DMA_to_Memory_avalon_dma_master_translator:av_write
	wire          dma_to_stream_avalon_dma_master_waitrequest;                                                                    // DMA_to_Stream_avalon_dma_master_translator:av_waitrequest -> DMA_to_Stream:master_waitrequest
	wire   [31:0] dma_to_stream_avalon_dma_master_address;                                                                        // DMA_to_Stream:master_address -> DMA_to_Stream_avalon_dma_master_translator:av_address
	wire          dma_to_stream_avalon_dma_master_lock;                                                                           // DMA_to_Stream:master_arbiterlock -> DMA_to_Stream_avalon_dma_master_translator:av_lock
	wire          dma_to_stream_avalon_dma_master_read;                                                                           // DMA_to_Stream:master_read -> DMA_to_Stream_avalon_dma_master_translator:av_read
	wire   [31:0] dma_to_stream_avalon_dma_master_readdata;                                                                       // DMA_to_Stream_avalon_dma_master_translator:av_readdata -> DMA_to_Stream:master_readdata
	wire          dma_to_stream_avalon_dma_master_readdatavalid;                                                                  // DMA_to_Stream_avalon_dma_master_translator:av_readdatavalid -> DMA_to_Stream:master_readdatavalid
	wire   [15:0] sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                     // SRAM_Controller_avalon_sram_slave_translator:av_writedata -> SRAM_Controller:writedata
	wire   [19:0] sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                       // SRAM_Controller_avalon_sram_slave_translator:av_address -> SRAM_Controller:address
	wire          sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                         // SRAM_Controller_avalon_sram_slave_translator:av_write -> SRAM_Controller:write
	wire          sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                          // SRAM_Controller_avalon_sram_slave_translator:av_read -> SRAM_Controller:read
	wire   [15:0] sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                      // SRAM_Controller:readdata -> SRAM_Controller_avalon_sram_slave_translator:av_readdata
	wire          sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                 // SRAM_Controller:readdatavalid -> SRAM_Controller_avalon_sram_slave_translator:av_readdatavalid
	wire    [1:0] sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                    // SRAM_Controller_avalon_sram_slave_translator:av_byteenable -> SRAM_Controller:byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                                        // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                                         // CPU_instruction_master_translator:uav_burstcount -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                                          // CPU_instruction_master_translator:uav_writedata -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [15:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                            // CPU_instruction_master_translator:uav_address -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                               // CPU_instruction_master_translator:uav_lock -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                              // CPU_instruction_master_translator:uav_write -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                               // CPU_instruction_master_translator:uav_read -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                                           // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                                        // CPU_instruction_master_translator:uav_debugaccess -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                                         // CPU_instruction_master_translator:uav_byteenable -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                      // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_instruction_master_translator:uav_readdatavalid
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                               // CPU_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                                // CPU_data_master_translator:uav_burstcount -> CPU_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                                 // CPU_data_master_translator:uav_writedata -> CPU_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [15:0] cpu_data_master_translator_avalon_universal_master_0_address;                                                   // CPU_data_master_translator:uav_address -> CPU_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                                      // CPU_data_master_translator:uav_lock -> CPU_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                                     // CPU_data_master_translator:uav_write -> CPU_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                                      // CPU_data_master_translator:uav_read -> CPU_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                                  // CPU_data_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                               // CPU_data_master_translator:uav_debugaccess -> CPU_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                                // CPU_data_master_translator:uav_byteenable -> CPU_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                             // CPU_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_data_master_translator:uav_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // CPU_jtag_debug_module_translator:uav_waitrequest -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> CPU_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> CPU_jtag_debug_module_translator:uav_writedata
	wire   [15:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                     // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> CPU_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                       // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> CPU_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> CPU_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> CPU_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // CPU_jtag_debug_module_translator:uav_readdata -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // CPU_jtag_debug_module_translator:uav_readdatavalid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CPU_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> CPU_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // Onchip_Memory_s1_translator:uav_waitrequest -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Onchip_Memory_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Onchip_Memory_s1_translator:uav_writedata
	wire   [15:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> Onchip_Memory_s1_translator:uav_address
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> Onchip_Memory_s1_translator:uav_write
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Onchip_Memory_s1_translator:uav_lock
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> Onchip_Memory_s1_translator:uav_read
	wire   [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // Onchip_Memory_s1_translator:uav_readdata -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // Onchip_Memory_s1_translator:uav_readdatavalid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Onchip_Memory_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Onchip_Memory_s1_translator:uav_byteenable
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // DMA_to_Memory_avalon_dma_control_slave_translator:uav_waitrequest -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> DMA_to_Memory_avalon_dma_control_slave_translator:uav_burstcount
	wire   [31:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> DMA_to_Memory_avalon_dma_control_slave_translator:uav_writedata
	wire   [15:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> DMA_to_Memory_avalon_dma_control_slave_translator:uav_address
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> DMA_to_Memory_avalon_dma_control_slave_translator:uav_write
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> DMA_to_Memory_avalon_dma_control_slave_translator:uav_lock
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> DMA_to_Memory_avalon_dma_control_slave_translator:uav_read
	wire   [31:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // DMA_to_Memory_avalon_dma_control_slave_translator:uav_readdata -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // DMA_to_Memory_avalon_dma_control_slave_translator:uav_readdatavalid -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> DMA_to_Memory_avalon_dma_control_slave_translator:uav_debugaccess
	wire    [3:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> DMA_to_Memory_avalon_dma_control_slave_translator:uav_byteenable
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // DMA_to_Stream_avalon_dma_control_slave_translator:uav_waitrequest -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> DMA_to_Stream_avalon_dma_control_slave_translator:uav_burstcount
	wire   [31:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> DMA_to_Stream_avalon_dma_control_slave_translator:uav_writedata
	wire   [15:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> DMA_to_Stream_avalon_dma_control_slave_translator:uav_address
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> DMA_to_Stream_avalon_dma_control_slave_translator:uav_write
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> DMA_to_Stream_avalon_dma_control_slave_translator:uav_lock
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> DMA_to_Stream_avalon_dma_control_slave_translator:uav_read
	wire   [31:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // DMA_to_Stream_avalon_dma_control_slave_translator:uav_readdata -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // DMA_to_Stream_avalon_dma_control_slave_translator:uav_readdatavalid -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> DMA_to_Stream_avalon_dma_control_slave_translator:uav_debugaccess
	wire    [3:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> DMA_to_Stream_avalon_dma_control_slave_translator:uav_byteenable
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Audio_Video_Config_avalon_av_config_slave_translator:uav_waitrequest -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Audio_Video_Config_avalon_av_config_slave_translator:uav_burstcount
	wire   [31:0] audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Audio_Video_Config_avalon_av_config_slave_translator:uav_writedata
	wire   [15:0] audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_address -> Audio_Video_Config_avalon_av_config_slave_translator:uav_address
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_write -> Audio_Video_Config_avalon_av_config_slave_translator:uav_write
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Audio_Video_Config_avalon_av_config_slave_translator:uav_lock
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_read -> Audio_Video_Config_avalon_av_config_slave_translator:uav_read
	wire   [31:0] audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // Audio_Video_Config_avalon_av_config_slave_translator:uav_readdata -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Audio_Video_Config_avalon_av_config_slave_translator:uav_readdatavalid -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Audio_Video_Config_avalon_av_config_slave_translator:uav_debugaccess
	wire    [3:0] audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Audio_Video_Config_avalon_av_config_slave_translator:uav_byteenable
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_waitrequest;                               // DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> DMA_to_Memory_avalon_dma_master_translator:uav_waitrequest
	wire    [2:0] dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_burstcount;                                // DMA_to_Memory_avalon_dma_master_translator:uav_burstcount -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_writedata;                                 // DMA_to_Memory_avalon_dma_master_translator:uav_writedata -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_address;                                   // DMA_to_Memory_avalon_dma_master_translator:uav_address -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_lock;                                      // DMA_to_Memory_avalon_dma_master_translator:uav_lock -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_write;                                     // DMA_to_Memory_avalon_dma_master_translator:uav_write -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_read;                                      // DMA_to_Memory_avalon_dma_master_translator:uav_read -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_readdata;                                  // DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> DMA_to_Memory_avalon_dma_master_translator:uav_readdata
	wire          dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_debugaccess;                               // DMA_to_Memory_avalon_dma_master_translator:uav_debugaccess -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_byteenable;                                // DMA_to_Memory_avalon_dma_master_translator:uav_byteenable -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid;                             // DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> DMA_to_Memory_avalon_dma_master_translator:uav_readdatavalid
	wire          dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_waitrequest;                               // DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> DMA_to_Stream_avalon_dma_master_translator:uav_waitrequest
	wire    [2:0] dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_burstcount;                                // DMA_to_Stream_avalon_dma_master_translator:uav_burstcount -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_writedata;                                 // DMA_to_Stream_avalon_dma_master_translator:uav_writedata -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_address;                                   // DMA_to_Stream_avalon_dma_master_translator:uav_address -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_lock;                                      // DMA_to_Stream_avalon_dma_master_translator:uav_lock -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_write;                                     // DMA_to_Stream_avalon_dma_master_translator:uav_write -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_read;                                      // DMA_to_Stream_avalon_dma_master_translator:uav_read -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_readdata;                                  // DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> DMA_to_Stream_avalon_dma_master_translator:uav_readdata
	wire          dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_debugaccess;                               // DMA_to_Stream_avalon_dma_master_translator:uav_debugaccess -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_byteenable;                                // DMA_to_Stream_avalon_dma_master_translator:uav_byteenable -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid;                             // DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> DMA_to_Stream_avalon_dma_master_translator:uav_readdatavalid
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // SRAM_Controller_avalon_sram_slave_translator:uav_waitrequest -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> SRAM_Controller_avalon_sram_slave_translator:uav_burstcount
	wire   [15:0] sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> SRAM_Controller_avalon_sram_slave_translator:uav_writedata
	wire   [31:0] sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> SRAM_Controller_avalon_sram_slave_translator:uav_address
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> SRAM_Controller_avalon_sram_slave_translator:uav_write
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> SRAM_Controller_avalon_sram_slave_translator:uav_lock
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> SRAM_Controller_avalon_sram_slave_translator:uav_read
	wire   [15:0] sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // SRAM_Controller_avalon_sram_slave_translator:uav_readdata -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // SRAM_Controller_avalon_sram_slave_translator:uav_readdatavalid -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SRAM_Controller_avalon_sram_slave_translator:uav_debugaccess
	wire    [1:0] sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> SRAM_Controller_avalon_sram_slave_translator:uav_byteenable
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                               // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                     // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                             // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire   [88:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                      // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                     // addr_router:sink_ready -> CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                      // CPU_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                            // CPU_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                    // CPU_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire   [88:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                             // CPU_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                            // addr_router_001:sink_ready -> CPU_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                       // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire   [88:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router:sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [88:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_001:sink_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [88:0] dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_002:sink_ready -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire   [88:0] dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_003:sink_ready -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire   [88:0] audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_004:sink_ready -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid;                            // DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [100:0] dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data;                             // DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_002:sink_ready -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid;                            // DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [100:0] dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data;                             // DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_003:sink_ready -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire   [82:0] sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_005:sink_ready -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                                              // burst_adapter:source0_endofpacket -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                    // burst_adapter:source0_valid -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                            // burst_adapter:source0_startofpacket -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] burst_adapter_source0_data;                                                                                     // burst_adapter:source0_data -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                    // SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [1:0] burst_adapter_source0_channel;                                                                                  // burst_adapter:source0_channel -> SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                 // rst_controller:reset_out -> Clock_Signals:reset
	wire          clock_signals_sys_clk_reset_reset;                                                                              // Clock_Signals:sys_reset_n -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire          cpu_jtag_debug_module_reset_reset;                                                                              // CPU:jtag_debug_module_resetrequest -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in2]
	wire          rst_controller_001_reset_out_reset;                                                                             // rst_controller_001:reset_out -> [Audio_Video_Config:reset, Audio_Video_Config_avalon_av_config_slave_translator:reset, Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:reset, Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CPU:reset_n, CPU_data_master_translator:reset, CPU_data_master_translator_avalon_universal_master_0_agent:reset, CPU_instruction_master_translator:reset, CPU_instruction_master_translator_avalon_universal_master_0_agent:reset, CPU_jtag_debug_module_translator:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Chroma_Resampler:reset, DMA_to_Memory:reset, DMA_to_Memory_avalon_dma_control_slave_translator:reset, DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:reset, DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, DMA_to_Memory_avalon_dma_master_translator:reset, DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:reset, DMA_to_Stream:reset, DMA_to_Stream_avalon_dma_control_slave_translator:reset, DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:reset, DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, DMA_to_Stream_avalon_dma_master_translator:reset, DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:reset, Dual_Clock_FIFO:reset_stream_in, Onchip_Memory:reset, Onchip_Memory_s1_translator:reset, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:reset, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RGB_Resampler_1:reset, SRAM_Controller:reset, SRAM_Controller_avalon_sram_slave_translator:reset, SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, SRAM_Controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Scaler_0:reset, Scaler_1:reset, Video_Clipper:reset, Video_Decoder:reset, YCrCb_to_RGB_2_0:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_005:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, irq_mapper:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, width_adapter:reset, width_adapter_001:reset]
	wire          rst_controller_002_reset_out_reset;                                                                             // rst_controller_002:reset_out -> [Dual_Clock_FIFO:reset_stream_out, VGA_Controller:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                      // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                              // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire   [88:0] cmd_xbar_demux_src0_data;                                                                                       // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire    [4:0] cmd_xbar_demux_src0_channel;                                                                                    // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                      // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                      // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                              // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire   [88:0] cmd_xbar_demux_src1_data;                                                                                       // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire    [4:0] cmd_xbar_demux_src1_channel;                                                                                    // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                      // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                            // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                  // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                          // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire   [88:0] cmd_xbar_demux_001_src0_data;                                                                                   // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire    [4:0] cmd_xbar_demux_001_src0_channel;                                                                                // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                  // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                            // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                  // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                          // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire   [88:0] cmd_xbar_demux_001_src1_data;                                                                                   // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire    [4:0] cmd_xbar_demux_001_src1_channel;                                                                                // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                  // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                            // cmd_xbar_demux_001:src2_endofpacket -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                  // cmd_xbar_demux_001:src2_valid -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                          // cmd_xbar_demux_001:src2_startofpacket -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_demux_001_src2_data;                                                                                   // cmd_xbar_demux_001:src2_data -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_001_src2_channel;                                                                                // cmd_xbar_demux_001:src2_channel -> DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                            // cmd_xbar_demux_001:src3_endofpacket -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                  // cmd_xbar_demux_001:src3_valid -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                          // cmd_xbar_demux_001:src3_startofpacket -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_demux_001_src3_data;                                                                                   // cmd_xbar_demux_001:src3_data -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_001_src3_channel;                                                                                // cmd_xbar_demux_001:src3_channel -> DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                            // cmd_xbar_demux_001:src4_endofpacket -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                  // cmd_xbar_demux_001:src4_valid -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                          // cmd_xbar_demux_001:src4_startofpacket -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_demux_001_src4_data;                                                                                   // cmd_xbar_demux_001:src4_data -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_001_src4_channel;                                                                                // cmd_xbar_demux_001:src4_channel -> Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                      // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                              // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire   [88:0] rsp_xbar_demux_src0_data;                                                                                       // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [4:0] rsp_xbar_demux_src0_channel;                                                                                    // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                      // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                      // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                              // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire   [88:0] rsp_xbar_demux_src1_data;                                                                                       // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [4:0] rsp_xbar_demux_src1_channel;                                                                                    // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                      // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                            // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                  // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                          // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src0_data;                                                                                   // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [4:0] rsp_xbar_demux_001_src0_channel;                                                                                // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                  // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                            // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                  // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                          // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src1_data;                                                                                   // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire    [4:0] rsp_xbar_demux_001_src1_channel;                                                                                // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                                  // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                            // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                  // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                          // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire   [88:0] rsp_xbar_demux_002_src0_data;                                                                                   // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire    [4:0] rsp_xbar_demux_002_src0_channel;                                                                                // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                  // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                            // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                  // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                          // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire   [88:0] rsp_xbar_demux_003_src0_data;                                                                                   // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire    [4:0] rsp_xbar_demux_003_src0_channel;                                                                                // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                  // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                            // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                  // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                          // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire   [88:0] rsp_xbar_demux_004_src0_data;                                                                                   // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire    [4:0] rsp_xbar_demux_004_src0_channel;                                                                                // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                  // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          addr_router_src_endofpacket;                                                                                    // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                                          // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                                  // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire   [88:0] addr_router_src_data;                                                                                           // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [4:0] addr_router_src_channel;                                                                                        // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                                          // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                   // rsp_xbar_mux:src_endofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                         // rsp_xbar_mux:src_valid -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                 // rsp_xbar_mux:src_startofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] rsp_xbar_mux_src_data;                                                                                          // rsp_xbar_mux:src_data -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_mux_src_channel;                                                                                       // rsp_xbar_mux:src_channel -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                                         // CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                                // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                      // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                              // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire   [88:0] addr_router_001_src_data;                                                                                       // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [4:0] addr_router_001_src_channel;                                                                                    // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                      // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                               // rsp_xbar_mux_001:src_endofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                     // rsp_xbar_mux_001:src_valid -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                             // rsp_xbar_mux_001:src_startofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] rsp_xbar_mux_001_src_data;                                                                                      // rsp_xbar_mux_001:src_data -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_mux_001_src_channel;                                                                                   // rsp_xbar_mux_001:src_channel -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                     // CPU_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                   // cmd_xbar_mux:src_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                         // cmd_xbar_mux:src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                 // cmd_xbar_mux:src_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_mux_src_data;                                                                                          // cmd_xbar_mux:src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_mux_src_channel;                                                                                       // cmd_xbar_mux:src_channel -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                         // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                      // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                            // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                    // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire   [88:0] id_router_src_data;                                                                                             // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [4:0] id_router_src_channel;                                                                                          // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                            // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                               // cmd_xbar_mux_001:src_endofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                     // cmd_xbar_mux_001:src_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                             // cmd_xbar_mux_001:src_startofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] cmd_xbar_mux_001_src_data;                                                                                      // cmd_xbar_mux_001:src_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_mux_001_src_channel;                                                                                   // cmd_xbar_mux_001:src_channel -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                     // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                                  // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                        // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [88:0] id_router_001_src_data;                                                                                         // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [4:0] id_router_001_src_channel;                                                                                      // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                        // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_001_src2_ready;                                                                                  // DMA_to_Memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire          id_router_002_src_endofpacket;                                                                                  // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                        // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                                // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [88:0] id_router_002_src_data;                                                                                         // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [4:0] id_router_002_src_channel;                                                                                      // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                        // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                                  // DMA_to_Stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_003_src_endofpacket;                                                                                  // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                        // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire   [88:0] id_router_003_src_data;                                                                                         // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [4:0] id_router_003_src_channel;                                                                                      // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                        // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                                  // Audio_Video_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                                  // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                        // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire   [88:0] id_router_004_src_data;                                                                                         // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [4:0] id_router_004_src_channel;                                                                                      // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                        // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                            // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                                  // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_005:sink0_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                          // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [100:0] cmd_xbar_demux_002_src0_data;                                                                                   // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_005:sink0_data
	wire    [1:0] cmd_xbar_demux_002_src0_channel;                                                                                // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                                  // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                            // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                                  // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_005:sink1_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                          // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [100:0] cmd_xbar_demux_003_src0_data;                                                                                   // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_005:sink1_data
	wire    [1:0] cmd_xbar_demux_003_src0_channel;                                                                                // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_005:sink1_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                                  // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                            // rsp_xbar_demux_005:src0_endofpacket -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                  // rsp_xbar_demux_005:src0_valid -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                          // rsp_xbar_demux_005:src0_startofpacket -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [100:0] rsp_xbar_demux_005_src0_data;                                                                                   // rsp_xbar_demux_005:src0_data -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] rsp_xbar_demux_005_src0_channel;                                                                                // rsp_xbar_demux_005:src0_channel -> DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                            // rsp_xbar_demux_005:src1_endofpacket -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                                  // rsp_xbar_demux_005:src1_valid -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                                          // rsp_xbar_demux_005:src1_startofpacket -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [100:0] rsp_xbar_demux_005_src1_data;                                                                                   // rsp_xbar_demux_005:src1_data -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] rsp_xbar_demux_005_src1_channel;                                                                                // rsp_xbar_demux_005:src1_channel -> DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_002_src_endofpacket;                                                                                // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                      // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                              // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [100:0] addr_router_002_src_data;                                                                                       // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [1:0] addr_router_002_src_channel;                                                                                    // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                      // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_005_src0_ready;                                                                                  // DMA_to_Memory_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_005:src0_ready
	wire          addr_router_003_src_endofpacket;                                                                                // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                                      // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                              // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [100:0] addr_router_003_src_data;                                                                                       // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire    [1:0] addr_router_003_src_channel;                                                                                    // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                                      // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_demux_005_src1_ready;                                                                                  // DMA_to_Stream_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_005:src1_ready
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                               // cmd_xbar_mux_005:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                                     // cmd_xbar_mux_005:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                             // cmd_xbar_mux_005:src_startofpacket -> width_adapter:in_startofpacket
	wire  [100:0] cmd_xbar_mux_005_src_data;                                                                                      // cmd_xbar_mux_005:src_data -> width_adapter:in_data
	wire    [1:0] cmd_xbar_mux_005_src_channel;                                                                                   // cmd_xbar_mux_005:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                                     // width_adapter:in_ready -> cmd_xbar_mux_005:src_ready
	wire          width_adapter_src_endofpacket;                                                                                  // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                        // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                                // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [82:0] width_adapter_src_data;                                                                                         // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                                        // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire    [1:0] width_adapter_src_channel;                                                                                      // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_005_src_endofpacket;                                                                                  // id_router_005:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_005_src_valid;                                                                                        // id_router_005:src_valid -> width_adapter_001:in_valid
	wire          id_router_005_src_startofpacket;                                                                                // id_router_005:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [82:0] id_router_005_src_data;                                                                                         // id_router_005:src_data -> width_adapter_001:in_data
	wire    [1:0] id_router_005_src_channel;                                                                                      // id_router_005:src_channel -> width_adapter_001:in_channel
	wire          id_router_005_src_ready;                                                                                        // width_adapter_001:in_ready -> id_router_005:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                              // width_adapter_001:out_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                                    // width_adapter_001:out_valid -> rsp_xbar_demux_005:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                            // width_adapter_001:out_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [100:0] width_adapter_001_src_data;                                                                                     // width_adapter_001:out_data -> rsp_xbar_demux_005:sink_data
	wire          width_adapter_001_src_ready;                                                                                    // rsp_xbar_demux_005:sink_ready -> width_adapter_001:out_ready
	wire    [1:0] width_adapter_001_src_channel;                                                                                  // width_adapter_001:out_channel -> rsp_xbar_demux_005:sink_channel
	wire   [31:0] cpu_d_irq_irq;                                                                                                  // irq_mapper:sender_irq -> CPU:d_irq

	niosII_system_Clock_Signals clock_signals (
		.CLOCK_50    (clk_clk),                           //       clk_in_primary.clk
		.reset       (rst_controller_reset_out_reset),    // clk_in_primary_reset.reset
		.sys_clk     (clock_signals_sys_clk_clk),         //              sys_clk.clk
		.sys_reset_n (clock_signals_sys_clk_reset_reset), //        sys_clk_reset.reset_n
		.VGA_CLK     (clock_signals_vga_clk_clk)          //              vga_clk.clk
	);

	niosII_system_Onchip_Memory onchip_memory (
		.clk        (clock_signals_sys_clk_clk),                                  //   clk1.clk
		.address    (onchip_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset)                          // reset1.reset
	);

	niosII_system_CPU cpu (
		.clk                                   (clock_signals_sys_clk_clk),                                          //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                                //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                                 //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	niosII_system_Video_Decoder video_decoder (
		.clk                      (clock_signals_sys_clk_clk),                         //           clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),                //     clock_reset_reset.reset
		.stream_out_ready         (video_decoder_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (video_decoder_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (video_decoder_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (video_decoder_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (video_decoder_avalon_decoder_source_data),          //                      .data
		.TD_CLK27                 (video_decoder_external_interface_TD_CLK27),         //    external_interface.export
		.TD_DATA                  (video_decoder_external_interface_TD_DATA),          //                      .export
		.TD_HS                    (video_decoder_external_interface_TD_HS),            //                      .export
		.TD_VS                    (video_decoder_external_interface_TD_VS),            //                      .export
		.TD_RESET                 (video_decoder_external_interface_TD_RESET),         //                      .export
		.overflow_flag            (video_decoder_external_interface_overflow_flag)     //                      .export
	);

	niosII_system_Video_Clipper video_clipper (
		.clk                      (clock_signals_sys_clk_clk),                         //           clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),                //     clock_reset_reset.reset
		.stream_in_data           (video_decoder_avalon_decoder_source_data),          //   avalon_clipper_sink.data
		.stream_in_startofpacket  (video_decoder_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_in_endofpacket    (video_decoder_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_in_valid          (video_decoder_avalon_decoder_source_valid),         //                      .valid
		.stream_in_ready          (video_decoder_avalon_decoder_source_ready),         //                      .ready
		.stream_out_ready         (video_clipper_avalon_clipper_source_ready),         // avalon_clipper_source.ready
		.stream_out_data          (video_clipper_avalon_clipper_source_data),          //                      .data
		.stream_out_startofpacket (video_clipper_avalon_clipper_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (video_clipper_avalon_clipper_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (video_clipper_avalon_clipper_source_valid)          //                      .valid
	);

	niosII_system_Chroma_Resampler chroma_resampler (
		.clk                      (clock_signals_sys_clk_clk),                           //          clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),                  //    clock_reset_reset.reset
		.stream_in_startofpacket  (scaler_0_avalon_scaler_source_startofpacket),         //   avalon_chroma_sink.startofpacket
		.stream_in_endofpacket    (scaler_0_avalon_scaler_source_endofpacket),           //                     .endofpacket
		.stream_in_valid          (scaler_0_avalon_scaler_source_valid),                 //                     .valid
		.stream_in_ready          (scaler_0_avalon_scaler_source_ready),                 //                     .ready
		.stream_in_data           (scaler_0_avalon_scaler_source_data),                  //                     .data
		.stream_out_ready         (chroma_resampler_avalon_chroma_source_ready),         // avalon_chroma_source.ready
		.stream_out_startofpacket (chroma_resampler_avalon_chroma_source_startofpacket), //                     .startofpacket
		.stream_out_endofpacket   (chroma_resampler_avalon_chroma_source_endofpacket),   //                     .endofpacket
		.stream_out_valid         (chroma_resampler_avalon_chroma_source_valid),         //                     .valid
		.stream_out_data          (chroma_resampler_avalon_chroma_source_data)           //                     .data
	);

	niosII_system_Scaler_0 scaler_0 (
		.clk                      (clock_signals_sys_clk_clk),                         //          clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),                //    clock_reset_reset.reset
		.stream_in_startofpacket  (video_clipper_avalon_clipper_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_clipper_avalon_clipper_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_clipper_avalon_clipper_source_valid),         //                     .valid
		.stream_in_ready          (video_clipper_avalon_clipper_source_ready),         //                     .ready
		.stream_in_data           (video_clipper_avalon_clipper_source_data),          //                     .data
		.stream_out_ready         (scaler_0_avalon_scaler_source_ready),               // avalon_scaler_source.ready
		.stream_out_startofpacket (scaler_0_avalon_scaler_source_startofpacket),       //                     .startofpacket
		.stream_out_endofpacket   (scaler_0_avalon_scaler_source_endofpacket),         //                     .endofpacket
		.stream_out_valid         (scaler_0_avalon_scaler_source_valid),               //                     .valid
		.stream_out_data          (scaler_0_avalon_scaler_source_data)                 //                     .data
	);

	niosII_system_SRAM_Controller sram_controller (
		.clk           (clock_signals_sys_clk_clk),                                                      //        clock_reset.clk
		.reset         (rst_controller_001_reset_out_reset),                                             //  clock_reset_reset.reset
		.SRAM_DQ       (sram_controller_external_interface_DQ),                                          // external_interface.export
		.SRAM_ADDR     (sram_controller_external_interface_ADDR),                                        //                   .export
		.SRAM_LB_N     (sram_controller_external_interface_LB_N),                                        //                   .export
		.SRAM_UB_N     (sram_controller_external_interface_UB_N),                                        //                   .export
		.SRAM_CE_N     (sram_controller_external_interface_CE_N),                                        //                   .export
		.SRAM_OE_N     (sram_controller_external_interface_OE_N),                                        //                   .export
		.SRAM_WE_N     (sram_controller_external_interface_WE_N),                                        //                   .export
		.address       (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	niosII_system_DMA_to_Memory dma_to_memory (
		.clk                  (clock_signals_sys_clk_clk),                                                        //              clock_reset.clk
		.reset                (rst_controller_001_reset_out_reset),                                               //        clock_reset_reset.reset
		.stream_data          (ycrcb_to_rgb_2_0_avalon_streaming_source_data),                                    //          avalon_dma_sink.data
		.stream_startofpacket (ycrcb_to_rgb_2_0_avalon_streaming_source_startofpacket),                           //                         .startofpacket
		.stream_endofpacket   (ycrcb_to_rgb_2_0_avalon_streaming_source_endofpacket),                             //                         .endofpacket
		.stream_valid         (ycrcb_to_rgb_2_0_avalon_streaming_source_valid),                                   //                         .valid
		.stream_ready         (ycrcb_to_rgb_2_0_avalon_streaming_source_ready),                                   //                         .ready
		.slave_address        (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable), //                         .byteenable
		.slave_read           (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),       //                         .read
		.slave_write          (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),      //                         .write
		.slave_writedata      (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),  //                         .writedata
		.slave_readdata       (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),   //                         .readdata
		.master_address       (dma_to_memory_avalon_dma_master_address),                                          //        avalon_dma_master.address
		.master_waitrequest   (dma_to_memory_avalon_dma_master_waitrequest),                                      //                         .waitrequest
		.master_write         (dma_to_memory_avalon_dma_master_write),                                            //                         .write
		.master_writedata     (dma_to_memory_avalon_dma_master_writedata)                                         //                         .writedata
	);

	niosII_system_DMA_to_Stream dma_to_stream (
		.clk                  (clock_signals_sys_clk_clk),                                                        //              clock_reset.clk
		.reset                (rst_controller_001_reset_out_reset),                                               //        clock_reset_reset.reset
		.master_address       (dma_to_stream_avalon_dma_master_address),                                          //        avalon_dma_master.address
		.master_waitrequest   (dma_to_stream_avalon_dma_master_waitrequest),                                      //                         .waitrequest
		.master_arbiterlock   (dma_to_stream_avalon_dma_master_lock),                                             //                         .lock
		.master_read          (dma_to_stream_avalon_dma_master_read),                                             //                         .read
		.master_readdata      (dma_to_stream_avalon_dma_master_readdata),                                         //                         .readdata
		.master_readdatavalid (dma_to_stream_avalon_dma_master_readdatavalid),                                    //                         .readdatavalid
		.slave_address        (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable), //                         .byteenable
		.slave_read           (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),       //                         .read
		.slave_write          (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),      //                         .write
		.slave_writedata      (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),  //                         .writedata
		.slave_readdata       (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),   //                         .readdata
		.stream_ready         (dma_to_stream_avalon_pixel_source_ready),                                          //      avalon_pixel_source.ready
		.stream_data          (dma_to_stream_avalon_pixel_source_data),                                           //                         .data
		.stream_startofpacket (dma_to_stream_avalon_pixel_source_startofpacket),                                  //                         .startofpacket
		.stream_endofpacket   (dma_to_stream_avalon_pixel_source_endofpacket),                                    //                         .endofpacket
		.stream_valid         (dma_to_stream_avalon_pixel_source_valid)                                           //                         .valid
	);

	niosII_system_VGA_Controller vga_controller (
		.clk           (clock_signals_vga_clk_clk),                             //        clock_reset.clk
		.reset         (rst_controller_002_reset_out_reset),                    //  clock_reset_reset.reset
		.data          (dual_clock_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (video_vga_controller_0_external_interface_CLK),         // external_interface.export
		.VGA_HS        (video_vga_controller_0_external_interface_HS),          //                   .export
		.VGA_VS        (video_vga_controller_0_external_interface_VS),          //                   .export
		.VGA_BLANK     (video_vga_controller_0_external_interface_BLANK),       //                   .export
		.VGA_SYNC      (video_vga_controller_0_external_interface_SYNC),        //                   .export
		.VGA_R         (video_vga_controller_0_external_interface_R),           //                   .export
		.VGA_G         (video_vga_controller_0_external_interface_G),           //                   .export
		.VGA_B         (video_vga_controller_0_external_interface_B)            //                   .export
	);

	niosII_system_Dual_Clock_FIFO dual_clock_fifo (
		.clk_stream_in            (clock_signals_sys_clk_clk),                             //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_001_reset_out_reset),                    //   clock_stream_in_reset.reset
		.clk_stream_out           (clock_signals_vga_clk_clk),                             //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                    //  clock_stream_out_reset.reset
		.stream_in_ready          (scaler_1_avalon_scaler_source_ready),                   //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (scaler_1_avalon_scaler_source_startofpacket),           //                        .startofpacket
		.stream_in_endofpacket    (scaler_1_avalon_scaler_source_endofpacket),             //                        .endofpacket
		.stream_in_valid          (scaler_1_avalon_scaler_source_valid),                   //                        .valid
		.stream_in_data           (scaler_1_avalon_scaler_source_data),                    //                        .data
		.stream_out_ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (dual_clock_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	niosII_system_Audio_Video_Config audio_video_config (
		.clk         (clock_signals_sys_clk_clk),                                                            //            clock_reset.clk
		.reset       (rst_controller_001_reset_out_reset),                                                   //      clock_reset_reset.reset
		.address     (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address),     // avalon_av_config_slave.address
		.byteenable  (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),  //                       .byteenable
		.read        (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read),        //                       .read
		.write       (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write),       //                       .write
		.writedata   (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),   //                       .writedata
		.readdata    (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),    //                       .readdata
		.waitrequest (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_video_config_external_interface_SDAT),                                           //     external_interface.export
		.I2C_SCLK    (audio_video_config_external_interface_SCLK)                                            //                       .export
	);

	YCrCb_444_to_24_RGB #(
		.IW  (23),
		.OW  (23),
		.EIW (1),
		.EOW (1)
	) ycrcb_to_rgb_2_0 (
		.clk                      (clock_signals_sys_clk_clk),                              //                   clock.clk
		.reset                    (rst_controller_001_reset_out_reset),                     //                   reset.reset
		.stream_in_data           (chroma_resampler_avalon_chroma_source_data),             //   avalon_streaming_sink.data
		.stream_in_startofpacket  (chroma_resampler_avalon_chroma_source_startofpacket),    //                        .startofpacket
		.stream_in_endofpacket    (chroma_resampler_avalon_chroma_source_endofpacket),      //                        .endofpacket
		.stream_in_valid          (chroma_resampler_avalon_chroma_source_valid),            //                        .valid
		.stream_in_ready          (chroma_resampler_avalon_chroma_source_ready),            //                        .ready
		.stream_out_ready         (ycrcb_to_rgb_2_0_avalon_streaming_source_ready),         // avalon_streaming_source.ready
		.stream_out_data          (ycrcb_to_rgb_2_0_avalon_streaming_source_data),          //                        .data
		.stream_out_startofpacket (ycrcb_to_rgb_2_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (ycrcb_to_rgb_2_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (ycrcb_to_rgb_2_0_avalon_streaming_source_valid)          //                        .valid
	);

	niosII_system_Scaler_1 scaler_1 (
		.clk                      (clock_signals_sys_clk_clk),                       //          clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),              //    clock_reset_reset.reset
		.stream_in_startofpacket  (rgb_resampler_1_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (rgb_resampler_1_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (rgb_resampler_1_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (rgb_resampler_1_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (rgb_resampler_1_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (scaler_1_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (scaler_1_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (scaler_1_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (scaler_1_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (scaler_1_avalon_scaler_source_data)               //                     .data
	);

	niosII_system_RGB_Resampler_1 rgb_resampler_1 (
		.clk                      (clock_signals_sys_clk_clk),                       //       clock_reset.clk
		.reset                    (rst_controller_001_reset_out_reset),              // clock_reset_reset.reset
		.stream_in_startofpacket  (dma_to_stream_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (dma_to_stream_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (dma_to_stream_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (dma_to_stream_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (dma_to_stream_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (rgb_resampler_1_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_resampler_1_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (rgb_resampler_1_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (rgb_resampler_1_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (rgb_resampler_1_avalon_rgb_source_data)           //                  .data
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                 //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                        //                     reset.reset
		.uav_address           (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_byteenable         (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_readdatavalid      (),                                                                          //               (terminated)
		.av_write              (1'b0),                                                                      //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_data_master_translator (
		.clk                   (clock_signals_sys_clk_clk),                                          //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                 //                     reset.reset
		.uav_address           (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_data_master_read),                                               //                          .read
		.av_readdata           (cpu_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_data_master_write),                                              //                          .write
		.av_writedata          (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_readdatavalid      (),                                                                   //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                               //                    reset.reset
		.uav_address           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_s1_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dma_to_memory_avalon_dma_control_slave_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                                //                    reset.reset
		.uav_address           (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (dma_to_memory_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer      (),                                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                                  //              (terminated)
		.av_lock               (),                                                                                                  //              (terminated)
		.av_chipselect         (),                                                                                                  //              (terminated)
		.av_clken              (),                                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dma_to_stream_avalon_dma_control_slave_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                                //                    reset.reset
		.uav_address           (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (dma_to_stream_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer      (),                                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                                  //              (terminated)
		.av_lock               (),                                                                                                  //              (terminated)
		.av_chipselect         (),                                                                                                  //              (terminated)
		.av_clken              (),                                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_video_config_avalon_av_config_slave_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                                   //                    reset.reset
		.uav_address           (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (audio_video_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                                     //              (terminated)
		.av_lock               (),                                                                                                     //              (terminated)
		.av_chipselect         (),                                                                                                     //              (terminated)
		.av_clken              (),                                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                                      //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_to_memory_avalon_dma_master_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                          //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                 //                     reset.reset
		.uav_address           (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (dma_to_memory_avalon_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (dma_to_memory_avalon_dma_master_waitrequest),                                        //                          .waitrequest
		.av_write              (dma_to_memory_avalon_dma_master_write),                                              //                          .write
		.av_writedata          (dma_to_memory_avalon_dma_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                                               //               (terminated)
		.av_read               (1'b0),                                                                               //               (terminated)
		.av_readdata           (),                                                                                   //               (terminated)
		.av_readdatavalid      (),                                                                                   //               (terminated)
		.av_lock               (1'b0),                                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                                               //               (terminated)
		.uav_clken             (),                                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_to_stream_avalon_dma_master_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                          //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                 //                     reset.reset
		.uav_address           (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (dma_to_stream_avalon_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (dma_to_stream_avalon_dma_master_waitrequest),                                        //                          .waitrequest
		.av_read               (dma_to_stream_avalon_dma_master_read),                                               //                          .read
		.av_readdata           (dma_to_stream_avalon_dma_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (dma_to_stream_avalon_dma_master_readdatavalid),                                      //                          .readdatavalid
		.av_lock               (dma_to_stream_avalon_dma_master_lock),                                               //                          .lock
		.av_burstcount         (1'b1),                                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                                               //               (terminated)
		.av_write              (1'b0),                                                                               //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                                               //               (terminated)
		.uav_clken             (),                                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (20),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sram_controller_avalon_sram_slave_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sram_controller_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer      (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_lock               (),                                                                                             //              (terminated)
		.av_chipselect         (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_debugaccess        (),                                                                                             //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_THREAD_ID_H           (79),
		.PKT_THREAD_ID_L           (79),
		.PKT_CACHE_H               (86),
		.PKT_CACHE_L               (83),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clock_signals_sys_clk_clk),                                                          //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.av_address       (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_src_valid),                                                             //        rp.valid
		.rp_data          (rsp_xbar_mux_src_data),                                                              //          .data
		.rp_channel       (rsp_xbar_mux_src_channel),                                                           //          .channel
		.rp_startofpacket (rsp_xbar_mux_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_src_endofpacket),                                                       //          .endofpacket
		.rp_ready         (rsp_xbar_mux_src_ready)                                                              //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_THREAD_ID_H           (79),
		.PKT_THREAD_ID_L           (79),
		.PKT_CACHE_H               (86),
		.PKT_CACHE_L               (83),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clock_signals_sys_clk_clk),                                                   //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.av_address       (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                  //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                   //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                          //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                            //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                   //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                          //                .channel
		.rf_sink_ready           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                          //       clk_reset.reset
		.m0_address              (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                                             //                .channel
		.rf_sink_ready           (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                          // clk_reset.reset
		.in_data           (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                                        // (terminated)
		.csr_readdata      (),                                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                        // (terminated)
		.almost_full_data  (),                                                                                                            // (terminated)
		.almost_empty_data (),                                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                                        // (terminated)
		.out_empty         (),                                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                                        // (terminated)
		.out_error         (),                                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                                        // (terminated)
		.out_channel       ()                                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                          //       clk_reset.reset
		.m0_address              (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                             //                .channel
		.rf_sink_ready           (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                          // clk_reset.reset
		.in_data           (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                                        // (terminated)
		.csr_readdata      (),                                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                        // (terminated)
		.almost_full_data  (),                                                                                                            // (terminated)
		.almost_empty_data (),                                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                                        // (terminated)
		.out_empty         (),                                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                                        // (terminated)
		.out_error         (),                                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                                        // (terminated)
		.out_channel       ()                                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                                                //                .channel
		.rf_sink_ready           (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                                           // (terminated)
		.csr_readdata      (),                                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                           // (terminated)
		.almost_full_data  (),                                                                                                               // (terminated)
		.almost_empty_data (),                                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                                           // (terminated)
		.out_empty         (),                                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                                           // (terminated)
		.out_error         (),                                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                                           // (terminated)
		.out_channel       ()                                                                                                                // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (90),
		.PKT_THREAD_ID_H           (91),
		.PKT_THREAD_ID_L           (91),
		.PKT_CACHE_H               (98),
		.PKT_CACHE_L               (95),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent (
		.clk              (clock_signals_sys_clk_clk),                                                                   //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.av_address       (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_005_src0_valid),                                                               //        rp.valid
		.rp_data          (rsp_xbar_demux_005_src0_data),                                                                //          .data
		.rp_channel       (rsp_xbar_demux_005_src0_channel),                                                             //          .channel
		.rp_startofpacket (rsp_xbar_demux_005_src0_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),                                                         //          .endofpacket
		.rp_ready         (rsp_xbar_demux_005_src0_ready)                                                                //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (90),
		.PKT_THREAD_ID_H           (91),
		.PKT_THREAD_ID_L           (91),
		.PKT_CACHE_H               (98),
		.PKT_CACHE_L               (95),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent (
		.clk              (clock_signals_sys_clk_clk),                                                                   //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.av_address       (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_005_src1_valid),                                                               //        rp.valid
		.rp_data          (rsp_xbar_demux_005_src1_data),                                                                //          .data
		.rp_channel       (rsp_xbar_demux_005_src1_channel),                                                             //          .channel
		.rp_startofpacket (rsp_xbar_demux_005_src1_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),                                                         //          .endofpacket
		.rp_ready         (rsp_xbar_demux_005_src1_ready)                                                                //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (71),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (72),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                            //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                            //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                             //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                                          //                .channel
		.rf_sink_ready           (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	niosII_system_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	niosII_system_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                              //          .endofpacket
	);

	niosII_system_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	niosII_system_id_router id_router_001 (
		.sink_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                     //       src.ready
		.src_valid          (id_router_001_src_valid),                                                     //          .valid
		.src_data           (id_router_001_src_data),                                                      //          .data
		.src_channel        (id_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                //          .endofpacket
	);

	niosII_system_id_router_002 id_router_002 (
		.sink_ready         (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_to_memory_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                                // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                           //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                           //          .valid
		.src_data           (id_router_002_src_data),                                                                            //          .data
		.src_channel        (id_router_002_src_channel),                                                                         //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                                   //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                                      //          .endofpacket
	);

	niosII_system_id_router_002 id_router_003 (
		.sink_ready         (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_to_stream_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                                // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                           //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                           //          .valid
		.src_data           (id_router_003_src_data),                                                                            //          .data
		.src_channel        (id_router_003_src_channel),                                                                         //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                                   //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                                      //          .endofpacket
	);

	niosII_system_id_router_002 id_router_004 (
		.sink_ready         (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_video_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                              //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                              //          .valid
		.src_data           (id_router_004_src_data),                                                                               //          .data
		.src_channel        (id_router_004_src_channel),                                                                            //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                                         //          .endofpacket
	);

	niosII_system_addr_router_002 addr_router_002 (
		.sink_ready         (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_to_memory_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                                   //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                                   //          .valid
		.src_data           (addr_router_002_src_data),                                                                    //          .data
		.src_channel        (addr_router_002_src_channel),                                                                 //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                              //          .endofpacket
	);

	niosII_system_addr_router_002 addr_router_003 (
		.sink_ready         (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_to_stream_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                                   //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                                   //          .valid
		.src_data           (addr_router_003_src_data),                                                                    //          .data
		.src_channel        (addr_router_003_src_channel),                                                                 //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                              //          .endofpacket
	);

	niosII_system_id_router_005 id_router_005 (
		.sink_ready         (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_controller_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                      //          .valid
		.src_data           (id_router_005_src_data),                                                                       //          .data
		.src_channel        (id_router_005_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                                 //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (2),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter (
		.clk                   (clock_signals_sys_clk_clk),           //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (~clock_signals_sys_clk_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (~clock_signals_sys_clk_reset_reset), // reset_in1.reset
		.reset_in2  (cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.clk        (clock_signals_sys_clk_clk),          //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~clock_signals_sys_clk_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                     // reset_in1.reset
		.reset_in2  (cpu_jtag_debug_module_reset_reset),  // reset_in2.reset
		.clk        (clock_signals_vga_clk_clk),          //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	niosII_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clock_signals_sys_clk_clk),          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (addr_router_src_ready),              //      sink.ready
		.sink_channel       (addr_router_src_channel),            //          .channel
		.sink_data          (addr_router_src_data),               //          .data
		.sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid         (addr_router_src_valid),              //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	niosII_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clock_signals_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clock_signals_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_demux rsp_xbar_demux (
		.clk                (clock_signals_sys_clk_clk),          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	niosII_system_cmd_xbar_demux rsp_xbar_demux_001 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clock_signals_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clock_signals_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux_005 cmd_xbar_mux_005 (
		.clk                 (clock_signals_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src0_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_005 rsp_xbar_demux_005 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (100),
		.IN_PKT_RESPONSE_STATUS_L      (99),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (101),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (82),
		.OUT_PKT_RESPONSE_STATUS_L     (81),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (83),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (clock_signals_sys_clk_clk),          //       clk.clk
		.reset                (rst_controller_001_reset_out_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_mux_005_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_005_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_005_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_005_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_005_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_005_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (82),
		.IN_PKT_RESPONSE_STATUS_L      (81),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (83),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (100),
		.OUT_PKT_RESPONSE_STATUS_L     (99),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (101),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (clock_signals_sys_clk_clk),           //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_005_src_valid),             //      sink.valid
		.in_channel           (id_router_005_src_channel),           //          .channel
		.in_startofpacket     (id_router_005_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_005_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_005_src_ready),             //          .ready
		.in_data              (id_router_005_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	niosII_system_irq_mapper irq_mapper (
		.clk        (clock_signals_sys_clk_clk),          //       clk.clk
		.reset      (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu_d_irq_irq)                       //    sender.irq
	);

endmodule
